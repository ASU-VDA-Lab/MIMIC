module real_jpeg_9743_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_314, n_11, n_14, n_313, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_314;
input n_11;
input n_14;
input n_313;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_1),
.A2(n_49),
.B1(n_64),
.B2(n_65),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_49),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_2),
.A2(n_11),
.B(n_28),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_3),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_77),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_77),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_77),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g98 ( 
.A(n_4),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_6),
.A2(n_35),
.B1(n_64),
.B2(n_65),
.Y(n_232)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_31),
.B(n_62),
.C(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_9),
.B(n_31),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_10),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_10),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_59),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_59),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_31),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_11),
.B(n_31),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_11),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_11),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_11),
.A2(n_27),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_11),
.B(n_27),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_11),
.B(n_50),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_121),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_12),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_108),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_108),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_108),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_14),
.A2(n_42),
.B1(n_64),
.B2(n_65),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_42),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_15),
.A2(n_64),
.B1(n_65),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_15),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_101),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_101),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_101),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_16),
.A2(n_64),
.B1(n_65),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_16),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_137),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_16),
.A2(n_27),
.B1(n_28),
.B2(n_137),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_16),
.A2(n_40),
.B1(n_41),
.B2(n_137),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_17),
.A2(n_64),
.B1(n_65),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_17),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_96),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_96),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_17),
.A2(n_40),
.B1(n_41),
.B2(n_96),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_84),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_82),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_69),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_69),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_51),
.B1(n_52),
.B2(n_68),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_25),
.A2(n_30),
.B1(n_55),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_25),
.A2(n_30),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_25),
.A2(n_30),
.B1(n_146),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_25),
.A2(n_30),
.B1(n_162),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_25),
.A2(n_30),
.B1(n_202),
.B2(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_25),
.A2(n_30),
.B1(n_213),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_25),
.A2(n_30),
.B1(n_239),
.B2(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_25),
.A2(n_30),
.B1(n_81),
.B2(n_257),
.Y(n_273)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_27),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_29),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_30),
.B(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_31),
.B(n_33),
.Y(n_150)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_32),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_44),
.B1(n_47),
.B2(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_45),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_41),
.A2(n_45),
.B(n_121),
.C(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_43),
.A2(n_50),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_47),
.B1(n_58),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_44),
.A2(n_47),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_44),
.A2(n_47),
.B1(n_217),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_44),
.A2(n_47),
.B1(n_242),
.B2(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_44),
.A2(n_47),
.B1(n_76),
.B2(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.C(n_60),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_54),
.B1(n_60),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_60),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_63),
.B(n_67),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_63),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_61),
.A2(n_63),
.B1(n_107),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_61),
.A2(n_63),
.B1(n_134),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_61),
.A2(n_63),
.B1(n_142),
.B2(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_61),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_61),
.A2(n_63),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_61),
.A2(n_63),
.B1(n_225),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_61),
.A2(n_63),
.B1(n_234),
.B2(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_61),
.A2(n_63),
.B1(n_67),
.B2(n_266),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_63),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_63),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_64),
.B(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_64),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.C(n_78),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_300),
.Y(n_305)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_75),
.C(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_75),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_75),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_78),
.B(n_305),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_297),
.A3(n_306),
.B1(n_309),
.B2(n_310),
.C(n_313),
.Y(n_84)
);

AOI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_250),
.A3(n_285),
.B1(n_291),
.B2(n_296),
.C(n_314),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_207),
.C(n_246),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_177),
.B(n_206),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_156),
.B(n_176),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_139),
.B(n_155),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_128),
.B(n_138),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_114),
.B(n_127),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_93),
.B(n_102),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_97),
.A2(n_98),
.B1(n_154),
.B2(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_118),
.B1(n_119),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_109),
.B2(n_113),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_113),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_122),
.B(n_126),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_120),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_119),
.B1(n_136),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_118),
.A2(n_119),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_118),
.A2(n_119),
.B1(n_188),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_118),
.A2(n_119),
.B1(n_222),
.B2(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_118),
.A2(n_119),
.B(n_232),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_130),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_140),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.CI(n_135),
.CON(n_131),
.SN(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_140),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_143),
.CI(n_147),
.CON(n_140),
.SN(n_140)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_145),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_152),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_158),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_169),
.B2(n_170),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_172),
.C(n_174),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_163),
.B1(n_164),
.B2(n_168),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_161),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_166),
.C(n_168),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_171),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_178),
.B(n_179),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_192),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_181),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_181),
.B(n_191),
.C(n_192),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_186),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_189),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_203),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_200),
.B2(n_201),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_200),
.C(n_203),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_205),
.Y(n_216)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_208),
.A2(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_227),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_209),
.B(n_227),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_220),
.C(n_226),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_219),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_218),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_212),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_SL g244 ( 
.A(n_214),
.B(n_218),
.C(n_219),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_226),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_223),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_244),
.B2(n_245),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_230),
.B(n_235),
.C(n_245),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_233),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_240),
.C(n_243),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_238),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_247),
.B(n_248),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_269),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_251),
.B(n_269),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_262),
.C(n_268),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_252),
.A2(n_253),
.B1(n_262),
.B2(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_258),
.C(n_261),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_256),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_262),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_264),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_263),
.A2(n_279),
.B(n_281),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_265),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_265),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_283),
.B2(n_284),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_276),
.C(n_284),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B(n_275),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_274),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_299),
.C(n_303),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_275),
.B(n_299),
.CI(n_303),
.CON(n_308),
.SN(n_308)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_281),
.B2(n_282),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_279),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_292),
.B(n_295),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_304),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_304),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_307),
.B(n_308),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_308),
.Y(n_312)
);


endmodule