module fake_jpeg_21179_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_29),
.B1(n_24),
.B2(n_31),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_48),
.B1(n_39),
.B2(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_47),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_29),
.B1(n_24),
.B2(n_32),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_29),
.B1(n_32),
.B2(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_63),
.A2(n_82),
.B1(n_53),
.B2(n_46),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_68),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_16),
.B1(n_31),
.B2(n_18),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_53),
.B1(n_41),
.B2(n_46),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_80),
.B1(n_85),
.B2(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_54),
.B(n_38),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_39),
.B1(n_16),
.B2(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_23),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_16),
.B1(n_22),
.B2(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_38),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_73),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_87),
.B(n_25),
.Y(n_125)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_47),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_75),
.Y(n_119)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_61),
.B1(n_87),
.B2(n_60),
.Y(n_121)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_111),
.B(n_112),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_83),
.B1(n_46),
.B2(n_74),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_135),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_61),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_124),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_88),
.B1(n_94),
.B2(n_104),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_86),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_122),
.A2(n_132),
.B(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_76),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_88),
.B(n_17),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_104),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_78),
.B1(n_83),
.B2(n_65),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_92),
.B(n_89),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_128),
.B(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_38),
.C(n_47),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_109),
.C(n_102),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_59),
.B1(n_44),
.B2(n_43),
.Y(n_131)
);

NAND2x1p5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_19),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_72),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_44),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_96),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_138),
.C(n_135),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_22),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_19),
.Y(n_142)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_110),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_142),
.B(n_125),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_149),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_92),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_146),
.B(n_161),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_111),
.C(n_108),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_155),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_94),
.C(n_95),
.Y(n_153)
);

AO22x2_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_103),
.B1(n_72),
.B2(n_106),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_160),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_21),
.B(n_27),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_142),
.B(n_118),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_21),
.B(n_103),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_163),
.C(n_151),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_98),
.B1(n_101),
.B2(n_107),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_93),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_166),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_107),
.B1(n_101),
.B2(n_98),
.Y(n_165)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_23),
.C(n_100),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_134),
.B1(n_115),
.B2(n_4),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_28),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_174),
.B(n_179),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_178),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_148),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_115),
.B(n_133),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_165),
.B1(n_144),
.B2(n_5),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_19),
.B1(n_23),
.B2(n_28),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_28),
.Y(n_189)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_19),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_191),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_193),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_26),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_194),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_201),
.A2(n_211),
.B1(n_213),
.B2(n_174),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_154),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_204),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_154),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_149),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_210),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_163),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_164),
.B1(n_155),
.B2(n_153),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_155),
.B1(n_166),
.B2(n_158),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_216),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_155),
.C(n_2),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_183),
.C(n_176),
.Y(n_229)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

OAI22x1_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_172),
.B1(n_177),
.B2(n_179),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_221),
.A2(n_216),
.B1(n_212),
.B2(n_207),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_224),
.Y(n_243)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_177),
.B(n_194),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_226),
.A2(n_213),
.B(n_199),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_211),
.A2(n_188),
.B1(n_175),
.B2(n_187),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_232),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_197),
.C(n_204),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_188),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_209),
.B(n_184),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_231),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_175),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_8),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_219),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_242),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_238),
.A2(n_229),
.B1(n_228),
.B2(n_210),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_182),
.B(n_191),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g242 ( 
.A(n_230),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_182),
.Y(n_244)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_221),
.B1(n_222),
.B2(n_185),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_245),
.A2(n_250),
.B1(n_8),
.B2(n_9),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_255),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_237),
.B1(n_240),
.B2(n_10),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_235),
.A2(n_218),
.B1(n_219),
.B2(n_5),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_253),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_218),
.B1(n_2),
.B2(n_5),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_0),
.C(n_6),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_255),
.C(n_247),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_0),
.B(n_7),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_251),
.B1(n_11),
.B2(n_12),
.Y(n_268)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_8),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_260),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_9),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_263),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_249),
.B(n_10),
.Y(n_262)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_254),
.B(n_245),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_259),
.B(n_257),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_10),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_259),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_271),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_263),
.B(n_11),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_266),
.B(n_267),
.C(n_268),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_273),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_13),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_275),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_14),
.Y(n_278)
);


endmodule