module fake_jpeg_16747_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx8_ASAP7_75t_SL g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_56),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_37),
.C(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_60),
.Y(n_83)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_44),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_51),
.B1(n_49),
.B2(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_50),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_46),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_85),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_42),
.Y(n_96)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_93),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_60),
.B1(n_45),
.B2(n_66),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_62),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_84),
.B1(n_48),
.B2(n_42),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_72),
.B1(n_83),
.B2(n_81),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_92),
.B(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_102),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_SL g105 ( 
.A1(n_97),
.A2(n_93),
.B(n_91),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_106),
.C(n_107),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_88),
.C(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_100),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_111),
.B1(n_99),
.B2(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_100),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_113),
.B(n_8),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_110),
.A2(n_22),
.B1(n_36),
.B2(n_10),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_26),
.CI(n_14),
.CON(n_116),
.SN(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

AOI21x1_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_116),
.B(n_15),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_28),
.B1(n_16),
.B2(n_18),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_73),
.A3(n_20),
.B1(n_21),
.B2(n_25),
.C1(n_27),
.C2(n_29),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_31),
.B(n_32),
.Y(n_121)
);


endmodule