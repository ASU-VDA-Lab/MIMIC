module fake_jpeg_17023_n_29 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

INVx3_ASAP7_75t_SL g10 ( 
.A(n_9),
.Y(n_10)
);

CKINVDCx14_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_L g12 ( 
.A1(n_3),
.A2(n_1),
.B1(n_8),
.B2(n_0),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_6),
.A2(n_9),
.B1(n_2),
.B2(n_8),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_18),
.C(n_11),
.Y(n_19)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_19),
.B(n_18),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_10),
.C(n_11),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_10),
.C(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_25),
.B1(n_13),
.B2(n_14),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_12),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_15),
.B1(n_20),
.B2(n_22),
.Y(n_27)
);

AOI322xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.C1(n_17),
.C2(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_26),
.Y(n_29)
);


endmodule