module fake_ariane_3140_n_5439 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_640, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_598, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_620, n_228, n_325, n_276, n_93, n_636, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_588, n_638, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_5439);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_640;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_5439;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_5402;
wire n_2182;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_2482;
wire n_1682;
wire n_958;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_786;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_3482;
wire n_5403;
wire n_823;
wire n_1900;
wire n_4268;
wire n_863;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_899;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_661;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_4476;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_1213;
wire n_2382;
wire n_780;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_1140;
wire n_3458;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5391;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_992;
wire n_966;
wire n_3549;
wire n_3914;
wire n_1692;
wire n_2611;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5179;
wire n_2435;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_4254;
wire n_646;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_670;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_5088;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_1053;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_4292;
wire n_2118;
wire n_688;
wire n_1490;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_1104;
wire n_986;
wire n_887;
wire n_2125;
wire n_1156;
wire n_5123;
wire n_4974;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1498;
wire n_1188;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_3944;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_655;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_951;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_704;
wire n_2958;
wire n_1714;
wire n_1044;
wire n_4429;
wire n_5435;
wire n_3340;
wire n_5053;
wire n_1243;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_811;
wire n_791;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_3450;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_906;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_3740;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_1517;
wire n_2647;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_3380;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_5377;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5426;
wire n_4093;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_2963;
wire n_2561;
wire n_1056;
wire n_674;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_848;
wire n_5125;
wire n_4922;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_724;
wire n_2931;
wire n_3433;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_3786;
wire n_875;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_793;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_3610;
wire n_2443;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5388;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_5196;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_3633;
wire n_857;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_840;
wire n_2324;
wire n_5283;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5040;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_5399;
wire n_658;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_1168;
wire n_4663;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3895;
wire n_3707;
wire n_1091;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_5304;
wire n_5437;
wire n_1581;
wire n_946;
wire n_3058;
wire n_757;
wire n_2047;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_5355;
wire n_998;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_963;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_4016;
wire n_3334;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_4591;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_1233;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_675;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_1169;
wire n_789;
wire n_3181;
wire n_1916;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_5360;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_2221;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_2634;
wire n_2746;
wire n_645;
wire n_5098;
wire n_721;
wire n_1084;
wire n_1276;
wire n_5145;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_2458;
wire n_3150;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_4498;
wire n_772;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_3234;
wire n_1351;
wire n_2216;
wire n_2426;
wire n_652;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_3391;
wire n_912;
wire n_4786;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_5408;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_967;
wire n_5130;
wire n_4175;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2601;
wire n_2172;
wire n_1880;
wire n_2365;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_1226;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_3257;
wire n_3730;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5159;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_926;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_855;
wire n_2059;
wire n_4713;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_5376;
wire n_3508;
wire n_4129;
wire n_1105;
wire n_3599;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_983;
wire n_699;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_729;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_3568;
wire n_3216;
wire n_2555;
wire n_2708;
wire n_735;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_3791;
wire n_982;
wire n_915;
wire n_2008;
wire n_4989;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_1171;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5256;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_3735;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_5364;
wire n_3302;
wire n_2486;
wire n_1897;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_5222;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_3408;
wire n_2884;
wire n_1293;
wire n_961;
wire n_726;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_5378;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5293;
wire n_779;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_3738;
wire n_894;
wire n_1380;
wire n_2020;
wire n_2310;
wire n_3600;
wire n_1023;
wire n_914;
wire n_689;
wire n_5382;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_4370;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_962;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_1968;
wire n_918;
wire n_5020;
wire n_673;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_4333;
wire n_5339;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_3481;
wire n_5101;
wire n_2236;
wire n_692;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_1204;
wire n_2428;
wire n_994;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_856;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_2402;
wire n_1458;
wire n_679;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_3687;
wire n_2787;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_2375;
wire n_3278;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_5143;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_5425;
wire n_5273;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_5002;
wire n_831;
wire n_3681;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_671;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_684;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_662;
wire n_3461;
wire n_1410;
wire n_2297;
wire n_939;
wire n_4203;
wire n_5400;
wire n_1325;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_3763;
wire n_933;
wire n_3499;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_5375;
wire n_5438;
wire n_1264;
wire n_4958;
wire n_1827;
wire n_4149;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_2423;
wire n_2208;
wire n_1421;
wire n_5422;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_1383;
wire n_4259;
wire n_2030;
wire n_850;
wire n_4299;
wire n_2407;
wire n_690;
wire n_5367;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_1246;
wire n_5265;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_1196;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_1187;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_766;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_665;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_672;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_821;
wire n_770;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_1112;
wire n_700;
wire n_4174;
wire n_5131;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_5333;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_712;
wire n_909;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_964;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_1095;
wire n_3078;
wire n_3971;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_677;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_5420;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_5406;
wire n_4328;
wire n_1854;
wire n_666;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_5428;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_1078;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_4766;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_5431;
wire n_643;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_686;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_5369;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5270;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_879;
wire n_4561;
wire n_1541;
wire n_3291;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_1185;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_1090;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_2692;
wire n_683;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_2645;
wire n_2553;
wire n_1420;
wire n_4711;
wire n_2749;
wire n_660;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_5223;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_1022;
wire n_3532;
wire n_5154;
wire n_2609;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_4138;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_697;
wire n_4620;
wire n_5397;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_880;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_975;
wire n_1645;
wire n_932;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_2465;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_4858;
wire n_1445;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_969;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_1271;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_1285;
wire n_733;
wire n_761;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_648;
wire n_3273;
wire n_2918;
wire n_835;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_654;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_977;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_723;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_4886;
wire n_5172;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1982;
wire n_5311;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_4483;
wire n_3061;
wire n_3504;
wire n_2587;
wire n_4693;
wire n_1043;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_664;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_2135;
wire n_4475;
wire n_5432;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_1988;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_4768;
wire n_1889;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_2727;
wire n_942;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_5418;
wire n_5019;
wire n_1819;
wire n_3095;
wire n_947;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_696;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2549;
wire n_2499;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_669;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_824;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_815;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_965;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_713;
wire n_3179;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_927;
wire n_3699;
wire n_706;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_5335;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_3276;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_647;
wire n_2027;
wire n_2932;
wire n_3118;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_1467;
wire n_5209;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_681;
wire n_3286;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_5219;
wire n_920;
wire n_3951;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_861;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_657;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_1030;
wire n_5181;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_876;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_3694;
wire n_771;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_3543;
wire n_2945;
wire n_1324;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_2698;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_2352;
wire n_5201;
wire n_790;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_4544;
wire n_1773;
wire n_3175;
wire n_2666;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_3790;
wire n_907;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_2174;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_2865;
wire n_973;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_5387;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_653;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_2169;
wire n_5133;
wire n_5305;
wire n_2175;
wire n_1625;
wire n_4578;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_2395;
wire n_2868;
wire n_4057;
wire n_1530;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_668;
wire n_2111;
wire n_3743;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_694;
wire n_4749;
wire n_1845;
wire n_921;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_741;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_865;
wire n_5034;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_1474;
wire n_937;
wire n_1631;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_1249;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

INVxp67_ASAP7_75t_L g643 ( 
.A(n_272),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_86),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_242),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_273),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_58),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_394),
.Y(n_648)
);

BUFx10_ASAP7_75t_L g649 ( 
.A(n_275),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_47),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_642),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_13),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_141),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_605),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_36),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_339),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_264),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_83),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_126),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_508),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_632),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_608),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_215),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_277),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_2),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_434),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_464),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_622),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_250),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_481),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_149),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_445),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_301),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_621),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_200),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_8),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_598),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_114),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_145),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_595),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_587),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_502),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_152),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_201),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_516),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_454),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_620),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_24),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_495),
.Y(n_689)
);

BUFx8_ASAP7_75t_SL g690 ( 
.A(n_562),
.Y(n_690)
);

CKINVDCx16_ASAP7_75t_R g691 ( 
.A(n_374),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_414),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_581),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_507),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_424),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_169),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_38),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_136),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_145),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_247),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_306),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_557),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_619),
.Y(n_703)
);

CKINVDCx16_ASAP7_75t_R g704 ( 
.A(n_422),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_512),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_623),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_176),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_106),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_334),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_377),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_147),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_614),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_27),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_618),
.Y(n_714)
);

CKINVDCx14_ASAP7_75t_R g715 ( 
.A(n_637),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_574),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_212),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_348),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_440),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_38),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_70),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_584),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_303),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_283),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_44),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_158),
.Y(n_726)
);

BUFx5_ASAP7_75t_L g727 ( 
.A(n_636),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_350),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_553),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_184),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_251),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_398),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_504),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_626),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_247),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_374),
.Y(n_736)
);

BUFx10_ASAP7_75t_L g737 ( 
.A(n_19),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_514),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_578),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_256),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_182),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_612),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_285),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_197),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_336),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_560),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_18),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_21),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_242),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_326),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_163),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_396),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_146),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_339),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_236),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_268),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_213),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_299),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_191),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_550),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_341),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_417),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_400),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_68),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_342),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_159),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_68),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_424),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_289),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_360),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_468),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_634),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_99),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_380),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_21),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_40),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_428),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_83),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_506),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_52),
.Y(n_780)
);

BUFx5_ASAP7_75t_L g781 ( 
.A(n_163),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_382),
.Y(n_782)
);

BUFx8_ASAP7_75t_SL g783 ( 
.A(n_51),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_453),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_521),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_546),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_303),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_162),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_67),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_395),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_178),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_2),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_596),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_485),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_84),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_209),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_531),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_324),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_453),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_326),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_50),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_153),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_600),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_106),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_104),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_299),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_455),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_402),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_489),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_79),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_97),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_532),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_476),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_444),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_624),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_458),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_349),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_180),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_358),
.Y(n_819)
);

BUFx8_ASAP7_75t_SL g820 ( 
.A(n_607),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_402),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_178),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_419),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_35),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_602),
.Y(n_825)
);

BUFx5_ASAP7_75t_L g826 ( 
.A(n_57),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_546),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_597),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_60),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_205),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_234),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_17),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_82),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_118),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_237),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_523),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_370),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_470),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_67),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_27),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_207),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_525),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_287),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_628),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_209),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_350),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_641),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_584),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_134),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_29),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_355),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_556),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_304),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_79),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_245),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_551),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_454),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_195),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_558),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_418),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_65),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_52),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_358),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_313),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_39),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_171),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_575),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_261),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_507),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_610),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_129),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_344),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_429),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_49),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_379),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_544),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_129),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_544),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_367),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_445),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_57),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_164),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_530),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_520),
.Y(n_884)
);

CKINVDCx14_ASAP7_75t_R g885 ( 
.A(n_630),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_354),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_329),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_498),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_601),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_604),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_150),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_569),
.Y(n_892)
);

CKINVDCx16_ASAP7_75t_R g893 ( 
.A(n_141),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_347),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_211),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_469),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_633),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_120),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_81),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_640),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_310),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_310),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_435),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_548),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_115),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_320),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_594),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_609),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_311),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_214),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_229),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_513),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_428),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_189),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_112),
.Y(n_915)
);

BUFx10_ASAP7_75t_L g916 ( 
.A(n_629),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_627),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_287),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_561),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_193),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_139),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_499),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_440),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_353),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_395),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_295),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_301),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_223),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_631),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_184),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_530),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_244),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_384),
.Y(n_933)
);

BUFx10_ASAP7_75t_L g934 ( 
.A(n_545),
.Y(n_934)
);

BUFx5_ASAP7_75t_L g935 ( 
.A(n_499),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_536),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_41),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_420),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_313),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_217),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_72),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_140),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_309),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_324),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_112),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_386),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_414),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_423),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_598),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_503),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_528),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_421),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_244),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_603),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_464),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_635),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_0),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_317),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_297),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_314),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_69),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_280),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_164),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_251),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_496),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_89),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_114),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_245),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_77),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_12),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_615),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_166),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_383),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_439),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_566),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_199),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_321),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_393),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_262),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_462),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_240),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_54),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_435),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_268),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_220),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_561),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_433),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_34),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_406),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_535),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_625),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_195),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_97),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_147),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_364),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_446),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_393),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_512),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_505),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_429),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_582),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_564),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_176),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_590),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_348),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_576),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_220),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_547),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_617),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_416),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_154),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_319),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_365),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_300),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_457),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_248),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_186),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_100),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_277),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_256),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_154),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_377),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_386),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_613),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_179),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_250),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_7),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_531),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_144),
.Y(n_1029)
);

BUFx10_ASAP7_75t_L g1030 ( 
.A(n_280),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_237),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_567),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_616),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_390),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_33),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_372),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_152),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_143),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_8),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_433),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_375),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_36),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_290),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_541),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_104),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_46),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_611),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_119),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_86),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_130),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_50),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_33),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_594),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_192),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_215),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_585),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_113),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_518),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_218),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_476),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_172),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_599),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_297),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_214),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_314),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_596),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_536),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_457),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_538),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_228),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_368),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_177),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_532),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_638),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_170),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_579),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_497),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_602),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_425),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_347),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_426),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_514),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_182),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_504),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_406),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_203),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_380),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_533),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_199),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_572),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_88),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_248),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_208),
.Y(n_1093)
);

BUFx10_ASAP7_75t_L g1094 ( 
.A(n_566),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_603),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_81),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_45),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_559),
.Y(n_1098)
);

BUFx5_ASAP7_75t_L g1099 ( 
.A(n_5),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_146),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_4),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_42),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_66),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_31),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_349),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_87),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_196),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_325),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_444),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_576),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_606),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_330),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_413),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_135),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_473),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_161),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_53),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_639),
.Y(n_1118)
);

BUFx10_ASAP7_75t_L g1119 ( 
.A(n_322),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_24),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_96),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_371),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_31),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_241),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_551),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_353),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_385),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_217),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_469),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_235),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_405),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_7),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_524),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_131),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_107),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_961),
.Y(n_1136)
);

INVxp67_ASAP7_75t_SL g1137 ( 
.A(n_961),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_690),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_703),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_783),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_916),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_961),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_916),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_916),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_683),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_961),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_781),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_651),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_683),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_998),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_781),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_917),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_916),
.Y(n_1153)
);

INVxp33_ASAP7_75t_SL g1154 ( 
.A(n_886),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_998),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_691),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_998),
.Y(n_1157)
);

CKINVDCx16_ASAP7_75t_R g1158 ( 
.A(n_691),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_704),
.Y(n_1159)
);

INVxp67_ASAP7_75t_L g1160 ( 
.A(n_787),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1069),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1069),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_704),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1069),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_718),
.Y(n_1165)
);

INVxp33_ASAP7_75t_L g1166 ( 
.A(n_1104),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_787),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_718),
.Y(n_1168)
);

CKINVDCx16_ASAP7_75t_R g1169 ( 
.A(n_747),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_797),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_747),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_733),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_688),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_733),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_773),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_893),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_781),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_773),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_861),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_861),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_797),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_893),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_820),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_945),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_945),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_949),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_949),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1019),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1019),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_871),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_715),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_781),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_L g1193 ( 
.A(n_677),
.B(n_0),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_720),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_885),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_644),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_871),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_877),
.Y(n_1198)
);

INVxp67_ASAP7_75t_SL g1199 ( 
.A(n_652),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_735),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_877),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_923),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_923),
.Y(n_1203)
);

INVxp33_ASAP7_75t_SL g1204 ( 
.A(n_1107),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_946),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_946),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_645),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_646),
.Y(n_1208)
);

CKINVDCx16_ASAP7_75t_R g1209 ( 
.A(n_649),
.Y(n_1209)
);

INVxp33_ASAP7_75t_SL g1210 ( 
.A(n_1012),
.Y(n_1210)
);

CKINVDCx16_ASAP7_75t_R g1211 ( 
.A(n_649),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_781),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_648),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_781),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_781),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_781),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_781),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1012),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_752),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1018),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_826),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_826),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_826),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_826),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1018),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_650),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_653),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_826),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_656),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_657),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_826),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_826),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_826),
.Y(n_1233)
);

NOR2xp67_ASAP7_75t_L g1234 ( 
.A(n_677),
.B(n_738),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_763),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_658),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_826),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_935),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_647),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_817),
.Y(n_1240)
);

NOR2xp67_ASAP7_75t_L g1241 ( 
.A(n_738),
.B(n_1),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_647),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_935),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_935),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_659),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_660),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_935),
.Y(n_1247)
);

BUFx5_ASAP7_75t_L g1248 ( 
.A(n_662),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_935),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_666),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_935),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_669),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_671),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_935),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_935),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_676),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_655),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_655),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_665),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_678),
.Y(n_1260)
);

INVxp33_ASAP7_75t_L g1261 ( 
.A(n_665),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_649),
.B(n_664),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_935),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_681),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_667),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_667),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_652),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_672),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_822),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_703),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_662),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_649),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_672),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_682),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_673),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_824),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_830),
.Y(n_1277)
);

CKINVDCx14_ASAP7_75t_R g1278 ( 
.A(n_664),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_673),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1099),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_679),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_679),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_684),
.Y(n_1283)
);

INVxp33_ASAP7_75t_L g1284 ( 
.A(n_684),
.Y(n_1284)
);

CKINVDCx16_ASAP7_75t_R g1285 ( 
.A(n_664),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_692),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_692),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_694),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_694),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_687),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_L g1291 ( 
.A(n_762),
.B(n_775),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1099),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_696),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_696),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_685),
.Y(n_1295)
);

INVxp33_ASAP7_75t_SL g1296 ( 
.A(n_686),
.Y(n_1296)
);

CKINVDCx14_ASAP7_75t_R g1297 ( 
.A(n_664),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_668),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_699),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_689),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_699),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_695),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1099),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_668),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_700),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_700),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_701),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_701),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_702),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1099),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_698),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_702),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_705),
.Y(n_1313)
);

INVxp67_ASAP7_75t_SL g1314 ( 
.A(n_652),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_687),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_705),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_710),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_841),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_713),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_707),
.Y(n_1320)
);

INVxp33_ASAP7_75t_SL g1321 ( 
.A(n_719),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_846),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_707),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_721),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_709),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_722),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_709),
.Y(n_1327)
);

INVxp33_ASAP7_75t_L g1328 ( 
.A(n_716),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_716),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1099),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_717),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_717),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_725),
.Y(n_1333)
);

INVxp33_ASAP7_75t_L g1334 ( 
.A(n_725),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_754),
.Y(n_1335)
);

BUFx2_ASAP7_75t_SL g1336 ( 
.A(n_742),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_754),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_723),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_757),
.Y(n_1339)
);

INVx4_ASAP7_75t_R g1340 ( 
.A(n_742),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_757),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_768),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_848),
.Y(n_1343)
);

CKINVDCx14_ASAP7_75t_R g1344 ( 
.A(n_670),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_726),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_728),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_729),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_768),
.Y(n_1348)
);

INVxp33_ASAP7_75t_L g1349 ( 
.A(n_776),
.Y(n_1349)
);

CKINVDCx16_ASAP7_75t_R g1350 ( 
.A(n_670),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1099),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_776),
.Y(n_1352)
);

INVxp67_ASAP7_75t_SL g1353 ( 
.A(n_652),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_777),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_777),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_778),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_778),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_782),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_730),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_782),
.Y(n_1360)
);

XNOR2x1_ASAP7_75t_L g1361 ( 
.A(n_1135),
.B(n_680),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1134),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_789),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1099),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_852),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_731),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_668),
.Y(n_1367)
);

INVxp67_ASAP7_75t_SL g1368 ( 
.A(n_652),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_652),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_789),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1134),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1099),
.Y(n_1372)
);

INVxp33_ASAP7_75t_L g1373 ( 
.A(n_791),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_791),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1133),
.Y(n_1375)
);

INVxp67_ASAP7_75t_SL g1376 ( 
.A(n_663),
.Y(n_1376)
);

INVxp67_ASAP7_75t_SL g1377 ( 
.A(n_663),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_732),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_792),
.Y(n_1379)
);

INVx4_ASAP7_75t_R g1380 ( 
.A(n_870),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_736),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_792),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1133),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_796),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_796),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1132),
.Y(n_1386)
);

INVxp67_ASAP7_75t_SL g1387 ( 
.A(n_663),
.Y(n_1387)
);

NOR2xp67_ASAP7_75t_L g1388 ( 
.A(n_762),
.B(n_1),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_798),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_798),
.Y(n_1390)
);

INVxp33_ASAP7_75t_SL g1391 ( 
.A(n_739),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_801),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_668),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_801),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_853),
.Y(n_1395)
);

CKINVDCx14_ASAP7_75t_R g1396 ( 
.A(n_670),
.Y(n_1396)
);

CKINVDCx16_ASAP7_75t_R g1397 ( 
.A(n_670),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1132),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1099),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1131),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_740),
.Y(n_1401)
);

INVxp33_ASAP7_75t_L g1402 ( 
.A(n_803),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_803),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_860),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_805),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_873),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_663),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_741),
.Y(n_1408)
);

INVxp67_ASAP7_75t_SL g1409 ( 
.A(n_663),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_805),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1131),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_807),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_734),
.Y(n_1413)
);

INVxp67_ASAP7_75t_SL g1414 ( 
.A(n_663),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_813),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_807),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_808),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_813),
.Y(n_1418)
);

CKINVDCx16_ASAP7_75t_R g1419 ( 
.A(n_708),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_668),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_813),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_813),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_808),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_814),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_743),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_744),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_814),
.Y(n_1427)
);

INVxp33_ASAP7_75t_SL g1428 ( 
.A(n_745),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_746),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_775),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_748),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_819),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_819),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_823),
.Y(n_1434)
);

INVxp33_ASAP7_75t_SL g1435 ( 
.A(n_749),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_823),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_750),
.Y(n_1437)
);

NOR2xp67_ASAP7_75t_L g1438 ( 
.A(n_804),
.B(n_849),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_825),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_876),
.Y(n_1440)
);

CKINVDCx16_ASAP7_75t_R g1441 ( 
.A(n_708),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_751),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_753),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_825),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_755),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_829),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_804),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_829),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_833),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_833),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_813),
.Y(n_1451)
);

CKINVDCx14_ASAP7_75t_R g1452 ( 
.A(n_708),
.Y(n_1452)
);

CKINVDCx16_ASAP7_75t_R g1453 ( 
.A(n_708),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_835),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_756),
.Y(n_1455)
);

CKINVDCx14_ASAP7_75t_R g1456 ( 
.A(n_737),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_835),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_836),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_813),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_758),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_828),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_836),
.Y(n_1462)
);

INVxp67_ASAP7_75t_SL g1463 ( 
.A(n_828),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_759),
.Y(n_1464)
);

CKINVDCx16_ASAP7_75t_R g1465 ( 
.A(n_737),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_839),
.Y(n_1466)
);

CKINVDCx14_ASAP7_75t_R g1467 ( 
.A(n_737),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_849),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_839),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_895),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_840),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_760),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_828),
.Y(n_1473)
);

INVxp33_ASAP7_75t_SL g1474 ( 
.A(n_761),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_904),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_764),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_765),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_840),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_828),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_843),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_828),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_766),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_828),
.Y(n_1483)
);

INVxp67_ASAP7_75t_SL g1484 ( 
.A(n_868),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_767),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_843),
.Y(n_1486)
);

CKINVDCx20_ASAP7_75t_R g1487 ( 
.A(n_964),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_845),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_771),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_845),
.Y(n_1490)
);

INVxp33_ASAP7_75t_SL g1491 ( 
.A(n_774),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_851),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_851),
.Y(n_1493)
);

INVxp67_ASAP7_75t_SL g1494 ( 
.A(n_868),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_854),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_854),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_857),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_780),
.Y(n_1498)
);

INVxp33_ASAP7_75t_L g1499 ( 
.A(n_857),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_863),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_868),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_868),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_863),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_865),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_865),
.Y(n_1505)
);

CKINVDCx16_ASAP7_75t_R g1506 ( 
.A(n_737),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_784),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_972),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_785),
.Y(n_1509)
);

INVxp33_ASAP7_75t_L g1510 ( 
.A(n_875),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_875),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_882),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_882),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_883),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_883),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_888),
.Y(n_1516)
);

INVxp33_ASAP7_75t_SL g1517 ( 
.A(n_786),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_888),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_788),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_734),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_1000),
.Y(n_1521)
);

CKINVDCx16_ASAP7_75t_R g1522 ( 
.A(n_779),
.Y(n_1522)
);

INVxp67_ASAP7_75t_SL g1523 ( 
.A(n_868),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_889),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_815),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_790),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_815),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_844),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_844),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_868),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1004),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_991),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_991),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1009),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1009),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_793),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1111),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1014),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_794),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1111),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1017),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_879),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_668),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_795),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1139),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1136),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1142),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1183),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1146),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1262),
.B(n_779),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1191),
.B(n_890),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1137),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1150),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1157),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1183),
.Y(n_1555)
);

INVxp33_ASAP7_75t_SL g1556 ( 
.A(n_1191),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1195),
.B(n_674),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1161),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1162),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1148),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1164),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1152),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1138),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1138),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1199),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_SL g1566 ( 
.A(n_1272),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1322),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1314),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1353),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1368),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1369),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1173),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1376),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1267),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1377),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1387),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1409),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1194),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1140),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1195),
.B(n_674),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1414),
.Y(n_1581)
);

CKINVDCx16_ASAP7_75t_R g1582 ( 
.A(n_1209),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1200),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1463),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1235),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1484),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1219),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1494),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1240),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1318),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1278),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1523),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1520),
.Y(n_1593)
);

CKINVDCx16_ASAP7_75t_R g1594 ( 
.A(n_1211),
.Y(n_1594)
);

CKINVDCx20_ASAP7_75t_R g1595 ( 
.A(n_1269),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1297),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1520),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1276),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1525),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1525),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1277),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1343),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1344),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1527),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1365),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_R g1606 ( 
.A(n_1396),
.B(n_654),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1452),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1456),
.Y(n_1608)
);

CKINVDCx20_ASAP7_75t_R g1609 ( 
.A(n_1395),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1267),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1404),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1527),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1528),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1528),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1529),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1508),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_1139),
.Y(n_1617)
);

INVxp67_ASAP7_75t_SL g1618 ( 
.A(n_1270),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1406),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1440),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1274),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_1470),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1521),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1475),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1529),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1487),
.Y(n_1626)
);

NOR2xp67_ASAP7_75t_L g1627 ( 
.A(n_1141),
.B(n_661),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1532),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1532),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1531),
.Y(n_1630)
);

CKINVDCx20_ASAP7_75t_R g1631 ( 
.A(n_1538),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1533),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1533),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1541),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1267),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1534),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1158),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1196),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1196),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1534),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1535),
.Y(n_1641)
);

INVxp33_ASAP7_75t_L g1642 ( 
.A(n_1361),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1535),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1537),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1207),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1207),
.Y(n_1646)
);

INVxp67_ASAP7_75t_L g1647 ( 
.A(n_1345),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1537),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1208),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1540),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1208),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1213),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1213),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1540),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1257),
.Y(n_1655)
);

NOR2xp67_ASAP7_75t_L g1656 ( 
.A(n_1141),
.B(n_706),
.Y(n_1656)
);

INVxp33_ASAP7_75t_L g1657 ( 
.A(n_1361),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1226),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1262),
.B(n_859),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1258),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1226),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1227),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1227),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1259),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1407),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1265),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1266),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1229),
.Y(n_1668)
);

NOR2xp67_ASAP7_75t_L g1669 ( 
.A(n_1143),
.B(n_712),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1229),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1230),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1268),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1407),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1415),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1336),
.B(n_897),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1169),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1230),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1467),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1270),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1273),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1156),
.Y(n_1681)
);

CKINVDCx16_ASAP7_75t_R g1682 ( 
.A(n_1285),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1275),
.Y(n_1683)
);

INVxp33_ASAP7_75t_SL g1684 ( 
.A(n_1143),
.Y(n_1684)
);

CKINVDCx20_ASAP7_75t_R g1685 ( 
.A(n_1350),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1279),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1397),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1236),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1281),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_1419),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1282),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1283),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1286),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1236),
.Y(n_1694)
);

CKINVDCx16_ASAP7_75t_R g1695 ( 
.A(n_1441),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1289),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1245),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1245),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1293),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1156),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1246),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1299),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1301),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1246),
.Y(n_1704)
);

CKINVDCx20_ASAP7_75t_R g1705 ( 
.A(n_1453),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1305),
.Y(n_1706)
);

CKINVDCx20_ASAP7_75t_R g1707 ( 
.A(n_1465),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1306),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1307),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1250),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1250),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1308),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1309),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1252),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1312),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_1506),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1522),
.Y(n_1717)
);

INVxp33_ASAP7_75t_L g1718 ( 
.A(n_1347),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1159),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1313),
.Y(n_1720)
);

INVxp67_ASAP7_75t_SL g1721 ( 
.A(n_1155),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1316),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1336),
.B(n_897),
.Y(n_1723)
);

CKINVDCx20_ASAP7_75t_R g1724 ( 
.A(n_1159),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1163),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1252),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1320),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1253),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1323),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1325),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1253),
.Y(n_1731)
);

CKINVDCx16_ASAP7_75t_R g1732 ( 
.A(n_1489),
.Y(n_1732)
);

INVxp67_ASAP7_75t_SL g1733 ( 
.A(n_1271),
.Y(n_1733)
);

NOR2xp67_ASAP7_75t_L g1734 ( 
.A(n_1144),
.B(n_714),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1327),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1144),
.B(n_1024),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1153),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1329),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1256),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1256),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_1163),
.Y(n_1741)
);

CKINVDCx20_ASAP7_75t_R g1742 ( 
.A(n_1171),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1331),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1332),
.Y(n_1744)
);

INVxp67_ASAP7_75t_SL g1745 ( 
.A(n_1271),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1260),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1153),
.B(n_1024),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_R g1748 ( 
.A(n_1260),
.B(n_772),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1333),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1264),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1264),
.Y(n_1751)
);

CKINVDCx20_ASAP7_75t_R g1752 ( 
.A(n_1171),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1295),
.Y(n_1753)
);

CKINVDCx20_ASAP7_75t_R g1754 ( 
.A(n_1176),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1335),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1337),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1339),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1341),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1295),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1342),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1300),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1348),
.Y(n_1762)
);

CKINVDCx20_ASAP7_75t_R g1763 ( 
.A(n_1176),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1300),
.Y(n_1764)
);

CKINVDCx20_ASAP7_75t_R g1765 ( 
.A(n_1182),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1352),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1302),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1355),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1356),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1302),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_1182),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1357),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1358),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1360),
.Y(n_1774)
);

CKINVDCx20_ASAP7_75t_R g1775 ( 
.A(n_1311),
.Y(n_1775)
);

CKINVDCx20_ASAP7_75t_R g1776 ( 
.A(n_1311),
.Y(n_1776)
);

NOR2xp67_ASAP7_75t_L g1777 ( 
.A(n_1272),
.B(n_1317),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_R g1778 ( 
.A(n_1317),
.B(n_847),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1362),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1370),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1371),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1374),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1375),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1379),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1382),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1296),
.B(n_1321),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1319),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_1319),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1383),
.Y(n_1789)
);

INVxp67_ASAP7_75t_SL g1790 ( 
.A(n_1290),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1384),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1296),
.B(n_1118),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1385),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_1324),
.Y(n_1794)
);

INVxp67_ASAP7_75t_L g1795 ( 
.A(n_1509),
.Y(n_1795)
);

INVxp67_ASAP7_75t_L g1796 ( 
.A(n_1526),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1386),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1389),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1390),
.Y(n_1799)
);

CKINVDCx20_ASAP7_75t_R g1800 ( 
.A(n_1324),
.Y(n_1800)
);

INVxp67_ASAP7_75t_SL g1801 ( 
.A(n_1290),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1536),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1392),
.Y(n_1803)
);

CKINVDCx20_ASAP7_75t_R g1804 ( 
.A(n_1326),
.Y(n_1804)
);

CKINVDCx20_ASAP7_75t_R g1805 ( 
.A(n_1326),
.Y(n_1805)
);

CKINVDCx20_ASAP7_75t_R g1806 ( 
.A(n_1338),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1394),
.Y(n_1807)
);

INVxp67_ASAP7_75t_L g1808 ( 
.A(n_1170),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1398),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1400),
.Y(n_1810)
);

INVxp33_ASAP7_75t_L g1811 ( 
.A(n_1166),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1403),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1321),
.B(n_1118),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1338),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1346),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1346),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1405),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1410),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1145),
.B(n_1125),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1411),
.Y(n_1820)
);

CKINVDCx20_ASAP7_75t_R g1821 ( 
.A(n_1359),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1248),
.B(n_900),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1359),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1412),
.Y(n_1824)
);

CKINVDCx20_ASAP7_75t_R g1825 ( 
.A(n_1366),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1416),
.Y(n_1826)
);

CKINVDCx20_ASAP7_75t_R g1827 ( 
.A(n_1366),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1378),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1378),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1381),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1417),
.Y(n_1831)
);

INVxp67_ASAP7_75t_SL g1832 ( 
.A(n_1315),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1381),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1423),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1315),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1220),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1401),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1424),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1401),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1408),
.Y(n_1840)
);

CKINVDCx20_ASAP7_75t_R g1841 ( 
.A(n_1408),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1427),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1432),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1544),
.Y(n_1844)
);

CKINVDCx20_ASAP7_75t_R g1845 ( 
.A(n_1425),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1425),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1145),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1426),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1248),
.B(n_908),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1433),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1434),
.Y(n_1851)
);

NOR2xp67_ASAP7_75t_L g1852 ( 
.A(n_1426),
.B(n_929),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1436),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1429),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1261),
.B(n_779),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1429),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1431),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1431),
.Y(n_1858)
);

INVxp67_ASAP7_75t_SL g1859 ( 
.A(n_1413),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1439),
.Y(n_1860)
);

CKINVDCx16_ASAP7_75t_R g1861 ( 
.A(n_1149),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1437),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1413),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1444),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1446),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1448),
.Y(n_1866)
);

NOR2xp67_ASAP7_75t_L g1867 ( 
.A(n_1437),
.B(n_956),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1212),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1449),
.Y(n_1869)
);

INVx1_ASAP7_75t_SL g1870 ( 
.A(n_1544),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1442),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1450),
.Y(n_1872)
);

INVxp33_ASAP7_75t_SL g1873 ( 
.A(n_1442),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1454),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1149),
.Y(n_1875)
);

CKINVDCx20_ASAP7_75t_R g1876 ( 
.A(n_1443),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1593),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1811),
.B(n_1443),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1597),
.Y(n_1879)
);

CKINVDCx20_ASAP7_75t_R g1880 ( 
.A(n_1572),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1550),
.B(n_1239),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1868),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1855),
.B(n_1445),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1574),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1679),
.B(n_1242),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1679),
.B(n_1287),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1792),
.A2(n_1210),
.B1(n_1204),
.B2(n_1154),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1777),
.B(n_1248),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1574),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1721),
.B(n_1552),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1610),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1610),
.Y(n_1892)
);

AND2x2_ASAP7_75t_R g1893 ( 
.A(n_1684),
.B(n_1876),
.Y(n_1893)
);

INVx2_ASAP7_75t_SL g1894 ( 
.A(n_1676),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1599),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1635),
.Y(n_1896)
);

BUFx6f_ASAP7_75t_L g1897 ( 
.A(n_1868),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1600),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1675),
.B(n_1248),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1861),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1733),
.B(n_1288),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1604),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1612),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1585),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1635),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1613),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1590),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1813),
.A2(n_1210),
.B1(n_1204),
.B2(n_1154),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1565),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1665),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1614),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1615),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1775),
.A2(n_1048),
.B1(n_1054),
.B2(n_1028),
.Y(n_1913)
);

CKINVDCx20_ASAP7_75t_R g1914 ( 
.A(n_1572),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1579),
.Y(n_1915)
);

OA21x2_ASAP7_75t_L g1916 ( 
.A1(n_1822),
.A2(n_1214),
.B(n_1212),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1578),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1786),
.A2(n_1428),
.B1(n_1435),
.B2(n_1391),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1723),
.B(n_1248),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1745),
.B(n_1248),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1568),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1569),
.B(n_1391),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1790),
.B(n_1248),
.Y(n_1923)
);

BUFx6f_ASAP7_75t_L g1924 ( 
.A(n_1570),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1801),
.B(n_1248),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1625),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1665),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1571),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1718),
.B(n_1847),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1628),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1673),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1875),
.B(n_1445),
.Y(n_1932)
);

BUFx6f_ASAP7_75t_L g1933 ( 
.A(n_1573),
.Y(n_1933)
);

CKINVDCx20_ASAP7_75t_R g1934 ( 
.A(n_1578),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1736),
.A2(n_1435),
.B1(n_1474),
.B2(n_1428),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1629),
.Y(n_1936)
);

OAI21x1_ASAP7_75t_L g1937 ( 
.A1(n_1849),
.A2(n_1151),
.B(n_1147),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1673),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1546),
.Y(n_1939)
);

NAND2xp33_ASAP7_75t_R g1940 ( 
.A(n_1848),
.B(n_1474),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1844),
.B(n_1455),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1548),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1832),
.B(n_1294),
.Y(n_1943)
);

CKINVDCx20_ASAP7_75t_R g1944 ( 
.A(n_1583),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1674),
.Y(n_1945)
);

AND2x2_ASAP7_75t_SL g1946 ( 
.A(n_1582),
.B(n_693),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1674),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1632),
.Y(n_1948)
);

INVxp33_ASAP7_75t_SL g1949 ( 
.A(n_1737),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1633),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1636),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1747),
.B(n_1491),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1640),
.Y(n_1953)
);

INVxp67_ASAP7_75t_L g1954 ( 
.A(n_1611),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1641),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1575),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1576),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1577),
.Y(n_1958)
);

OAI22xp5_ASAP7_75t_SL g1959 ( 
.A1(n_1775),
.A2(n_1060),
.B1(n_1108),
.B2(n_1056),
.Y(n_1959)
);

AOI22x1_ASAP7_75t_SL g1960 ( 
.A1(n_1567),
.A2(n_1113),
.B1(n_800),
.B2(n_802),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1555),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1643),
.Y(n_1962)
);

INVx3_ASAP7_75t_L g1963 ( 
.A(n_1547),
.Y(n_1963)
);

INVx5_ASAP7_75t_L g1964 ( 
.A(n_1659),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1644),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1648),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1650),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1581),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1560),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1654),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1549),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1835),
.B(n_1455),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1584),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1870),
.B(n_1460),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1748),
.B(n_1778),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1859),
.B(n_1524),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1586),
.Y(n_1977)
);

XNOR2xp5_ASAP7_75t_L g1978 ( 
.A(n_1583),
.B(n_1460),
.Y(n_1978)
);

AOI22x1_ASAP7_75t_SL g1979 ( 
.A1(n_1587),
.A2(n_1589),
.B1(n_1598),
.B2(n_1595),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1863),
.B(n_1464),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1616),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1588),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1637),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1592),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1808),
.B(n_1464),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1553),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1655),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1554),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1836),
.B(n_1472),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1659),
.B(n_1354),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1659),
.B(n_1363),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1557),
.B(n_1472),
.Y(n_1992)
);

OA21x2_ASAP7_75t_L g1993 ( 
.A1(n_1558),
.A2(n_1215),
.B(n_1214),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1660),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1664),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1580),
.B(n_1476),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1559),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1545),
.B(n_1476),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1561),
.Y(n_1999)
);

CKINVDCx20_ASAP7_75t_R g2000 ( 
.A(n_1587),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1666),
.Y(n_2001)
);

INVxp67_ASAP7_75t_L g2002 ( 
.A(n_1623),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1621),
.B(n_1477),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1562),
.Y(n_2004)
);

BUFx6f_ASAP7_75t_L g2005 ( 
.A(n_1667),
.Y(n_2005)
);

INVx3_ASAP7_75t_L g2006 ( 
.A(n_1672),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1680),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1683),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1686),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1689),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1787),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_1732),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1624),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1626),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1630),
.Y(n_2015)
);

AND2x4_ASAP7_75t_L g2016 ( 
.A(n_1617),
.B(n_1234),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1618),
.B(n_1477),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1551),
.B(n_1482),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1634),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_SL g2020 ( 
.A1(n_1776),
.A2(n_1517),
.B1(n_1491),
.B2(n_1167),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1691),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1692),
.B(n_1291),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1693),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1696),
.B(n_1438),
.Y(n_2024)
);

CKINVDCx8_ASAP7_75t_R g2025 ( 
.A(n_1594),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1647),
.B(n_1482),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1699),
.Y(n_2027)
);

NAND2x1p5_ASAP7_75t_L g2028 ( 
.A(n_1702),
.B(n_1193),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1563),
.Y(n_2029)
);

BUFx2_ASAP7_75t_L g2030 ( 
.A(n_1637),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1627),
.B(n_1485),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1795),
.B(n_1485),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1656),
.B(n_1498),
.Y(n_2033)
);

INVx2_ASAP7_75t_SL g2034 ( 
.A(n_1591),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1564),
.Y(n_2035)
);

OAI22xp5_ASAP7_75t_SL g2036 ( 
.A1(n_1776),
.A2(n_1517),
.B1(n_1181),
.B2(n_1160),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1703),
.Y(n_2037)
);

OAI22xp5_ASAP7_75t_SL g2038 ( 
.A1(n_1788),
.A2(n_1507),
.B1(n_1498),
.B2(n_1519),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1706),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1708),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1709),
.Y(n_2041)
);

CKINVDCx6p67_ASAP7_75t_R g2042 ( 
.A(n_1788),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1591),
.Y(n_2043)
);

AND2x6_ASAP7_75t_L g2044 ( 
.A(n_1712),
.B(n_675),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_1713),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1715),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_1566),
.B(n_1507),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1720),
.Y(n_2048)
);

OAI22xp5_ASAP7_75t_SL g2049 ( 
.A1(n_1794),
.A2(n_1519),
.B1(n_1539),
.B2(n_1225),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_L g2050 ( 
.A(n_1566),
.B(n_1539),
.Y(n_2050)
);

BUFx6f_ASAP7_75t_L g2051 ( 
.A(n_1722),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1727),
.Y(n_2052)
);

AND2x6_ASAP7_75t_L g2053 ( 
.A(n_1729),
.B(n_675),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1730),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1735),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_1738),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1743),
.Y(n_2057)
);

NOR2xp67_ASAP7_75t_L g2058 ( 
.A(n_1596),
.B(n_1165),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1669),
.B(n_1430),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1744),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1749),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1566),
.B(n_1168),
.Y(n_2062)
);

INVx3_ASAP7_75t_L g2063 ( 
.A(n_1755),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1796),
.B(n_1218),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1734),
.B(n_1430),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1596),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1852),
.B(n_1867),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_SL g2068 ( 
.A1(n_1794),
.A2(n_1804),
.B1(n_1805),
.B2(n_1800),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1756),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1757),
.B(n_1447),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1758),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1760),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1762),
.Y(n_2073)
);

INVx3_ASAP7_75t_L g2074 ( 
.A(n_1766),
.Y(n_2074)
);

BUFx8_ASAP7_75t_L g2075 ( 
.A(n_1819),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1768),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1769),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1772),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1773),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1774),
.B(n_1447),
.Y(n_2080)
);

BUFx6f_ASAP7_75t_L g2081 ( 
.A(n_1779),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1780),
.Y(n_2082)
);

OA21x2_ASAP7_75t_L g2083 ( 
.A1(n_1781),
.A2(n_1216),
.B(n_1215),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1782),
.B(n_1468),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1783),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1784),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1785),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1789),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1791),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_1793),
.B(n_1172),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1848),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_1797),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1603),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1798),
.Y(n_2094)
);

BUFx3_ASAP7_75t_L g2095 ( 
.A(n_1799),
.Y(n_2095)
);

CKINVDCx20_ASAP7_75t_R g2096 ( 
.A(n_1589),
.Y(n_2096)
);

NOR2xp67_ASAP7_75t_L g2097 ( 
.A(n_1603),
.B(n_1174),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1803),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1807),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1809),
.Y(n_2100)
);

BUFx6f_ASAP7_75t_L g2101 ( 
.A(n_1810),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1607),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1812),
.Y(n_2103)
);

BUFx2_ASAP7_75t_L g2104 ( 
.A(n_1719),
.Y(n_2104)
);

AOI22x1_ASAP7_75t_SL g2105 ( 
.A1(n_1595),
.A2(n_806),
.B1(n_809),
.B2(n_799),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1802),
.B(n_1218),
.Y(n_2106)
);

INVx3_ASAP7_75t_L g2107 ( 
.A(n_1817),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1818),
.Y(n_2108)
);

AND2x4_ASAP7_75t_L g2109 ( 
.A(n_1820),
.B(n_1241),
.Y(n_2109)
);

CKINVDCx20_ASAP7_75t_R g2110 ( 
.A(n_1598),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1824),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1826),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1684),
.B(n_879),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1831),
.Y(n_2114)
);

INVx2_ASAP7_75t_SL g2115 ( 
.A(n_1607),
.Y(n_2115)
);

OAI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_1737),
.A2(n_1388),
.B1(n_943),
.B2(n_643),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1834),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1838),
.Y(n_2118)
);

OAI22xp5_ASAP7_75t_SL g2119 ( 
.A1(n_1800),
.A2(n_1225),
.B1(n_1328),
.B2(n_1284),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1608),
.B(n_1334),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_1608),
.B(n_1349),
.Y(n_2121)
);

BUFx6f_ASAP7_75t_L g2122 ( 
.A(n_1842),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1843),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1850),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1851),
.Y(n_2125)
);

OAI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_1873),
.A2(n_837),
.B1(n_862),
.B2(n_812),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_1678),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1853),
.Y(n_2128)
);

BUFx6f_ASAP7_75t_L g2129 ( 
.A(n_1860),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_L g2130 ( 
.A(n_1864),
.B(n_1175),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1865),
.B(n_1468),
.Y(n_2131)
);

AND2x4_ASAP7_75t_L g2132 ( 
.A(n_1866),
.B(n_1513),
.Y(n_2132)
);

CKINVDCx20_ASAP7_75t_R g2133 ( 
.A(n_1601),
.Y(n_2133)
);

BUFx3_ASAP7_75t_L g2134 ( 
.A(n_1869),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1872),
.B(n_1216),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1678),
.Y(n_2136)
);

NAND3xp33_ASAP7_75t_L g2137 ( 
.A(n_1638),
.B(n_1645),
.C(n_1639),
.Y(n_2137)
);

INVxp67_ASAP7_75t_L g2138 ( 
.A(n_1681),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_1606),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1874),
.Y(n_2140)
);

AOI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_1873),
.A2(n_878),
.B1(n_930),
.B2(n_711),
.Y(n_2141)
);

BUFx2_ASAP7_75t_L g2142 ( 
.A(n_1719),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_SL g2143 ( 
.A(n_1682),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_1646),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_1649),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1815),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1857),
.Y(n_2147)
);

OAI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_1556),
.A2(n_850),
.B1(n_869),
.B2(n_818),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1700),
.Y(n_2149)
);

INVx5_ASAP7_75t_L g2150 ( 
.A(n_1695),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1651),
.B(n_1217),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1652),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1653),
.Y(n_2153)
);

AOI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_1854),
.A2(n_968),
.B1(n_1001),
.B2(n_952),
.Y(n_2154)
);

BUFx6f_ASAP7_75t_L g2155 ( 
.A(n_1658),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_1854),
.B(n_1373),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1661),
.B(n_1217),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_1662),
.Y(n_2158)
);

AOI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_1856),
.A2(n_1042),
.B1(n_1072),
.B2(n_1040),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1663),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1668),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1670),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1671),
.B(n_1221),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_1677),
.B(n_1221),
.Y(n_2164)
);

INVxp67_ASAP7_75t_L g2165 ( 
.A(n_1856),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1688),
.Y(n_2166)
);

BUFx3_ASAP7_75t_L g2167 ( 
.A(n_1694),
.Y(n_2167)
);

BUFx6f_ASAP7_75t_L g2168 ( 
.A(n_1697),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1698),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1701),
.B(n_1222),
.Y(n_2170)
);

BUFx6f_ASAP7_75t_L g2171 ( 
.A(n_1704),
.Y(n_2171)
);

CKINVDCx20_ASAP7_75t_R g2172 ( 
.A(n_1601),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1710),
.Y(n_2173)
);

AND2x6_ASAP7_75t_L g2174 ( 
.A(n_1556),
.B(n_693),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1711),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1714),
.B(n_1222),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1726),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1728),
.B(n_1223),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1731),
.B(n_1223),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_1739),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1740),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_1746),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1750),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1751),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1858),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_1753),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_1759),
.B(n_879),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1761),
.B(n_1224),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_1858),
.B(n_1402),
.Y(n_2189)
);

INVx3_ASAP7_75t_L g2190 ( 
.A(n_1764),
.Y(n_2190)
);

CKINVDCx16_ASAP7_75t_R g2191 ( 
.A(n_1804),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1767),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1770),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1814),
.Y(n_2194)
);

CKINVDCx11_ASAP7_75t_R g2195 ( 
.A(n_1805),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_1862),
.B(n_1871),
.Y(n_2196)
);

OR2x2_ASAP7_75t_L g2197 ( 
.A(n_1862),
.B(n_1190),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1816),
.Y(n_2198)
);

BUFx6f_ASAP7_75t_L g2199 ( 
.A(n_1823),
.Y(n_2199)
);

HB1xp67_ASAP7_75t_L g2200 ( 
.A(n_1871),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_L g2201 ( 
.A(n_1828),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1829),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1830),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1833),
.Y(n_2204)
);

AOI22xp5_ASAP7_75t_L g2205 ( 
.A1(n_1837),
.A2(n_1109),
.B1(n_810),
.B2(n_821),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_1839),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1840),
.B(n_1224),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1806),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1806),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_1821),
.B(n_1503),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1821),
.Y(n_2211)
);

OAI22xp5_ASAP7_75t_SL g2212 ( 
.A1(n_1825),
.A2(n_1499),
.B1(n_1510),
.B2(n_864),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1825),
.Y(n_2213)
);

BUFx8_ASAP7_75t_L g2214 ( 
.A(n_1685),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1827),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1827),
.Y(n_2216)
);

INVx6_ASAP7_75t_L g2217 ( 
.A(n_1841),
.Y(n_2217)
);

BUFx6f_ASAP7_75t_L g2218 ( 
.A(n_1841),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_1642),
.B(n_1197),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1845),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1845),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1846),
.Y(n_2222)
);

BUFx6f_ASAP7_75t_L g2223 ( 
.A(n_1846),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1657),
.B(n_1228),
.Y(n_2224)
);

BUFx6f_ASAP7_75t_L g2225 ( 
.A(n_1876),
.Y(n_2225)
);

AND2x4_ASAP7_75t_L g2226 ( 
.A(n_1724),
.B(n_1511),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1724),
.Y(n_2227)
);

BUFx6f_ASAP7_75t_L g2228 ( 
.A(n_1685),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1725),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1725),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1687),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_1687),
.Y(n_2232)
);

OAI22xp5_ASAP7_75t_SL g2233 ( 
.A1(n_1602),
.A2(n_866),
.B1(n_887),
.B2(n_832),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_1690),
.B(n_1198),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_L g2235 ( 
.A(n_1690),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_1741),
.B(n_1518),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1705),
.B(n_1228),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1741),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1742),
.Y(n_2239)
);

AND2x2_ASAP7_75t_SL g2240 ( 
.A(n_1705),
.B(n_1007),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_1707),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_1742),
.B(n_879),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_1602),
.Y(n_2243)
);

BUFx3_ASAP7_75t_L g2244 ( 
.A(n_1707),
.Y(n_2244)
);

NAND2xp33_ASAP7_75t_L g2245 ( 
.A(n_1752),
.B(n_727),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1752),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_1754),
.B(n_1457),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1754),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_1716),
.Y(n_2249)
);

AND2x4_ASAP7_75t_L g2250 ( 
.A(n_1763),
.B(n_1458),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1763),
.Y(n_2251)
);

OA21x2_ASAP7_75t_L g2252 ( 
.A1(n_1765),
.A2(n_1232),
.B(n_1231),
.Y(n_2252)
);

BUFx2_ASAP7_75t_L g2253 ( 
.A(n_1765),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1771),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1716),
.B(n_1231),
.Y(n_2255)
);

XNOR2xp5_ASAP7_75t_L g2256 ( 
.A(n_1605),
.B(n_1380),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_1882),
.B(n_1232),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1910),
.Y(n_2258)
);

INVx4_ASAP7_75t_L g2259 ( 
.A(n_1882),
.Y(n_2259)
);

BUFx6f_ASAP7_75t_L g2260 ( 
.A(n_1882),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_2245),
.A2(n_1771),
.B1(n_1717),
.B2(n_975),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1909),
.Y(n_2262)
);

NAND2x1p5_ASAP7_75t_L g2263 ( 
.A(n_2083),
.B(n_1993),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_1910),
.Y(n_2264)
);

AOI22xp5_ASAP7_75t_L g2265 ( 
.A1(n_2245),
.A2(n_2174),
.B1(n_1922),
.B2(n_1952),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1909),
.Y(n_2266)
);

OAI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_2018),
.A2(n_827),
.B1(n_831),
.B2(n_816),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1909),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2156),
.B(n_2189),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1909),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1921),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1921),
.Y(n_2272)
);

HB1xp67_ASAP7_75t_L g2273 ( 
.A(n_1900),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_1927),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_1882),
.B(n_1233),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_L g2276 ( 
.A(n_1992),
.B(n_834),
.Y(n_2276)
);

BUFx2_ASAP7_75t_L g2277 ( 
.A(n_1900),
.Y(n_2277)
);

CKINVDCx5p33_ASAP7_75t_R g2278 ( 
.A(n_1904),
.Y(n_2278)
);

INVxp67_ASAP7_75t_L g2279 ( 
.A(n_1878),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1927),
.Y(n_2280)
);

INVx3_ASAP7_75t_L g2281 ( 
.A(n_1897),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1921),
.Y(n_2282)
);

INVx3_ASAP7_75t_L g2283 ( 
.A(n_1897),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1921),
.Y(n_2284)
);

INVx3_ASAP7_75t_L g2285 ( 
.A(n_1897),
.Y(n_2285)
);

OAI21x1_ASAP7_75t_L g2286 ( 
.A1(n_1937),
.A2(n_1151),
.B(n_1147),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1931),
.Y(n_2287)
);

AOI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2174),
.A2(n_1717),
.B1(n_975),
.B2(n_1015),
.Y(n_2288)
);

BUFx2_ASAP7_75t_L g2289 ( 
.A(n_2012),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1924),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1924),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_1897),
.B(n_1233),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_2005),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1924),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1924),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_2151),
.B(n_1237),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_2005),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_1931),
.Y(n_2298)
);

INVxp67_ASAP7_75t_L g2299 ( 
.A(n_1929),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1928),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1928),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1928),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2157),
.B(n_1237),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_1938),
.Y(n_2304)
);

AO22x1_ASAP7_75t_L g2305 ( 
.A1(n_2174),
.A2(n_2044),
.B1(n_2053),
.B2(n_1964),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1928),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1933),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1938),
.Y(n_2308)
);

BUFx2_ASAP7_75t_L g2309 ( 
.A(n_2012),
.Y(n_2309)
);

OAI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_1996),
.A2(n_842),
.B1(n_855),
.B2(n_838),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_1945),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1933),
.Y(n_2312)
);

OAI22xp5_ASAP7_75t_SL g2313 ( 
.A1(n_1913),
.A2(n_1609),
.B1(n_1619),
.B2(n_1605),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1933),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2163),
.B(n_1238),
.Y(n_2315)
);

INVx3_ASAP7_75t_L g2316 ( 
.A(n_1993),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2164),
.B(n_1238),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_2005),
.Y(n_2318)
);

CKINVDCx8_ASAP7_75t_R g2319 ( 
.A(n_2150),
.Y(n_2319)
);

INVx1_ASAP7_75t_SL g2320 ( 
.A(n_1907),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_1945),
.Y(n_2321)
);

AOI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2174),
.A2(n_1015),
.B1(n_1053),
.B2(n_859),
.Y(n_2322)
);

INVx1_ASAP7_75t_SL g2323 ( 
.A(n_1981),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_1947),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1933),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1956),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_1947),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1956),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1956),
.Y(n_2329)
);

BUFx6f_ASAP7_75t_L g2330 ( 
.A(n_2005),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_1884),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1956),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1957),
.Y(n_2333)
);

INVx3_ASAP7_75t_L g2334 ( 
.A(n_1993),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1884),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_1964),
.B(n_1462),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_1957),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_1889),
.Y(n_2338)
);

HB1xp67_ASAP7_75t_L g2339 ( 
.A(n_2243),
.Y(n_2339)
);

INVx3_ASAP7_75t_L g2340 ( 
.A(n_1986),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_1957),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_1890),
.B(n_1053),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1957),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1958),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1890),
.B(n_1088),
.Y(n_2345)
);

BUFx3_ASAP7_75t_L g2346 ( 
.A(n_2150),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_1958),
.Y(n_2347)
);

INVx3_ASAP7_75t_L g2348 ( 
.A(n_1986),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1958),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2170),
.B(n_1088),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1958),
.Y(n_2351)
);

CKINVDCx5p33_ASAP7_75t_R g2352 ( 
.A(n_1942),
.Y(n_2352)
);

NAND3xp33_ASAP7_75t_L g2353 ( 
.A(n_1887),
.B(n_1202),
.C(n_1201),
.Y(n_2353)
);

BUFx3_ASAP7_75t_L g2354 ( 
.A(n_2150),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1889),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1968),
.Y(n_2356)
);

INVxp67_ASAP7_75t_L g2357 ( 
.A(n_2120),
.Y(n_2357)
);

INVx3_ASAP7_75t_L g2358 ( 
.A(n_1986),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1968),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_1891),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1968),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2176),
.B(n_697),
.Y(n_2362)
);

OAI22xp5_ASAP7_75t_SL g2363 ( 
.A1(n_1959),
.A2(n_1619),
.B1(n_1620),
.B2(n_1609),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_1881),
.B(n_1178),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_SL g2365 ( 
.A(n_2025),
.B(n_1620),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_1968),
.Y(n_2366)
);

HB1xp67_ASAP7_75t_L g2367 ( 
.A(n_2243),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1891),
.Y(n_2368)
);

HB1xp67_ASAP7_75t_L g2369 ( 
.A(n_1894),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2174),
.A2(n_1033),
.B1(n_1047),
.B2(n_971),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1984),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_1984),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2178),
.B(n_697),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_1892),
.Y(n_2374)
);

BUFx6f_ASAP7_75t_L g2375 ( 
.A(n_2039),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1984),
.Y(n_2376)
);

HB1xp67_ASAP7_75t_L g2377 ( 
.A(n_2210),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_1892),
.Y(n_2378)
);

HB1xp67_ASAP7_75t_L g2379 ( 
.A(n_2210),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2179),
.B(n_724),
.Y(n_2380)
);

AND2x4_ASAP7_75t_L g2381 ( 
.A(n_1964),
.B(n_1466),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_1896),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_1896),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2188),
.B(n_724),
.Y(n_2384)
);

BUFx6f_ASAP7_75t_L g2385 ( 
.A(n_2039),
.Y(n_2385)
);

NAND2xp33_ASAP7_75t_SL g2386 ( 
.A(n_2155),
.B(n_769),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_1905),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1984),
.Y(n_2388)
);

HB1xp67_ASAP7_75t_L g2389 ( 
.A(n_2210),
.Y(n_2389)
);

INVx3_ASAP7_75t_L g2390 ( 
.A(n_1986),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_1988),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2207),
.B(n_769),
.Y(n_2392)
);

BUFx6f_ASAP7_75t_L g2393 ( 
.A(n_2039),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_1881),
.B(n_1179),
.Y(n_2394)
);

INVxp67_ASAP7_75t_L g2395 ( 
.A(n_2121),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_1905),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_1881),
.B(n_1180),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2006),
.B(n_770),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2006),
.B(n_770),
.Y(n_2399)
);

AOI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_1922),
.A2(n_1074),
.B1(n_856),
.B2(n_867),
.Y(n_2400)
);

CKINVDCx8_ASAP7_75t_R g2401 ( 
.A(n_2150),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1973),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_1899),
.B(n_1919),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_1973),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_1952),
.A2(n_858),
.B1(n_874),
.B2(n_872),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2083),
.Y(n_2406)
);

INVx1_ASAP7_75t_SL g2407 ( 
.A(n_1880),
.Y(n_2407)
);

BUFx8_ASAP7_75t_L g2408 ( 
.A(n_2143),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2083),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_1951),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_1951),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1977),
.Y(n_2412)
);

BUFx2_ASAP7_75t_L g2413 ( 
.A(n_2226),
.Y(n_2413)
);

INVx3_ASAP7_75t_L g2414 ( 
.A(n_1988),
.Y(n_2414)
);

OAI22xp5_ASAP7_75t_SL g2415 ( 
.A1(n_2068),
.A2(n_1631),
.B1(n_1622),
.B2(n_1205),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_1964),
.B(n_1243),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_1988),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_1966),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_2226),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1977),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_1988),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_1982),
.Y(n_2422)
);

AND2x2_ASAP7_75t_SL g2423 ( 
.A(n_2240),
.B(n_811),
.Y(n_2423)
);

INVx1_ASAP7_75t_SL g2424 ( 
.A(n_1880),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_1982),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_1966),
.Y(n_2426)
);

BUFx6f_ASAP7_75t_L g2427 ( 
.A(n_2039),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_1967),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_1967),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_1970),
.Y(n_2430)
);

NAND2xp33_ASAP7_75t_L g2431 ( 
.A(n_2155),
.B(n_727),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2063),
.B(n_811),
.Y(n_2432)
);

OAI22xp5_ASAP7_75t_SL g2433 ( 
.A1(n_1914),
.A2(n_1631),
.B1(n_1622),
.B2(n_1206),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_1970),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_1990),
.B(n_1184),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_2155),
.B(n_1243),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_1997),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1997),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_1999),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_1990),
.B(n_1185),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_SL g2441 ( 
.A(n_2155),
.B(n_1249),
.Y(n_2441)
);

HB1xp67_ASAP7_75t_L g2442 ( 
.A(n_2226),
.Y(n_2442)
);

INVx3_ASAP7_75t_L g2443 ( 
.A(n_2045),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_1999),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2001),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2001),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2045),
.Y(n_2447)
);

AND2x6_ASAP7_75t_L g2448 ( 
.A(n_1990),
.B(n_954),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_1991),
.B(n_1186),
.Y(n_2449)
);

OAI22xp5_ASAP7_75t_L g2450 ( 
.A1(n_1908),
.A2(n_880),
.B1(n_884),
.B2(n_881),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2007),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_1971),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_1971),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2007),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2009),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2009),
.Y(n_2456)
);

XNOR2x2_ASAP7_75t_L g2457 ( 
.A(n_2242),
.B(n_1203),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2010),
.Y(n_2458)
);

INVx3_ASAP7_75t_L g2459 ( 
.A(n_2045),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2063),
.B(n_954),
.Y(n_2460)
);

NAND2xp33_ASAP7_75t_SL g2461 ( 
.A(n_2168),
.B(n_984),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2010),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2021),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2074),
.B(n_984),
.Y(n_2464)
);

BUFx8_ASAP7_75t_L g2465 ( 
.A(n_2143),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_L g2466 ( 
.A(n_2224),
.B(n_891),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2021),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2048),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2048),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2052),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2167),
.B(n_1469),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2052),
.Y(n_2472)
);

AOI22xp5_ASAP7_75t_L g2473 ( 
.A1(n_2113),
.A2(n_892),
.B1(n_898),
.B2(n_896),
.Y(n_2473)
);

HB1xp67_ASAP7_75t_L g2474 ( 
.A(n_2236),
.Y(n_2474)
);

CKINVDCx8_ASAP7_75t_R g2475 ( 
.A(n_2191),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2061),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2061),
.Y(n_2477)
);

OAI22xp33_ASAP7_75t_L g2478 ( 
.A1(n_1935),
.A2(n_1007),
.B1(n_1071),
.B2(n_993),
.Y(n_2478)
);

BUFx2_ASAP7_75t_L g2479 ( 
.A(n_2236),
.Y(n_2479)
);

INVxp67_ASAP7_75t_L g2480 ( 
.A(n_1941),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2072),
.Y(n_2481)
);

INVx1_ASAP7_75t_SL g2482 ( 
.A(n_1914),
.Y(n_2482)
);

NAND2xp33_ASAP7_75t_SL g2483 ( 
.A(n_2168),
.B(n_993),
.Y(n_2483)
);

BUFx6f_ASAP7_75t_SL g2484 ( 
.A(n_2167),
.Y(n_2484)
);

BUFx6f_ASAP7_75t_L g2485 ( 
.A(n_2045),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2168),
.B(n_1249),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2072),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2073),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2073),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2074),
.B(n_1071),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2076),
.Y(n_2491)
);

BUFx6f_ASAP7_75t_L g2492 ( 
.A(n_2051),
.Y(n_2492)
);

BUFx6f_ASAP7_75t_L g2493 ( 
.A(n_2051),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_SL g2494 ( 
.A(n_2168),
.B(n_1251),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2076),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_2182),
.B(n_1471),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2086),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2086),
.Y(n_2498)
);

INVx3_ASAP7_75t_L g2499 ( 
.A(n_2051),
.Y(n_2499)
);

NAND2xp33_ASAP7_75t_SL g2500 ( 
.A(n_2171),
.B(n_1081),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2087),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2087),
.Y(n_2502)
);

AND2x2_ASAP7_75t_L g2503 ( 
.A(n_1991),
.B(n_1187),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2088),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2088),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2094),
.Y(n_2506)
);

BUFx2_ASAP7_75t_L g2507 ( 
.A(n_2236),
.Y(n_2507)
);

NOR2x1_ASAP7_75t_L g2508 ( 
.A(n_1975),
.B(n_1188),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2094),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2098),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2098),
.Y(n_2511)
);

INVx3_ASAP7_75t_L g2512 ( 
.A(n_2051),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2099),
.Y(n_2513)
);

AOI22xp5_ASAP7_75t_L g2514 ( 
.A1(n_2113),
.A2(n_902),
.B1(n_903),
.B2(n_901),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2099),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2092),
.B(n_1081),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2112),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2112),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2114),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2182),
.B(n_2095),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2114),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2117),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2117),
.Y(n_2523)
);

BUFx6f_ASAP7_75t_L g2524 ( 
.A(n_2054),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_1991),
.B(n_1189),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2123),
.Y(n_2526)
);

AND2x2_ASAP7_75t_SL g2527 ( 
.A(n_2240),
.B(n_889),
.Y(n_2527)
);

INVx3_ASAP7_75t_L g2528 ( 
.A(n_2054),
.Y(n_2528)
);

AOI22xp5_ASAP7_75t_L g2529 ( 
.A1(n_1883),
.A2(n_906),
.B1(n_907),
.B2(n_905),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2123),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_1974),
.B(n_1478),
.Y(n_2531)
);

AOI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_1901),
.A2(n_910),
.B1(n_913),
.B2(n_909),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2124),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2124),
.Y(n_2534)
);

BUFx2_ASAP7_75t_L g2535 ( 
.A(n_2247),
.Y(n_2535)
);

HB1xp67_ASAP7_75t_L g2536 ( 
.A(n_2247),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2054),
.Y(n_2537)
);

INVxp67_ASAP7_75t_L g2538 ( 
.A(n_1985),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2054),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2056),
.Y(n_2540)
);

AND2x4_ASAP7_75t_L g2541 ( 
.A(n_2095),
.B(n_2134),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_1877),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_1879),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_1895),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_1898),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2092),
.B(n_894),
.Y(n_2546)
);

AOI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_1901),
.A2(n_915),
.B1(n_918),
.B2(n_914),
.Y(n_2547)
);

NOR2x1_ASAP7_75t_L g2548 ( 
.A(n_1975),
.B(n_1480),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2056),
.Y(n_2549)
);

AOI22xp5_ASAP7_75t_L g2550 ( 
.A1(n_1901),
.A2(n_920),
.B1(n_922),
.B2(n_919),
.Y(n_2550)
);

INVx3_ASAP7_75t_L g2551 ( 
.A(n_2056),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_1943),
.B(n_1486),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2056),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_1902),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2078),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_1903),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_1906),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_1911),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_1912),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2078),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2078),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_1943),
.B(n_1976),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_2171),
.B(n_2186),
.Y(n_2563)
);

BUFx6f_ASAP7_75t_L g2564 ( 
.A(n_2078),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_1926),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2247),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2081),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2081),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2081),
.Y(n_2569)
);

NAND2xp33_ASAP7_75t_L g2570 ( 
.A(n_2171),
.B(n_2186),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_SL g2571 ( 
.A(n_2171),
.B(n_1251),
.Y(n_2571)
);

AOI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_1943),
.A2(n_926),
.B1(n_927),
.B2(n_924),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2081),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2089),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_1930),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_SL g2576 ( 
.A(n_2186),
.B(n_1254),
.Y(n_2576)
);

CKINVDCx8_ASAP7_75t_R g2577 ( 
.A(n_1942),
.Y(n_2577)
);

HB1xp67_ASAP7_75t_L g2578 ( 
.A(n_2250),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2089),
.Y(n_2579)
);

BUFx6f_ASAP7_75t_L g2580 ( 
.A(n_2089),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_1936),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2089),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2101),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2186),
.B(n_1254),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_1948),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_L g2586 ( 
.A(n_2101),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2101),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_SL g2588 ( 
.A(n_2199),
.B(n_1255),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_1950),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_1953),
.Y(n_2590)
);

BUFx6f_ASAP7_75t_L g2591 ( 
.A(n_2101),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_1955),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2122),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2122),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2107),
.B(n_894),
.Y(n_2595)
);

AOI22xp5_ASAP7_75t_L g2596 ( 
.A1(n_1976),
.A2(n_931),
.B1(n_932),
.B2(n_928),
.Y(n_2596)
);

INVx3_ASAP7_75t_L g2597 ( 
.A(n_2122),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2199),
.B(n_1255),
.Y(n_2598)
);

BUFx3_ASAP7_75t_L g2599 ( 
.A(n_2199),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_2122),
.Y(n_2600)
);

BUFx2_ASAP7_75t_L g2601 ( 
.A(n_2250),
.Y(n_2601)
);

CKINVDCx8_ASAP7_75t_R g2602 ( 
.A(n_1961),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_1962),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_1965),
.Y(n_2604)
);

HB1xp67_ASAP7_75t_L g2605 ( 
.A(n_2250),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_1987),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_1994),
.Y(n_2607)
);

BUFx6f_ASAP7_75t_L g2608 ( 
.A(n_2129),
.Y(n_2608)
);

HB1xp67_ASAP7_75t_L g2609 ( 
.A(n_1978),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_1995),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_1961),
.Y(n_2611)
);

AND2x4_ASAP7_75t_L g2612 ( 
.A(n_2134),
.B(n_1488),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2008),
.Y(n_2613)
);

AND2x6_ASAP7_75t_L g2614 ( 
.A(n_1976),
.B(n_899),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2023),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2107),
.B(n_899),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2027),
.Y(n_2617)
);

INVx1_ASAP7_75t_SL g2618 ( 
.A(n_1917),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2037),
.Y(n_2619)
);

HB1xp67_ASAP7_75t_L g2620 ( 
.A(n_1969),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2040),
.Y(n_2621)
);

INVx1_ASAP7_75t_SL g2622 ( 
.A(n_1917),
.Y(n_2622)
);

BUFx8_ASAP7_75t_L g2623 ( 
.A(n_1983),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2041),
.Y(n_2624)
);

AOI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_2252),
.A2(n_936),
.B1(n_938),
.B2(n_933),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2129),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2046),
.Y(n_2627)
);

INVxp67_ASAP7_75t_L g2628 ( 
.A(n_1989),
.Y(n_2628)
);

INVx1_ASAP7_75t_SL g2629 ( 
.A(n_1934),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2055),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_1939),
.B(n_911),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2057),
.Y(n_2632)
);

AND2x2_ASAP7_75t_L g2633 ( 
.A(n_2064),
.B(n_1490),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2060),
.Y(n_2634)
);

HB1xp67_ASAP7_75t_L g2635 ( 
.A(n_1969),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2129),
.Y(n_2636)
);

BUFx6f_ASAP7_75t_L g2637 ( 
.A(n_2129),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2069),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_2199),
.B(n_727),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2140),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_2004),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2071),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2276),
.B(n_2047),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2562),
.B(n_2132),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2402),
.Y(n_2645)
);

INVx1_ASAP7_75t_SL g2646 ( 
.A(n_2289),
.Y(n_2646)
);

AND2x4_ASAP7_75t_L g2647 ( 
.A(n_2562),
.B(n_2132),
.Y(n_2647)
);

AO22x2_ASAP7_75t_L g2648 ( 
.A1(n_2527),
.A2(n_2242),
.B1(n_1979),
.B2(n_2230),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2331),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2276),
.B(n_2047),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2404),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2331),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2412),
.Y(n_2653)
);

BUFx6f_ASAP7_75t_L g2654 ( 
.A(n_2385),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_2265),
.B(n_2201),
.Y(n_2655)
);

BUFx3_ASAP7_75t_L g2656 ( 
.A(n_2408),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2335),
.Y(n_2657)
);

NAND2x1p5_ASAP7_75t_L g2658 ( 
.A(n_2346),
.B(n_2201),
.Y(n_2658)
);

NAND3xp33_ASAP7_75t_L g2659 ( 
.A(n_2278),
.B(n_2185),
.C(n_2180),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2531),
.B(n_2050),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2335),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2420),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2338),
.Y(n_2663)
);

CKINVDCx14_ASAP7_75t_R g2664 ( 
.A(n_2278),
.Y(n_2664)
);

AND2x6_ASAP7_75t_L g2665 ( 
.A(n_2385),
.B(n_2201),
.Y(n_2665)
);

OR2x6_ASAP7_75t_L g2666 ( 
.A(n_2413),
.B(n_2217),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2338),
.Y(n_2667)
);

BUFx6f_ASAP7_75t_SL g2668 ( 
.A(n_2527),
.Y(n_2668)
);

BUFx4f_ASAP7_75t_L g2669 ( 
.A(n_2289),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2422),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2355),
.Y(n_2671)
);

AOI22xp33_ASAP7_75t_SL g2672 ( 
.A1(n_2423),
.A2(n_2119),
.B1(n_1946),
.B2(n_2212),
.Y(n_2672)
);

NAND2x1p5_ASAP7_75t_L g2673 ( 
.A(n_2346),
.B(n_2201),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2355),
.Y(n_2674)
);

BUFx2_ASAP7_75t_L g2675 ( 
.A(n_2309),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2360),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2531),
.B(n_2050),
.Y(n_2677)
);

INVxp67_ASAP7_75t_SL g2678 ( 
.A(n_2385),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2466),
.B(n_2153),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2425),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2606),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2466),
.B(n_2153),
.Y(n_2682)
);

OR2x2_ASAP7_75t_L g2683 ( 
.A(n_2407),
.B(n_2424),
.Y(n_2683)
);

AOI22xp33_ASAP7_75t_L g2684 ( 
.A1(n_2423),
.A2(n_2252),
.B1(n_2053),
.B2(n_2044),
.Y(n_2684)
);

CKINVDCx5p33_ASAP7_75t_R g2685 ( 
.A(n_2352),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_2352),
.Y(n_2686)
);

AOI22xp33_ASAP7_75t_SL g2687 ( 
.A1(n_2614),
.A2(n_1946),
.B1(n_2049),
.B2(n_2075),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2607),
.Y(n_2688)
);

AOI22xp33_ASAP7_75t_L g2689 ( 
.A1(n_2614),
.A2(n_2252),
.B1(n_2053),
.B2(n_2044),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_2385),
.B(n_2203),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2360),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2610),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2269),
.B(n_2196),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2269),
.B(n_2106),
.Y(n_2694)
);

AOI22xp33_ASAP7_75t_L g2695 ( 
.A1(n_2614),
.A2(n_2053),
.B1(n_2044),
.B2(n_2140),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2613),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2615),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_L g2698 ( 
.A(n_2538),
.B(n_2628),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2617),
.Y(n_2699)
);

AND2x6_ASAP7_75t_L g2700 ( 
.A(n_2385),
.B(n_2203),
.Y(n_2700)
);

BUFx3_ASAP7_75t_L g2701 ( 
.A(n_2408),
.Y(n_2701)
);

CKINVDCx20_ASAP7_75t_R g2702 ( 
.A(n_2611),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_L g2703 ( 
.A(n_2480),
.B(n_2279),
.Y(n_2703)
);

INVx5_ASAP7_75t_L g2704 ( 
.A(n_2427),
.Y(n_2704)
);

OAI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2542),
.A2(n_1949),
.B1(n_2165),
.B2(n_2161),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2619),
.Y(n_2706)
);

HB1xp67_ASAP7_75t_L g2707 ( 
.A(n_2309),
.Y(n_2707)
);

INVx5_ASAP7_75t_L g2708 ( 
.A(n_2427),
.Y(n_2708)
);

AO21x2_ASAP7_75t_L g2709 ( 
.A1(n_2403),
.A2(n_2639),
.B(n_2286),
.Y(n_2709)
);

INVx3_ASAP7_75t_L g2710 ( 
.A(n_2259),
.Y(n_2710)
);

AND2x6_ASAP7_75t_L g2711 ( 
.A(n_2427),
.B(n_2203),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2621),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_2427),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2624),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_SL g2715 ( 
.A(n_2427),
.B(n_2203),
.Y(n_2715)
);

INVx1_ASAP7_75t_SL g2716 ( 
.A(n_2277),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2627),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_SL g2718 ( 
.A(n_2320),
.B(n_1915),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_2524),
.B(n_2206),
.Y(n_2719)
);

BUFx2_ASAP7_75t_L g2720 ( 
.A(n_2277),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2630),
.Y(n_2721)
);

NOR2xp33_ASAP7_75t_L g2722 ( 
.A(n_2357),
.B(n_1949),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2632),
.Y(n_2723)
);

AND3x1_ASAP7_75t_L g2724 ( 
.A(n_2365),
.B(n_2215),
.C(n_2208),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2552),
.B(n_2161),
.Y(n_2725)
);

INVx1_ASAP7_75t_SL g2726 ( 
.A(n_2482),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2634),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2638),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2642),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_SL g2730 ( 
.A(n_2323),
.B(n_1915),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2633),
.B(n_2091),
.Y(n_2731)
);

INVxp67_ASAP7_75t_SL g2732 ( 
.A(n_2524),
.Y(n_2732)
);

AND2x4_ASAP7_75t_L g2733 ( 
.A(n_2354),
.B(n_2132),
.Y(n_2733)
);

AND2x2_ASAP7_75t_L g2734 ( 
.A(n_2633),
.B(n_2091),
.Y(n_2734)
);

INVx3_ASAP7_75t_L g2735 ( 
.A(n_2259),
.Y(n_2735)
);

BUFx3_ASAP7_75t_L g2736 ( 
.A(n_2408),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2552),
.B(n_2200),
.Y(n_2737)
);

INVx4_ASAP7_75t_L g2738 ( 
.A(n_2354),
.Y(n_2738)
);

INVx4_ASAP7_75t_L g2739 ( 
.A(n_2484),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2543),
.Y(n_2740)
);

BUFx2_ASAP7_75t_L g2741 ( 
.A(n_2273),
.Y(n_2741)
);

INVx4_ASAP7_75t_L g2742 ( 
.A(n_2484),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_SL g2743 ( 
.A(n_2524),
.B(n_2206),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_2611),
.Y(n_2744)
);

INVx6_ASAP7_75t_L g2745 ( 
.A(n_2465),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2299),
.B(n_2200),
.Y(n_2746)
);

AND2x4_ASAP7_75t_L g2747 ( 
.A(n_2520),
.B(n_2206),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2413),
.B(n_2003),
.Y(n_2748)
);

OAI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_2544),
.A2(n_2183),
.B1(n_2184),
.B2(n_2181),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2479),
.B(n_2026),
.Y(n_2750)
);

BUFx6f_ASAP7_75t_L g2751 ( 
.A(n_2524),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2368),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_SL g2753 ( 
.A(n_2524),
.B(n_2206),
.Y(n_2753)
);

INVx2_ASAP7_75t_SL g2754 ( 
.A(n_2369),
.Y(n_2754)
);

BUFx3_ASAP7_75t_L g2755 ( 
.A(n_2465),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2545),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2479),
.B(n_2032),
.Y(n_2757)
);

INVx3_ASAP7_75t_L g2758 ( 
.A(n_2259),
.Y(n_2758)
);

INVx2_ASAP7_75t_SL g2759 ( 
.A(n_2520),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_L g2760 ( 
.A(n_2395),
.B(n_2237),
.Y(n_2760)
);

INVx3_ASAP7_75t_L g2761 ( 
.A(n_2564),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2554),
.Y(n_2762)
);

INVxp67_ASAP7_75t_L g2763 ( 
.A(n_2614),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2556),
.Y(n_2764)
);

CKINVDCx5p33_ASAP7_75t_R g2765 ( 
.A(n_2577),
.Y(n_2765)
);

AND2x6_ASAP7_75t_L g2766 ( 
.A(n_2564),
.B(n_2144),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_L g2767 ( 
.A(n_2261),
.B(n_2255),
.Y(n_2767)
);

INVx4_ASAP7_75t_L g2768 ( 
.A(n_2484),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2614),
.B(n_2181),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2368),
.Y(n_2770)
);

INVx4_ASAP7_75t_L g2771 ( 
.A(n_2520),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2557),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_SL g2773 ( 
.A(n_2564),
.B(n_2144),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2558),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2471),
.B(n_1972),
.Y(n_2775)
);

OR2x6_ASAP7_75t_L g2776 ( 
.A(n_2507),
.B(n_2217),
.Y(n_2776)
);

INVx1_ASAP7_75t_SL g2777 ( 
.A(n_2618),
.Y(n_2777)
);

INVx2_ASAP7_75t_SL g2778 ( 
.A(n_2623),
.Y(n_2778)
);

AOI22xp33_ASAP7_75t_L g2779 ( 
.A1(n_2614),
.A2(n_2053),
.B1(n_2044),
.B2(n_2140),
.Y(n_2779)
);

BUFx4_ASAP7_75t_L g2780 ( 
.A(n_2465),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2564),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2559),
.Y(n_2782)
);

NOR2xp33_ASAP7_75t_L g2783 ( 
.A(n_2471),
.B(n_1980),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2507),
.B(n_2185),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_2457),
.A2(n_2140),
.B1(n_2233),
.B2(n_2036),
.Y(n_2785)
);

HB1xp67_ASAP7_75t_L g2786 ( 
.A(n_2535),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2374),
.Y(n_2787)
);

OR2x6_ASAP7_75t_L g2788 ( 
.A(n_2535),
.B(n_2217),
.Y(n_2788)
);

INVx4_ASAP7_75t_L g2789 ( 
.A(n_2541),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2565),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2374),
.Y(n_2791)
);

NOR2xp33_ASAP7_75t_L g2792 ( 
.A(n_2471),
.B(n_2146),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2378),
.Y(n_2793)
);

INVx4_ASAP7_75t_SL g2794 ( 
.A(n_2448),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2378),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2382),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2612),
.B(n_2342),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2601),
.B(n_1932),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2496),
.B(n_2146),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2382),
.Y(n_2800)
);

INVx3_ASAP7_75t_L g2801 ( 
.A(n_2564),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2383),
.Y(n_2802)
);

BUFx8_ASAP7_75t_SL g2803 ( 
.A(n_2601),
.Y(n_2803)
);

INVx8_ASAP7_75t_L g2804 ( 
.A(n_2448),
.Y(n_2804)
);

INVx4_ASAP7_75t_L g2805 ( 
.A(n_2541),
.Y(n_2805)
);

NAND3xp33_ASAP7_75t_L g2806 ( 
.A(n_2400),
.B(n_2162),
.C(n_1940),
.Y(n_2806)
);

XOR2x2_ASAP7_75t_L g2807 ( 
.A(n_2313),
.B(n_2363),
.Y(n_2807)
);

HB1xp67_ASAP7_75t_L g2808 ( 
.A(n_2377),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2612),
.B(n_2183),
.Y(n_2809)
);

CKINVDCx5p33_ASAP7_75t_R g2810 ( 
.A(n_2577),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2575),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2364),
.B(n_1954),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2581),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2612),
.B(n_2184),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_R g2815 ( 
.A(n_2602),
.B(n_2029),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2585),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2345),
.B(n_2192),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_SL g2818 ( 
.A(n_2608),
.B(n_2145),
.Y(n_2818)
);

NAND3x1_ASAP7_75t_L g2819 ( 
.A(n_2288),
.B(n_2211),
.C(n_2209),
.Y(n_2819)
);

NOR2xp33_ASAP7_75t_L g2820 ( 
.A(n_2496),
.B(n_2192),
.Y(n_2820)
);

AND2x4_ASAP7_75t_L g2821 ( 
.A(n_2599),
.B(n_1885),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2589),
.Y(n_2822)
);

BUFx10_ASAP7_75t_L g2823 ( 
.A(n_2496),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2383),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_L g2825 ( 
.A(n_2379),
.B(n_2204),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2387),
.Y(n_2826)
);

INVx6_ASAP7_75t_L g2827 ( 
.A(n_2623),
.Y(n_2827)
);

BUFx6f_ASAP7_75t_L g2828 ( 
.A(n_2608),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_SL g2829 ( 
.A(n_2608),
.B(n_2293),
.Y(n_2829)
);

BUFx6f_ASAP7_75t_L g2830 ( 
.A(n_2608),
.Y(n_2830)
);

INVx4_ASAP7_75t_L g2831 ( 
.A(n_2541),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2387),
.Y(n_2832)
);

INVx4_ASAP7_75t_L g2833 ( 
.A(n_2599),
.Y(n_2833)
);

INVx2_ASAP7_75t_SL g2834 ( 
.A(n_2623),
.Y(n_2834)
);

BUFx3_ASAP7_75t_L g2835 ( 
.A(n_2319),
.Y(n_2835)
);

BUFx2_ASAP7_75t_L g2836 ( 
.A(n_2622),
.Y(n_2836)
);

AOI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2457),
.A2(n_2077),
.B1(n_2082),
.B2(n_2079),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2590),
.B(n_2204),
.Y(n_2838)
);

AOI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_2570),
.A2(n_1940),
.B1(n_2160),
.B2(n_2152),
.Y(n_2839)
);

OR2x6_ASAP7_75t_L g2840 ( 
.A(n_2415),
.B(n_2218),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2396),
.Y(n_2841)
);

NAND2x1p5_ASAP7_75t_L g2842 ( 
.A(n_2608),
.B(n_1939),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2364),
.B(n_2002),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2592),
.Y(n_2844)
);

INVx1_ASAP7_75t_SL g2845 ( 
.A(n_2629),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2603),
.Y(n_2846)
);

NAND2x1p5_ASAP7_75t_L g2847 ( 
.A(n_2293),
.B(n_1963),
.Y(n_2847)
);

AOI22xp33_ASAP7_75t_L g2848 ( 
.A1(n_2604),
.A2(n_2100),
.B1(n_2103),
.B2(n_2085),
.Y(n_2848)
);

BUFx2_ASAP7_75t_L g2849 ( 
.A(n_2339),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_SL g2850 ( 
.A(n_2293),
.B(n_2145),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2452),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2452),
.Y(n_2852)
);

INVx4_ASAP7_75t_L g2853 ( 
.A(n_2448),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2362),
.B(n_2158),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2453),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2453),
.Y(n_2856)
);

INVx3_ASAP7_75t_L g2857 ( 
.A(n_2293),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2373),
.B(n_2158),
.Y(n_2858)
);

NOR2xp33_ASAP7_75t_L g2859 ( 
.A(n_2389),
.B(n_1998),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_SL g2860 ( 
.A(n_2297),
.B(n_2318),
.Y(n_2860)
);

INVx3_ASAP7_75t_L g2861 ( 
.A(n_2297),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2396),
.Y(n_2862)
);

INVx4_ASAP7_75t_L g2863 ( 
.A(n_2448),
.Y(n_2863)
);

INVxp33_ASAP7_75t_SL g2864 ( 
.A(n_2620),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2454),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2380),
.B(n_2190),
.Y(n_2866)
);

INVx6_ASAP7_75t_L g2867 ( 
.A(n_2336),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2454),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2456),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2456),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2458),
.Y(n_2871)
);

AND2x2_ASAP7_75t_SL g2872 ( 
.A(n_2570),
.B(n_2431),
.Y(n_2872)
);

AND2x4_ASAP7_75t_L g2873 ( 
.A(n_2435),
.B(n_1885),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2458),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2462),
.Y(n_2875)
);

AND2x4_ASAP7_75t_L g2876 ( 
.A(n_2435),
.B(n_1885),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_SL g2877 ( 
.A(n_2297),
.B(n_2190),
.Y(n_2877)
);

NOR2xp33_ASAP7_75t_L g2878 ( 
.A(n_2419),
.B(n_2017),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2384),
.B(n_1886),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2392),
.B(n_1886),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_SL g2881 ( 
.A(n_2297),
.B(n_2318),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2462),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2467),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2258),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2258),
.Y(n_2885)
);

AND2x6_ASAP7_75t_L g2886 ( 
.A(n_2406),
.B(n_1886),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2467),
.Y(n_2887)
);

AOI22xp33_ASAP7_75t_L g2888 ( 
.A1(n_2448),
.A2(n_2111),
.B1(n_2118),
.B2(n_2108),
.Y(n_2888)
);

OR2x2_ASAP7_75t_L g2889 ( 
.A(n_2609),
.B(n_2104),
.Y(n_2889)
);

AND2x2_ASAP7_75t_L g2890 ( 
.A(n_2394),
.B(n_2219),
.Y(n_2890)
);

NAND2x1p5_ASAP7_75t_L g2891 ( 
.A(n_2318),
.B(n_1963),
.Y(n_2891)
);

INVxp67_ASAP7_75t_L g2892 ( 
.A(n_2394),
.Y(n_2892)
);

OAI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2350),
.A2(n_2011),
.B1(n_2169),
.B2(n_2166),
.Y(n_2893)
);

CKINVDCx5p33_ASAP7_75t_R g2894 ( 
.A(n_2602),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2336),
.B(n_2062),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2336),
.B(n_2062),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2264),
.Y(n_2897)
);

OR2x6_ASAP7_75t_L g2898 ( 
.A(n_2305),
.B(n_2218),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2381),
.B(n_2016),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2381),
.B(n_2016),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2264),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2397),
.B(n_2197),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2468),
.Y(n_2903)
);

BUFx6f_ASAP7_75t_SL g2904 ( 
.A(n_2448),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2274),
.Y(n_2905)
);

OR2x6_ASAP7_75t_L g2906 ( 
.A(n_2305),
.B(n_2218),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2468),
.Y(n_2907)
);

OR2x2_ASAP7_75t_L g2908 ( 
.A(n_2367),
.B(n_2142),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2501),
.Y(n_2909)
);

HB1xp67_ASAP7_75t_L g2910 ( 
.A(n_2442),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2381),
.B(n_2016),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2274),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2501),
.Y(n_2913)
);

BUFx3_ASAP7_75t_L g2914 ( 
.A(n_2319),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2397),
.B(n_2125),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2502),
.Y(n_2916)
);

NAND2xp33_ASAP7_75t_SL g2917 ( 
.A(n_2563),
.B(n_2029),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2502),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2440),
.B(n_2128),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2280),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2504),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2280),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2440),
.B(n_2090),
.Y(n_2923)
);

INVx5_ASAP7_75t_L g2924 ( 
.A(n_2318),
.Y(n_2924)
);

BUFx6f_ASAP7_75t_L g2925 ( 
.A(n_2260),
.Y(n_2925)
);

NAND3xp33_ASAP7_75t_L g2926 ( 
.A(n_2267),
.B(n_2035),
.C(n_2019),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_SL g2927 ( 
.A(n_2330),
.B(n_1920),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2504),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2287),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_SL g2930 ( 
.A(n_2475),
.B(n_2004),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2505),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2287),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_SL g2933 ( 
.A(n_2330),
.B(n_1923),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2449),
.B(n_2035),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2298),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2505),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2511),
.Y(n_2937)
);

AOI22xp5_ASAP7_75t_L g2938 ( 
.A1(n_2478),
.A2(n_2175),
.B1(n_2177),
.B2(n_2173),
.Y(n_2938)
);

BUFx2_ASAP7_75t_L g2939 ( 
.A(n_2635),
.Y(n_2939)
);

NAND3xp33_ASAP7_75t_L g2940 ( 
.A(n_2310),
.B(n_2019),
.C(n_2014),
.Y(n_2940)
);

CKINVDCx5p33_ASAP7_75t_R g2941 ( 
.A(n_2475),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2298),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2511),
.Y(n_2943)
);

INVx3_ASAP7_75t_L g2944 ( 
.A(n_2330),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2304),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2515),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2304),
.Y(n_2947)
);

BUFx3_ASAP7_75t_L g2948 ( 
.A(n_2401),
.Y(n_2948)
);

OAI21xp33_ASAP7_75t_L g2949 ( 
.A1(n_2405),
.A2(n_1918),
.B(n_2126),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2515),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2523),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2523),
.Y(n_2952)
);

AND2x2_ASAP7_75t_L g2953 ( 
.A(n_2449),
.B(n_2234),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2308),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2503),
.B(n_2090),
.Y(n_2955)
);

BUFx10_ASAP7_75t_L g2956 ( 
.A(n_2641),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2526),
.Y(n_2957)
);

OR2x2_ASAP7_75t_L g2958 ( 
.A(n_2474),
.B(n_2253),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2526),
.Y(n_2959)
);

AND2x4_ASAP7_75t_L g2960 ( 
.A(n_2503),
.B(n_2109),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2533),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2308),
.Y(n_2962)
);

OR2x6_ASAP7_75t_L g2963 ( 
.A(n_2433),
.B(n_2218),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2533),
.Y(n_2964)
);

NOR2xp33_ASAP7_75t_L g2965 ( 
.A(n_2536),
.B(n_2059),
.Y(n_2965)
);

BUFx4f_ASAP7_75t_L g2966 ( 
.A(n_2525),
.Y(n_2966)
);

OAI22xp5_ASAP7_75t_L g2967 ( 
.A1(n_2340),
.A2(n_2193),
.B1(n_2198),
.B2(n_2194),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2534),
.Y(n_2968)
);

CKINVDCx20_ASAP7_75t_R g2969 ( 
.A(n_2401),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_SL g2970 ( 
.A(n_2330),
.B(n_1925),
.Y(n_2970)
);

INVx2_ASAP7_75t_SL g2971 ( 
.A(n_2525),
.Y(n_2971)
);

OR2x6_ASAP7_75t_L g2972 ( 
.A(n_2566),
.B(n_2223),
.Y(n_2972)
);

NAND2xp33_ASAP7_75t_SL g2973 ( 
.A(n_2563),
.B(n_2139),
.Y(n_2973)
);

CKINVDCx20_ASAP7_75t_R g2974 ( 
.A(n_2578),
.Y(n_2974)
);

AND2x6_ASAP7_75t_L g2975 ( 
.A(n_2406),
.B(n_2202),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2311),
.Y(n_2976)
);

INVx5_ASAP7_75t_L g2977 ( 
.A(n_2375),
.Y(n_2977)
);

AND2x4_ASAP7_75t_L g2978 ( 
.A(n_2605),
.B(n_2109),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_2260),
.Y(n_2979)
);

BUFx3_ASAP7_75t_L g2980 ( 
.A(n_2260),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2375),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_L g2982 ( 
.A(n_2532),
.B(n_2065),
.Y(n_2982)
);

INVx4_ASAP7_75t_L g2983 ( 
.A(n_2375),
.Y(n_2983)
);

BUFx2_ASAP7_75t_L g2984 ( 
.A(n_2386),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2311),
.Y(n_2985)
);

NOR2xp33_ASAP7_75t_L g2986 ( 
.A(n_2547),
.B(n_2147),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2546),
.B(n_2130),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2321),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2321),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2534),
.Y(n_2990)
);

BUFx6f_ASAP7_75t_SL g2991 ( 
.A(n_2260),
.Y(n_2991)
);

INVx3_ASAP7_75t_L g2992 ( 
.A(n_2375),
.Y(n_2992)
);

INVx4_ASAP7_75t_L g2993 ( 
.A(n_2393),
.Y(n_2993)
);

OR2x2_ASAP7_75t_L g2994 ( 
.A(n_2353),
.B(n_2213),
.Y(n_2994)
);

BUFx3_ASAP7_75t_L g2995 ( 
.A(n_2393),
.Y(n_2995)
);

INVx3_ASAP7_75t_L g2996 ( 
.A(n_2393),
.Y(n_2996)
);

AND2x6_ASAP7_75t_L g2997 ( 
.A(n_2409),
.B(n_2109),
.Y(n_2997)
);

AOI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2322),
.A2(n_2137),
.B1(n_2187),
.B2(n_2020),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_2529),
.B(n_2215),
.Y(n_2999)
);

HB1xp67_ASAP7_75t_L g3000 ( 
.A(n_2393),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2550),
.B(n_2149),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2324),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2595),
.B(n_2130),
.Y(n_3003)
);

INVx4_ASAP7_75t_SL g3004 ( 
.A(n_2485),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2410),
.Y(n_3005)
);

BUFx8_ASAP7_75t_SL g3006 ( 
.A(n_2616),
.Y(n_3006)
);

INVxp67_ASAP7_75t_SL g3007 ( 
.A(n_2409),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2410),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2572),
.B(n_2031),
.Y(n_3009)
);

NOR2xp33_ASAP7_75t_SL g3010 ( 
.A(n_2548),
.B(n_2013),
.Y(n_3010)
);

AND2x6_ASAP7_75t_L g3011 ( 
.A(n_2485),
.B(n_2228),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2631),
.B(n_2028),
.Y(n_3012)
);

BUFx3_ASAP7_75t_L g3013 ( 
.A(n_2485),
.Y(n_3013)
);

AOI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2386),
.A2(n_2187),
.B1(n_2139),
.B2(n_2138),
.Y(n_3014)
);

OR2x2_ASAP7_75t_L g3015 ( 
.A(n_2450),
.B(n_2213),
.Y(n_3015)
);

NOR2xp33_ASAP7_75t_L g3016 ( 
.A(n_2596),
.B(n_2033),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2324),
.Y(n_3017)
);

BUFx6f_ASAP7_75t_L g3018 ( 
.A(n_2485),
.Y(n_3018)
);

CKINVDCx16_ASAP7_75t_R g3019 ( 
.A(n_2461),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2411),
.Y(n_3020)
);

INVx2_ASAP7_75t_SL g3021 ( 
.A(n_2508),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_SL g3022 ( 
.A(n_2492),
.B(n_1888),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2473),
.B(n_2208),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2411),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2327),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2418),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2418),
.Y(n_3027)
);

BUFx6f_ASAP7_75t_L g3028 ( 
.A(n_2492),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2649),
.Y(n_3029)
);

INVx2_ASAP7_75t_SL g3030 ( 
.A(n_2669),
.Y(n_3030)
);

NOR2xp33_ASAP7_75t_L g3031 ( 
.A(n_2643),
.B(n_2216),
.Y(n_3031)
);

NOR2xp33_ASAP7_75t_L g3032 ( 
.A(n_2650),
.B(n_2216),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2681),
.Y(n_3033)
);

NOR3xp33_ASAP7_75t_L g3034 ( 
.A(n_2949),
.B(n_2038),
.C(n_2220),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2649),
.Y(n_3035)
);

NAND2x1p5_ASAP7_75t_L g3036 ( 
.A(n_2853),
.B(n_2492),
.Y(n_3036)
);

BUFx6f_ASAP7_75t_SL g3037 ( 
.A(n_2656),
.Y(n_3037)
);

NOR2xp67_ASAP7_75t_L g3038 ( 
.A(n_2659),
.B(n_2015),
.Y(n_3038)
);

AOI22xp33_ASAP7_75t_L g3039 ( 
.A1(n_2672),
.A2(n_2426),
.B1(n_2625),
.B2(n_2438),
.Y(n_3039)
);

BUFx2_ASAP7_75t_L g3040 ( 
.A(n_2669),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2667),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2688),
.Y(n_3042)
);

OR2x2_ASAP7_75t_L g3043 ( 
.A(n_2646),
.B(n_2030),
.Y(n_3043)
);

NAND3xp33_ASAP7_75t_L g3044 ( 
.A(n_2982),
.B(n_2141),
.C(n_2221),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2667),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_SL g3046 ( 
.A(n_2966),
.B(n_2223),
.Y(n_3046)
);

NOR2xp33_ASAP7_75t_L g3047 ( 
.A(n_2660),
.B(n_2221),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2676),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_SL g3049 ( 
.A(n_2966),
.B(n_2722),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_SL g3050 ( 
.A(n_2722),
.B(n_2223),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2692),
.Y(n_3051)
);

BUFx6f_ASAP7_75t_L g3052 ( 
.A(n_2654),
.Y(n_3052)
);

NOR2xp67_ASAP7_75t_L g3053 ( 
.A(n_2765),
.B(n_2034),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2696),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2697),
.Y(n_3055)
);

HB1xp67_ASAP7_75t_L g3056 ( 
.A(n_2707),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2676),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2760),
.B(n_2767),
.Y(n_3058)
);

NOR2xp33_ASAP7_75t_L g3059 ( 
.A(n_2677),
.B(n_2227),
.Y(n_3059)
);

INVxp67_ASAP7_75t_L g3060 ( 
.A(n_2707),
.Y(n_3060)
);

INVx2_ASAP7_75t_SL g3061 ( 
.A(n_2827),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2718),
.B(n_2223),
.Y(n_3062)
);

NOR2x1p5_ASAP7_75t_L g3063 ( 
.A(n_2656),
.B(n_2042),
.Y(n_3063)
);

INVxp67_ASAP7_75t_SL g3064 ( 
.A(n_3007),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2699),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2760),
.B(n_2070),
.Y(n_3066)
);

AOI22xp5_ASAP7_75t_L g3067 ( 
.A1(n_2767),
.A2(n_2230),
.B1(n_2248),
.B2(n_2227),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2731),
.B(n_2080),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2734),
.B(n_2084),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2800),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2775),
.B(n_2131),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2706),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2775),
.B(n_2028),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_SL g3074 ( 
.A(n_2730),
.B(n_2225),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2800),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2934),
.B(n_2225),
.Y(n_3076)
);

NOR2xp33_ASAP7_75t_L g3077 ( 
.A(n_2679),
.B(n_2248),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2802),
.Y(n_3078)
);

INVx2_ASAP7_75t_SL g3079 ( 
.A(n_2827),
.Y(n_3079)
);

HB1xp67_ASAP7_75t_L g3080 ( 
.A(n_2786),
.Y(n_3080)
);

AOI22xp33_ASAP7_75t_L g3081 ( 
.A1(n_2672),
.A2(n_2426),
.B1(n_2439),
.B2(n_2437),
.Y(n_3081)
);

NOR2xp33_ASAP7_75t_L g3082 ( 
.A(n_2682),
.B(n_2222),
.Y(n_3082)
);

BUFx3_ASAP7_75t_L g3083 ( 
.A(n_2701),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2802),
.Y(n_3084)
);

OR2x2_ASAP7_75t_L g3085 ( 
.A(n_2716),
.B(n_2244),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2712),
.Y(n_3086)
);

INVx2_ASAP7_75t_L g3087 ( 
.A(n_2832),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2783),
.B(n_2444),
.Y(n_3088)
);

AOI22xp33_ASAP7_75t_L g3089 ( 
.A1(n_2648),
.A2(n_2446),
.B1(n_2451),
.B2(n_2445),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2783),
.B(n_2455),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2923),
.B(n_2463),
.Y(n_3091)
);

AOI22xp33_ASAP7_75t_L g3092 ( 
.A1(n_2648),
.A2(n_2470),
.B1(n_2472),
.B2(n_2469),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_SL g3093 ( 
.A(n_2784),
.B(n_2225),
.Y(n_3093)
);

INVx8_ASAP7_75t_L g3094 ( 
.A(n_3011),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_SL g3095 ( 
.A(n_2815),
.B(n_2930),
.Y(n_3095)
);

BUFx6f_ASAP7_75t_L g3096 ( 
.A(n_2835),
.Y(n_3096)
);

NOR2xp33_ASAP7_75t_L g3097 ( 
.A(n_2982),
.B(n_2644),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_2902),
.B(n_2225),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2955),
.B(n_2476),
.Y(n_3099)
);

AND2x2_ASAP7_75t_L g3100 ( 
.A(n_2953),
.B(n_2154),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2714),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2717),
.Y(n_3102)
);

NAND3xp33_ASAP7_75t_L g3103 ( 
.A(n_2785),
.B(n_3016),
.C(n_3009),
.Y(n_3103)
);

NOR2xp33_ASAP7_75t_SL g3104 ( 
.A(n_2685),
.B(n_1934),
.Y(n_3104)
);

AND2x4_ASAP7_75t_L g3105 ( 
.A(n_2644),
.B(n_2340),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2694),
.B(n_2477),
.Y(n_3106)
);

NAND2x1_ASAP7_75t_L g3107 ( 
.A(n_2665),
.B(n_2700),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_2832),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2721),
.Y(n_3109)
);

INVx4_ASAP7_75t_L g3110 ( 
.A(n_2991),
.Y(n_3110)
);

NOR2xp33_ASAP7_75t_L g3111 ( 
.A(n_2647),
.B(n_2229),
.Y(n_3111)
);

INVx2_ASAP7_75t_SL g3112 ( 
.A(n_2827),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2890),
.B(n_2481),
.Y(n_3113)
);

CKINVDCx20_ASAP7_75t_R g3114 ( 
.A(n_2702),
.Y(n_3114)
);

AND2x6_ASAP7_75t_SL g3115 ( 
.A(n_2963),
.B(n_2238),
.Y(n_3115)
);

INVx2_ASAP7_75t_SL g3116 ( 
.A(n_2745),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2723),
.Y(n_3117)
);

INVxp67_ASAP7_75t_L g3118 ( 
.A(n_2675),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2820),
.B(n_2487),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2820),
.B(n_2488),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2727),
.Y(n_3121)
);

INVx8_ASAP7_75t_L g3122 ( 
.A(n_3011),
.Y(n_3122)
);

BUFx8_ASAP7_75t_L g3123 ( 
.A(n_2720),
.Y(n_3123)
);

INVxp67_ASAP7_75t_L g3124 ( 
.A(n_2741),
.Y(n_3124)
);

BUFx3_ASAP7_75t_L g3125 ( 
.A(n_2701),
.Y(n_3125)
);

INVx2_ASAP7_75t_SL g3126 ( 
.A(n_2745),
.Y(n_3126)
);

NOR2xp33_ASAP7_75t_L g3127 ( 
.A(n_2647),
.B(n_2693),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2841),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2792),
.B(n_2489),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_2841),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2792),
.B(n_2491),
.Y(n_3131)
);

NAND2xp33_ASAP7_75t_L g3132 ( 
.A(n_2766),
.B(n_2043),
.Y(n_3132)
);

HB1xp67_ASAP7_75t_L g3133 ( 
.A(n_2786),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2799),
.B(n_2495),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_SL g3135 ( 
.A(n_2815),
.B(n_2228),
.Y(n_3135)
);

NAND2xp33_ASAP7_75t_L g3136 ( 
.A(n_2766),
.B(n_2043),
.Y(n_3136)
);

INVxp67_ASAP7_75t_L g3137 ( 
.A(n_2799),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2862),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_2737),
.B(n_2239),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2859),
.B(n_2497),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2705),
.B(n_2228),
.Y(n_3141)
);

NAND2xp33_ASAP7_75t_L g3142 ( 
.A(n_2766),
.B(n_2066),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2862),
.Y(n_3143)
);

BUFx6f_ASAP7_75t_L g3144 ( 
.A(n_2654),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_SL g3145 ( 
.A(n_2754),
.B(n_2839),
.Y(n_3145)
);

OR2x6_ASAP7_75t_L g3146 ( 
.A(n_2804),
.B(n_2228),
.Y(n_3146)
);

INVx2_ASAP7_75t_SL g3147 ( 
.A(n_2745),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2897),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2728),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2729),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2859),
.B(n_2498),
.Y(n_3151)
);

BUFx8_ASAP7_75t_L g3152 ( 
.A(n_2836),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2740),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2878),
.B(n_2506),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2756),
.Y(n_3155)
);

BUFx6f_ASAP7_75t_L g3156 ( 
.A(n_2654),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_SL g3157 ( 
.A(n_2821),
.B(n_2231),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_SL g3158 ( 
.A(n_2821),
.B(n_2231),
.Y(n_3158)
);

INVx3_ASAP7_75t_L g3159 ( 
.A(n_2665),
.Y(n_3159)
);

NAND2xp33_ASAP7_75t_L g3160 ( 
.A(n_2766),
.B(n_2066),
.Y(n_3160)
);

OAI221xp5_ASAP7_75t_L g3161 ( 
.A1(n_2785),
.A2(n_2159),
.B1(n_2205),
.B2(n_2251),
.C(n_2246),
.Y(n_3161)
);

INVx2_ASAP7_75t_SL g3162 ( 
.A(n_2736),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2762),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_SL g3164 ( 
.A(n_2873),
.B(n_2241),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2878),
.B(n_2509),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_SL g3166 ( 
.A(n_2873),
.B(n_2241),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2764),
.Y(n_3167)
);

AO22x1_ASAP7_75t_L g3168 ( 
.A1(n_2686),
.A2(n_2075),
.B1(n_2214),
.B2(n_2102),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2892),
.B(n_2725),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_2876),
.B(n_2254),
.Y(n_3170)
);

AOI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_2648),
.A2(n_2513),
.B1(n_2517),
.B2(n_2510),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2772),
.Y(n_3172)
);

AOI221xp5_ASAP7_75t_L g3173 ( 
.A1(n_2986),
.A2(n_2116),
.B1(n_1495),
.B2(n_1496),
.C(n_1493),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2897),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2901),
.Y(n_3175)
);

AOI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_3009),
.A2(n_2093),
.B1(n_2127),
.B2(n_2102),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2774),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2901),
.Y(n_3178)
);

OR2x6_ASAP7_75t_L g3179 ( 
.A(n_2804),
.B(n_2231),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2782),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2892),
.B(n_2518),
.Y(n_3181)
);

AND2x2_ASAP7_75t_L g3182 ( 
.A(n_2812),
.B(n_2244),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2965),
.B(n_2519),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2965),
.B(n_2521),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_SL g3185 ( 
.A(n_2876),
.B(n_2231),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2915),
.B(n_2522),
.Y(n_3186)
);

OAI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_2987),
.A2(n_2370),
.B1(n_2067),
.B2(n_2348),
.Y(n_3187)
);

BUFx3_ASAP7_75t_L g3188 ( 
.A(n_2736),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_3003),
.A2(n_2403),
.B(n_2303),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_2843),
.B(n_2232),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_SL g3191 ( 
.A(n_2810),
.B(n_2235),
.Y(n_3191)
);

AND2x4_ASAP7_75t_L g3192 ( 
.A(n_2747),
.B(n_2771),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2797),
.B(n_2530),
.Y(n_3193)
);

NOR3xp33_ASAP7_75t_L g3194 ( 
.A(n_2806),
.B(n_2483),
.C(n_2461),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2919),
.B(n_2022),
.Y(n_3195)
);

INVxp67_ASAP7_75t_SL g3196 ( 
.A(n_3007),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_2894),
.B(n_2235),
.Y(n_3197)
);

OAI22xp5_ASAP7_75t_L g3198 ( 
.A1(n_3016),
.A2(n_2348),
.B1(n_2358),
.B2(n_2340),
.Y(n_3198)
);

AOI22xp5_ASAP7_75t_L g3199 ( 
.A1(n_2986),
.A2(n_2093),
.B1(n_2136),
.B2(n_2127),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2920),
.Y(n_3200)
);

AND2x4_ASAP7_75t_L g3201 ( 
.A(n_2747),
.B(n_2771),
.Y(n_3201)
);

OAI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_2998),
.A2(n_2514),
.B1(n_2399),
.B2(n_2432),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2790),
.Y(n_3203)
);

NOR2x1_ASAP7_75t_L g3204 ( 
.A(n_2969),
.B(n_2436),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_2698),
.B(n_2022),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2698),
.B(n_2022),
.Y(n_3206)
);

BUFx6f_ASAP7_75t_L g3207 ( 
.A(n_2835),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2920),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2811),
.Y(n_3209)
);

OR2x2_ASAP7_75t_L g3210 ( 
.A(n_2889),
.B(n_2232),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2879),
.B(n_2024),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2880),
.B(n_2024),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2825),
.B(n_2024),
.Y(n_3213)
);

AOI22xp33_ASAP7_75t_L g3214 ( 
.A1(n_2687),
.A2(n_2429),
.B1(n_2430),
.B2(n_2428),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_2825),
.B(n_2398),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2971),
.B(n_2460),
.Y(n_3216)
);

OAI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_2817),
.A2(n_2303),
.B(n_2296),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2932),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_3001),
.B(n_2464),
.Y(n_3219)
);

OAI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_2854),
.A2(n_2358),
.B1(n_2390),
.B2(n_2348),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_3001),
.B(n_2490),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_2655),
.A2(n_2315),
.B(n_2296),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2813),
.Y(n_3223)
);

XOR2xp5_ASAP7_75t_L g3224 ( 
.A(n_2702),
.B(n_2256),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_L g3225 ( 
.A(n_2748),
.B(n_2232),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2816),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2703),
.B(n_2516),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2822),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_SL g3229 ( 
.A(n_2733),
.B(n_2232),
.Y(n_3229)
);

NOR2xp33_ASAP7_75t_L g3230 ( 
.A(n_2750),
.B(n_2235),
.Y(n_3230)
);

NOR2xp33_ASAP7_75t_L g3231 ( 
.A(n_2757),
.B(n_2235),
.Y(n_3231)
);

BUFx2_ASAP7_75t_SL g3232 ( 
.A(n_2969),
.Y(n_3232)
);

INVx4_ASAP7_75t_L g3233 ( 
.A(n_2991),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2844),
.Y(n_3234)
);

INVx2_ASAP7_75t_SL g3235 ( 
.A(n_2755),
.Y(n_3235)
);

INVxp67_ASAP7_75t_L g3236 ( 
.A(n_2703),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2798),
.B(n_2434),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2960),
.B(n_2136),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2960),
.B(n_2058),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2846),
.Y(n_3240)
);

OAI221xp5_ASAP7_75t_L g3241 ( 
.A1(n_3015),
.A2(n_2148),
.B1(n_2115),
.B2(n_2097),
.C(n_2483),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_SL g3242 ( 
.A(n_2733),
.B(n_2864),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2809),
.B(n_2262),
.Y(n_3243)
);

NAND2xp33_ASAP7_75t_L g3244 ( 
.A(n_2766),
.B(n_2492),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_2932),
.Y(n_3245)
);

OR2x2_ASAP7_75t_L g3246 ( 
.A(n_2908),
.B(n_2241),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2645),
.Y(n_3247)
);

OR2x2_ASAP7_75t_L g3248 ( 
.A(n_2958),
.B(n_2241),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2651),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2814),
.B(n_2266),
.Y(n_3250)
);

AOI22xp33_ASAP7_75t_L g3251 ( 
.A1(n_2687),
.A2(n_2270),
.B1(n_2271),
.B2(n_2268),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2746),
.B(n_2899),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_2942),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2900),
.B(n_2272),
.Y(n_3254)
);

AOI22xp5_ASAP7_75t_L g3255 ( 
.A1(n_2974),
.A2(n_2075),
.B1(n_1944),
.B2(n_2000),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_2911),
.B(n_2282),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_2789),
.B(n_2284),
.Y(n_3257)
);

NAND2xp33_ASAP7_75t_L g3258 ( 
.A(n_2665),
.B(n_2493),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_2789),
.B(n_2290),
.Y(n_3259)
);

BUFx2_ASAP7_75t_L g3260 ( 
.A(n_2666),
.Y(n_3260)
);

INVx2_ASAP7_75t_SL g3261 ( 
.A(n_2755),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2805),
.B(n_2831),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_SL g3263 ( 
.A(n_2744),
.B(n_2249),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2805),
.B(n_2291),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2653),
.Y(n_3265)
);

BUFx6f_ASAP7_75t_L g3266 ( 
.A(n_2654),
.Y(n_3266)
);

AOI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_2974),
.A2(n_1944),
.B1(n_2096),
.B2(n_2000),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2662),
.Y(n_3268)
);

OAI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_2927),
.A2(n_2317),
.B(n_2315),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2670),
.Y(n_3270)
);

NOR2xp33_ASAP7_75t_L g3271 ( 
.A(n_2858),
.B(n_2249),
.Y(n_3271)
);

NOR2xp33_ASAP7_75t_L g3272 ( 
.A(n_2866),
.B(n_2249),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2680),
.Y(n_3273)
);

NOR3xp33_ASAP7_75t_L g3274 ( 
.A(n_2926),
.B(n_2500),
.C(n_2195),
.Y(n_3274)
);

AOI22xp5_ASAP7_75t_L g3275 ( 
.A1(n_2726),
.A2(n_2777),
.B1(n_2845),
.B2(n_2893),
.Y(n_3275)
);

AOI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_3010),
.A2(n_2096),
.B1(n_2133),
.B2(n_2110),
.Y(n_3276)
);

NOR2xp33_ASAP7_75t_L g3277 ( 
.A(n_2994),
.B(n_3012),
.Y(n_3277)
);

BUFx6f_ASAP7_75t_L g3278 ( 
.A(n_2713),
.Y(n_3278)
);

NOR2xp33_ASAP7_75t_L g3279 ( 
.A(n_2668),
.B(n_2249),
.Y(n_3279)
);

AND2x4_ASAP7_75t_L g3280 ( 
.A(n_2914),
.B(n_2459),
.Y(n_3280)
);

NOR2xp33_ASAP7_75t_L g3281 ( 
.A(n_2668),
.B(n_2436),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_2831),
.B(n_2294),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_SL g3283 ( 
.A(n_2823),
.B(n_2493),
.Y(n_3283)
);

NOR2xp33_ASAP7_75t_L g3284 ( 
.A(n_2978),
.B(n_2808),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2851),
.Y(n_3285)
);

NOR2xp33_ASAP7_75t_L g3286 ( 
.A(n_2978),
.B(n_2441),
.Y(n_3286)
);

OR2x2_ASAP7_75t_L g3287 ( 
.A(n_2683),
.B(n_2110),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2759),
.B(n_2295),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2942),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_SL g3290 ( 
.A(n_2823),
.B(n_2493),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2852),
.Y(n_3291)
);

INVx3_ASAP7_75t_L g3292 ( 
.A(n_2665),
.Y(n_3292)
);

NOR2xp33_ASAP7_75t_L g3293 ( 
.A(n_2808),
.B(n_2441),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_2954),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2999),
.B(n_2838),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_2954),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2855),
.Y(n_3297)
);

NOR2xp67_ASAP7_75t_L g3298 ( 
.A(n_2739),
.B(n_2486),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3023),
.B(n_2300),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_2914),
.B(n_2301),
.Y(n_3300)
);

BUFx3_ASAP7_75t_L g3301 ( 
.A(n_2941),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_2948),
.B(n_2302),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_2962),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_2940),
.B(n_2493),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_2948),
.B(n_2306),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_2856),
.Y(n_3306)
);

INVxp67_ASAP7_75t_SL g3307 ( 
.A(n_2678),
.Y(n_3307)
);

O2A1O1Ixp33_ASAP7_75t_L g3308 ( 
.A1(n_2655),
.A2(n_2317),
.B(n_2494),
.C(n_2486),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_2666),
.B(n_2133),
.Y(n_3309)
);

OR2x6_ASAP7_75t_L g3310 ( 
.A(n_2804),
.B(n_2580),
.Y(n_3310)
);

NAND2xp33_ASAP7_75t_L g3311 ( 
.A(n_2665),
.B(n_2580),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_2886),
.B(n_2307),
.Y(n_3312)
);

AOI22xp5_ASAP7_75t_L g3313 ( 
.A1(n_2939),
.A2(n_2172),
.B1(n_2500),
.B2(n_2214),
.Y(n_3313)
);

NOR2xp33_ASAP7_75t_L g3314 ( 
.A(n_2910),
.B(n_2494),
.Y(n_3314)
);

BUFx2_ASAP7_75t_L g3315 ( 
.A(n_2666),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_2886),
.B(n_2312),
.Y(n_3316)
);

NOR2xp33_ASAP7_75t_L g3317 ( 
.A(n_2910),
.B(n_2571),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_2886),
.B(n_2314),
.Y(n_3318)
);

BUFx3_ASAP7_75t_L g3319 ( 
.A(n_2849),
.Y(n_3319)
);

INVx2_ASAP7_75t_SL g3320 ( 
.A(n_2780),
.Y(n_3320)
);

OR2x6_ASAP7_75t_L g3321 ( 
.A(n_2776),
.B(n_2580),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2865),
.Y(n_3322)
);

INVxp67_ASAP7_75t_L g3323 ( 
.A(n_2886),
.Y(n_3323)
);

AOI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_2776),
.A2(n_2172),
.B1(n_2214),
.B2(n_2571),
.Y(n_3324)
);

OR2x2_ASAP7_75t_L g3325 ( 
.A(n_2776),
.B(n_2576),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_2886),
.B(n_2325),
.Y(n_3326)
);

AND2x2_ASAP7_75t_L g3327 ( 
.A(n_2788),
.B(n_2195),
.Y(n_3327)
);

BUFx8_ASAP7_75t_L g3328 ( 
.A(n_2778),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_2938),
.B(n_2326),
.Y(n_3329)
);

NAND2xp33_ASAP7_75t_L g3330 ( 
.A(n_2700),
.B(n_2580),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2848),
.B(n_2328),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2848),
.B(n_2329),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_2962),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_2868),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2749),
.B(n_2895),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2869),
.Y(n_3336)
);

INVx1_ASAP7_75t_SL g3337 ( 
.A(n_2803),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_2896),
.B(n_2332),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_2870),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_2988),
.Y(n_3340)
);

BUFx3_ASAP7_75t_L g3341 ( 
.A(n_2956),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3011),
.B(n_2333),
.Y(n_3342)
);

NOR2x1p5_ASAP7_75t_L g3343 ( 
.A(n_2739),
.B(n_1893),
.Y(n_3343)
);

A2O1A1Ixp33_ASAP7_75t_L g3344 ( 
.A1(n_2769),
.A2(n_2584),
.B(n_2588),
.C(n_2576),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2871),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3011),
.B(n_2337),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_SL g3347 ( 
.A(n_3014),
.B(n_2586),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_SL g3348 ( 
.A(n_3019),
.B(n_2586),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_2988),
.Y(n_3349)
);

AOI22xp33_ASAP7_75t_L g3350 ( 
.A1(n_2840),
.A2(n_2341),
.B1(n_2344),
.B2(n_2343),
.Y(n_3350)
);

BUFx6f_ASAP7_75t_L g3351 ( 
.A(n_2713),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_2874),
.Y(n_3352)
);

NOR2xp33_ASAP7_75t_L g3353 ( 
.A(n_2788),
.B(n_2584),
.Y(n_3353)
);

BUFx6f_ASAP7_75t_L g3354 ( 
.A(n_2713),
.Y(n_3354)
);

INVxp67_ASAP7_75t_L g3355 ( 
.A(n_2997),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_SL g3356 ( 
.A(n_2967),
.B(n_2586),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_3011),
.B(n_2347),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_SL g3358 ( 
.A(n_2888),
.B(n_2586),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_L g3359 ( 
.A1(n_2840),
.A2(n_2684),
.B1(n_2807),
.B2(n_2963),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_3017),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2837),
.B(n_2349),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_3017),
.Y(n_3362)
);

CKINVDCx5p33_ASAP7_75t_R g3363 ( 
.A(n_2664),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_2837),
.B(n_2351),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_L g3365 ( 
.A(n_2788),
.B(n_2588),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3025),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_SL g3367 ( 
.A(n_2888),
.B(n_2591),
.Y(n_3367)
);

INVx2_ASAP7_75t_L g3368 ( 
.A(n_3025),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_SL g3369 ( 
.A(n_2956),
.B(n_2591),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_SL g3370 ( 
.A(n_2984),
.B(n_2591),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2652),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_2875),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_SL g3373 ( 
.A(n_2924),
.B(n_2591),
.Y(n_3373)
);

OR2x2_ASAP7_75t_L g3374 ( 
.A(n_2972),
.B(n_2598),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_2657),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_2661),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_2882),
.Y(n_3377)
);

NAND2xp33_ASAP7_75t_L g3378 ( 
.A(n_2700),
.B(n_2600),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_2663),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3371),
.Y(n_3380)
);

INVx2_ASAP7_75t_L g3381 ( 
.A(n_3375),
.Y(n_3381)
);

HB1xp67_ASAP7_75t_L g3382 ( 
.A(n_3056),
.Y(n_3382)
);

OAI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_3103),
.A2(n_2872),
.B(n_2927),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3058),
.B(n_2997),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3033),
.Y(n_3385)
);

INVx4_ASAP7_75t_L g3386 ( 
.A(n_3094),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3376),
.Y(n_3387)
);

INVx3_ASAP7_75t_L g3388 ( 
.A(n_3094),
.Y(n_3388)
);

AND2x2_ASAP7_75t_L g3389 ( 
.A(n_3100),
.B(n_3098),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3219),
.B(n_3221),
.Y(n_3390)
);

AOI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3199),
.A2(n_2664),
.B1(n_2917),
.B2(n_2819),
.Y(n_3391)
);

OAI22xp5_ASAP7_75t_SL g3392 ( 
.A1(n_3176),
.A2(n_2840),
.B1(n_2963),
.B2(n_2724),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3379),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3042),
.Y(n_3394)
);

AND2x4_ASAP7_75t_L g3395 ( 
.A(n_3192),
.B(n_2742),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_3236),
.B(n_2803),
.Y(n_3396)
);

BUFx3_ASAP7_75t_L g3397 ( 
.A(n_3152),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_SL g3398 ( 
.A(n_3097),
.B(n_2924),
.Y(n_3398)
);

AND2x4_ASAP7_75t_L g3399 ( 
.A(n_3192),
.B(n_2742),
.Y(n_3399)
);

INVx3_ASAP7_75t_L g3400 ( 
.A(n_3094),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3051),
.Y(n_3401)
);

CKINVDCx5p33_ASAP7_75t_R g3402 ( 
.A(n_3114),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3029),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3054),
.Y(n_3404)
);

INVx3_ASAP7_75t_L g3405 ( 
.A(n_3122),
.Y(n_3405)
);

NOR2x1p5_ASAP7_75t_L g3406 ( 
.A(n_3238),
.B(n_2768),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3055),
.Y(n_3407)
);

INVx4_ASAP7_75t_L g3408 ( 
.A(n_3122),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_3035),
.Y(n_3409)
);

A2O1A1Ixp33_ASAP7_75t_L g3410 ( 
.A1(n_3031),
.A2(n_2917),
.B(n_2973),
.C(n_2684),
.Y(n_3410)
);

AND2x2_ASAP7_75t_SL g3411 ( 
.A(n_3359),
.B(n_3214),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_SL g3412 ( 
.A(n_3097),
.B(n_2924),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3056),
.B(n_2972),
.Y(n_3413)
);

AOI22xp33_ASAP7_75t_L g3414 ( 
.A1(n_3359),
.A2(n_2997),
.B1(n_2898),
.B2(n_2906),
.Y(n_3414)
);

BUFx6f_ASAP7_75t_L g3415 ( 
.A(n_3122),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3065),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_3041),
.Y(n_3417)
);

AO22x1_ASAP7_75t_L g3418 ( 
.A1(n_3034),
.A2(n_2834),
.B1(n_2768),
.B2(n_2711),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_3045),
.Y(n_3419)
);

AOI22xp5_ASAP7_75t_L g3420 ( 
.A1(n_3139),
.A2(n_2867),
.B1(n_2972),
.B2(n_2763),
.Y(n_3420)
);

OAI22xp5_ASAP7_75t_SL g3421 ( 
.A1(n_3161),
.A2(n_2906),
.B1(n_2898),
.B2(n_3006),
.Y(n_3421)
);

INVx2_ASAP7_75t_SL g3422 ( 
.A(n_3152),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_SL g3423 ( 
.A(n_3236),
.B(n_2924),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_3073),
.B(n_2977),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3048),
.Y(n_3425)
);

AOI22xp5_ASAP7_75t_L g3426 ( 
.A1(n_3139),
.A2(n_2867),
.B1(n_2763),
.B2(n_2973),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_3276),
.B(n_3071),
.Y(n_3427)
);

AND2x2_ASAP7_75t_SL g3428 ( 
.A(n_3214),
.B(n_2853),
.Y(n_3428)
);

INVx2_ASAP7_75t_SL g3429 ( 
.A(n_3123),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3064),
.B(n_2997),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3057),
.Y(n_3431)
);

AOI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_3064),
.A2(n_2872),
.B(n_2933),
.Y(n_3432)
);

BUFx3_ASAP7_75t_L g3433 ( 
.A(n_3319),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3070),
.Y(n_3434)
);

NAND2x1p5_ASAP7_75t_L g3435 ( 
.A(n_3107),
.B(n_2977),
.Y(n_3435)
);

BUFx3_ASAP7_75t_L g3436 ( 
.A(n_3123),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_3075),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3196),
.B(n_2997),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3196),
.B(n_2887),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_SL g3440 ( 
.A(n_3137),
.B(n_2977),
.Y(n_3440)
);

AOI22xp33_ASAP7_75t_L g3441 ( 
.A1(n_3081),
.A2(n_2898),
.B1(n_2906),
.B2(n_2689),
.Y(n_3441)
);

INVx6_ASAP7_75t_L g3442 ( 
.A(n_3328),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3295),
.B(n_2903),
.Y(n_3443)
);

NOR2xp33_ASAP7_75t_L g3444 ( 
.A(n_3066),
.B(n_3006),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3072),
.Y(n_3445)
);

AND2x4_ASAP7_75t_L g3446 ( 
.A(n_3201),
.B(n_3004),
.Y(n_3446)
);

AOI22xp5_ASAP7_75t_L g3447 ( 
.A1(n_3111),
.A2(n_2867),
.B1(n_2975),
.B2(n_2711),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3078),
.Y(n_3448)
);

INVx2_ASAP7_75t_SL g3449 ( 
.A(n_3096),
.Y(n_3449)
);

INVx2_ASAP7_75t_SL g3450 ( 
.A(n_3096),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_SL g3451 ( 
.A(n_3137),
.B(n_2977),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3088),
.B(n_2883),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3086),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3081),
.A2(n_2689),
.B1(n_2779),
.B2(n_2695),
.Y(n_3454)
);

AND2x4_ASAP7_75t_L g3455 ( 
.A(n_3201),
.B(n_3004),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3101),
.Y(n_3456)
);

NOR2xp33_ASAP7_75t_L g3457 ( 
.A(n_3049),
.B(n_2105),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3102),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3090),
.B(n_2907),
.Y(n_3459)
);

NOR2x1p5_ASAP7_75t_L g3460 ( 
.A(n_3083),
.B(n_2738),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_SL g3461 ( 
.A(n_3213),
.B(n_2704),
.Y(n_3461)
);

INVx5_ASAP7_75t_L g3462 ( 
.A(n_3321),
.Y(n_3462)
);

INVx4_ASAP7_75t_L g3463 ( 
.A(n_3110),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3140),
.B(n_2909),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3151),
.B(n_2913),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3154),
.B(n_2916),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3109),
.Y(n_3467)
);

NAND3xp33_ASAP7_75t_L g3468 ( 
.A(n_3034),
.B(n_2431),
.C(n_2639),
.Y(n_3468)
);

AND2x4_ASAP7_75t_L g3469 ( 
.A(n_3105),
.B(n_3004),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3165),
.B(n_2918),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3117),
.Y(n_3471)
);

AOI22xp5_ASAP7_75t_L g3472 ( 
.A1(n_3111),
.A2(n_2975),
.B1(n_2700),
.B2(n_2711),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_R g3473 ( 
.A(n_3363),
.B(n_2700),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3121),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_3031),
.B(n_2704),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3149),
.Y(n_3476)
);

OAI22xp5_ASAP7_75t_L g3477 ( 
.A1(n_3044),
.A2(n_2779),
.B1(n_2695),
.B2(n_2863),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_SL g3478 ( 
.A(n_3032),
.B(n_2704),
.Y(n_3478)
);

NOR3xp33_ASAP7_75t_L g3479 ( 
.A(n_3241),
.B(n_2715),
.C(n_2690),
.Y(n_3479)
);

NOR2xp33_ASAP7_75t_L g3480 ( 
.A(n_3267),
.B(n_1960),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3091),
.B(n_3099),
.Y(n_3481)
);

AOI22xp5_ASAP7_75t_L g3482 ( 
.A1(n_3170),
.A2(n_2975),
.B1(n_2711),
.B2(n_2598),
.Y(n_3482)
);

INVx3_ASAP7_75t_L g3483 ( 
.A(n_3310),
.Y(n_3483)
);

OR2x2_ASAP7_75t_L g3484 ( 
.A(n_3287),
.B(n_2658),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3182),
.B(n_779),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3150),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3084),
.Y(n_3487)
);

INVx5_ASAP7_75t_L g3488 ( 
.A(n_3321),
.Y(n_3488)
);

A2O1A1Ixp33_ASAP7_75t_L g3489 ( 
.A1(n_3032),
.A2(n_2877),
.B(n_2850),
.C(n_2715),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3153),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3087),
.Y(n_3491)
);

AOI22xp33_ASAP7_75t_L g3492 ( 
.A1(n_3089),
.A2(n_2904),
.B1(n_2975),
.B2(n_2928),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_SL g3493 ( 
.A(n_3104),
.B(n_2704),
.Y(n_3493)
);

BUFx6f_ASAP7_75t_L g3494 ( 
.A(n_3096),
.Y(n_3494)
);

BUFx3_ASAP7_75t_L g3495 ( 
.A(n_3125),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_R g3496 ( 
.A(n_3040),
.B(n_2711),
.Y(n_3496)
);

INVx1_ASAP7_75t_SL g3497 ( 
.A(n_3085),
.Y(n_3497)
);

HB1xp67_ASAP7_75t_L g3498 ( 
.A(n_3124),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3183),
.B(n_3184),
.Y(n_3499)
);

INVxp67_ASAP7_75t_SL g3500 ( 
.A(n_3307),
.Y(n_3500)
);

BUFx6f_ASAP7_75t_L g3501 ( 
.A(n_3207),
.Y(n_3501)
);

AND2x4_ASAP7_75t_SL g3502 ( 
.A(n_3110),
.B(n_2738),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_3108),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3128),
.Y(n_3504)
);

INVx4_ASAP7_75t_L g3505 ( 
.A(n_3233),
.Y(n_3505)
);

AND2x2_ASAP7_75t_L g3506 ( 
.A(n_3080),
.B(n_934),
.Y(n_3506)
);

INVx3_ASAP7_75t_L g3507 ( 
.A(n_3310),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3215),
.B(n_2921),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_SL g3509 ( 
.A(n_3205),
.B(n_2708),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_3130),
.Y(n_3510)
);

INVx3_ASAP7_75t_L g3511 ( 
.A(n_3310),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_3138),
.Y(n_3512)
);

INVx3_ASAP7_75t_L g3513 ( 
.A(n_3159),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3186),
.B(n_2931),
.Y(n_3514)
);

INVx3_ASAP7_75t_L g3515 ( 
.A(n_3159),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3155),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3163),
.Y(n_3517)
);

INVx2_ASAP7_75t_SL g3518 ( 
.A(n_3207),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3193),
.B(n_2936),
.Y(n_3519)
);

INVx5_ASAP7_75t_L g3520 ( 
.A(n_3321),
.Y(n_3520)
);

A2O1A1Ixp33_ASAP7_75t_L g3521 ( 
.A1(n_3082),
.A2(n_2877),
.B(n_2850),
.C(n_2719),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3335),
.B(n_2937),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3167),
.Y(n_3523)
);

OAI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3068),
.A2(n_2863),
.B1(n_2673),
.B2(n_2658),
.Y(n_3524)
);

INVx4_ASAP7_75t_L g3525 ( 
.A(n_3233),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3143),
.Y(n_3526)
);

A2O1A1Ixp33_ASAP7_75t_L g3527 ( 
.A1(n_3082),
.A2(n_2719),
.B(n_2743),
.C(n_2690),
.Y(n_3527)
);

CKINVDCx5p33_ASAP7_75t_R g3528 ( 
.A(n_3301),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3172),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3148),
.Y(n_3530)
);

AND2x2_ASAP7_75t_L g3531 ( 
.A(n_3080),
.B(n_934),
.Y(n_3531)
);

AND2x4_ASAP7_75t_L g3532 ( 
.A(n_3105),
.B(n_2794),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3174),
.Y(n_3533)
);

BUFx3_ASAP7_75t_L g3534 ( 
.A(n_3188),
.Y(n_3534)
);

BUFx8_ASAP7_75t_L g3535 ( 
.A(n_3037),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3175),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3177),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_SL g3538 ( 
.A(n_3206),
.B(n_2708),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3119),
.B(n_2943),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3178),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3180),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3200),
.Y(n_3542)
);

OR2x2_ASAP7_75t_L g3543 ( 
.A(n_3043),
.B(n_2673),
.Y(n_3543)
);

INVx2_ASAP7_75t_SL g3544 ( 
.A(n_3207),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3120),
.B(n_3129),
.Y(n_3545)
);

AND2x4_ASAP7_75t_L g3546 ( 
.A(n_3280),
.B(n_2794),
.Y(n_3546)
);

BUFx6f_ASAP7_75t_L g3547 ( 
.A(n_3052),
.Y(n_3547)
);

OAI221xp5_ASAP7_75t_L g3548 ( 
.A1(n_3173),
.A2(n_1500),
.B1(n_1504),
.B2(n_1497),
.C(n_1492),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3203),
.Y(n_3549)
);

AND2x2_ASAP7_75t_L g3550 ( 
.A(n_3133),
.B(n_934),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3131),
.B(n_2946),
.Y(n_3551)
);

A2O1A1Ixp33_ASAP7_75t_L g3552 ( 
.A1(n_3077),
.A2(n_2753),
.B(n_2743),
.C(n_2818),
.Y(n_3552)
);

INVx3_ASAP7_75t_L g3553 ( 
.A(n_3292),
.Y(n_3553)
);

OR2x2_ASAP7_75t_L g3554 ( 
.A(n_3133),
.B(n_2950),
.Y(n_3554)
);

OAI22xp5_ASAP7_75t_L g3555 ( 
.A1(n_3069),
.A2(n_2847),
.B1(n_2891),
.B2(n_2842),
.Y(n_3555)
);

BUFx2_ASAP7_75t_L g3556 ( 
.A(n_3124),
.Y(n_3556)
);

INVx1_ASAP7_75t_SL g3557 ( 
.A(n_3248),
.Y(n_3557)
);

INVx3_ASAP7_75t_L g3558 ( 
.A(n_3292),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3134),
.B(n_2951),
.Y(n_3559)
);

AOI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_3258),
.A2(n_2970),
.B(n_2933),
.Y(n_3560)
);

BUFx6f_ASAP7_75t_L g3561 ( 
.A(n_3052),
.Y(n_3561)
);

AOI22xp33_ASAP7_75t_L g3562 ( 
.A1(n_3089),
.A2(n_2904),
.B1(n_2975),
.B2(n_2957),
.Y(n_3562)
);

INVx5_ASAP7_75t_L g3563 ( 
.A(n_3146),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3209),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3223),
.Y(n_3565)
);

OAI22xp5_ASAP7_75t_L g3566 ( 
.A1(n_3169),
.A2(n_2847),
.B1(n_2891),
.B2(n_2842),
.Y(n_3566)
);

NOR2x1p5_ASAP7_75t_L g3567 ( 
.A(n_3341),
.B(n_2833),
.Y(n_3567)
);

BUFx6f_ASAP7_75t_L g3568 ( 
.A(n_3052),
.Y(n_3568)
);

NOR2xp33_ASAP7_75t_L g3569 ( 
.A(n_3118),
.B(n_3021),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_SL g3570 ( 
.A(n_3277),
.B(n_2708),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3277),
.B(n_2952),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3226),
.Y(n_3572)
);

INVx5_ASAP7_75t_L g3573 ( 
.A(n_3146),
.Y(n_3573)
);

AOI22xp33_ASAP7_75t_L g3574 ( 
.A1(n_3092),
.A2(n_2961),
.B1(n_2964),
.B2(n_2959),
.Y(n_3574)
);

AND3x2_ASAP7_75t_SL g3575 ( 
.A(n_3168),
.B(n_1340),
.C(n_2537),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3228),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_3208),
.Y(n_3577)
);

AOI22xp33_ASAP7_75t_L g3578 ( 
.A1(n_3092),
.A2(n_2990),
.B1(n_3005),
.B2(n_2968),
.Y(n_3578)
);

AND2x2_ASAP7_75t_SL g3579 ( 
.A(n_3251),
.B(n_2833),
.Y(n_3579)
);

AND2x2_ASAP7_75t_SL g3580 ( 
.A(n_3251),
.B(n_3000),
.Y(n_3580)
);

NAND3xp33_ASAP7_75t_L g3581 ( 
.A(n_3047),
.B(n_2753),
.C(n_2773),
.Y(n_3581)
);

INVx2_ASAP7_75t_L g3582 ( 
.A(n_3218),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3299),
.B(n_3008),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_SL g3584 ( 
.A(n_3077),
.B(n_2708),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_SL g3585 ( 
.A(n_3252),
.B(n_2713),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3338),
.B(n_3020),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3227),
.B(n_3039),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3234),
.Y(n_3588)
);

HB1xp67_ASAP7_75t_L g3589 ( 
.A(n_3118),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3245),
.Y(n_3590)
);

HB1xp67_ASAP7_75t_L g3591 ( 
.A(n_3060),
.Y(n_3591)
);

AND2x4_ASAP7_75t_L g3592 ( 
.A(n_3280),
.B(n_2794),
.Y(n_3592)
);

INVxp67_ASAP7_75t_SL g3593 ( 
.A(n_3307),
.Y(n_3593)
);

OAI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_3039),
.A2(n_2818),
.B1(n_2773),
.B2(n_911),
.Y(n_3594)
);

NAND2x1_ASAP7_75t_L g3595 ( 
.A(n_3052),
.B(n_2761),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3253),
.Y(n_3596)
);

CKINVDCx5p33_ASAP7_75t_R g3597 ( 
.A(n_3037),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3189),
.B(n_3024),
.Y(n_3598)
);

BUFx2_ASAP7_75t_L g3599 ( 
.A(n_3309),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3189),
.B(n_3329),
.Y(n_3600)
);

INVx4_ASAP7_75t_L g3601 ( 
.A(n_3144),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3289),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3047),
.B(n_3026),
.Y(n_3603)
);

INVx2_ASAP7_75t_SL g3604 ( 
.A(n_3328),
.Y(n_3604)
);

AOI22xp33_ASAP7_75t_L g3605 ( 
.A1(n_3171),
.A2(n_3027),
.B1(n_2359),
.B2(n_2361),
.Y(n_3605)
);

AOI22xp33_ASAP7_75t_L g3606 ( 
.A1(n_3171),
.A2(n_2366),
.B1(n_2371),
.B2(n_2356),
.Y(n_3606)
);

INVx2_ASAP7_75t_L g3607 ( 
.A(n_3294),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3059),
.B(n_2678),
.Y(n_3608)
);

AOI22xp33_ASAP7_75t_L g3609 ( 
.A1(n_3170),
.A2(n_2376),
.B1(n_2388),
.B2(n_2372),
.Y(n_3609)
);

AOI22xp5_ASAP7_75t_L g3610 ( 
.A1(n_3127),
.A2(n_2732),
.B1(n_2358),
.B2(n_2391),
.Y(n_3610)
);

AOI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3127),
.A2(n_2732),
.B1(n_2390),
.B2(n_2414),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3240),
.Y(n_3612)
);

BUFx8_ASAP7_75t_L g3613 ( 
.A(n_3320),
.Y(n_3613)
);

INVxp33_ASAP7_75t_L g3614 ( 
.A(n_3224),
.Y(n_3614)
);

AOI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_3311),
.A2(n_3378),
.B(n_3330),
.Y(n_3615)
);

AND2x4_ASAP7_75t_L g3616 ( 
.A(n_3146),
.B(n_2995),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3247),
.Y(n_3617)
);

INVx1_ASAP7_75t_SL g3618 ( 
.A(n_3246),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3249),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_SL g3620 ( 
.A(n_3060),
.B(n_2751),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_3244),
.A2(n_2970),
.B(n_2829),
.Y(n_3621)
);

AND2x4_ASAP7_75t_L g3622 ( 
.A(n_3179),
.B(n_2995),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3265),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3268),
.Y(n_3624)
);

BUFx10_ASAP7_75t_L g3625 ( 
.A(n_3063),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_3132),
.A2(n_2829),
.B(n_2709),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3059),
.B(n_3000),
.Y(n_3627)
);

NOR2xp33_ASAP7_75t_L g3628 ( 
.A(n_3284),
.B(n_2857),
.Y(n_3628)
);

INVx3_ASAP7_75t_L g3629 ( 
.A(n_3144),
.Y(n_3629)
);

INVx3_ASAP7_75t_L g3630 ( 
.A(n_3144),
.Y(n_3630)
);

HB1xp67_ASAP7_75t_L g3631 ( 
.A(n_3284),
.Y(n_3631)
);

OR2x6_ASAP7_75t_L g3632 ( 
.A(n_3179),
.B(n_3232),
.Y(n_3632)
);

AND2x2_ASAP7_75t_L g3633 ( 
.A(n_3190),
.B(n_934),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3270),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3296),
.Y(n_3635)
);

BUFx3_ASAP7_75t_L g3636 ( 
.A(n_3162),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3243),
.B(n_2761),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3273),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3285),
.Y(n_3639)
);

AND2x2_ASAP7_75t_SL g3640 ( 
.A(n_3136),
.B(n_2983),
.Y(n_3640)
);

CKINVDCx5p33_ASAP7_75t_R g3641 ( 
.A(n_3337),
.Y(n_3641)
);

AOI22xp33_ASAP7_75t_L g3642 ( 
.A1(n_3195),
.A2(n_2674),
.B1(n_2691),
.B2(n_2671),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3250),
.B(n_2801),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3291),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3254),
.B(n_2801),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3303),
.Y(n_3646)
);

AND2x6_ASAP7_75t_SL g3647 ( 
.A(n_3327),
.B(n_912),
.Y(n_3647)
);

AOI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3211),
.A2(n_2770),
.B1(n_2787),
.B2(n_2752),
.Y(n_3648)
);

NOR2xp33_ASAP7_75t_R g3649 ( 
.A(n_3030),
.B(n_2925),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3297),
.Y(n_3650)
);

NAND2xp33_ASAP7_75t_L g3651 ( 
.A(n_3262),
.B(n_2751),
.Y(n_3651)
);

AOI21xp5_ASAP7_75t_L g3652 ( 
.A1(n_3142),
.A2(n_2709),
.B(n_2860),
.Y(n_3652)
);

AOI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3225),
.A2(n_2390),
.B1(n_2414),
.B2(n_2391),
.Y(n_3653)
);

CKINVDCx5p33_ASAP7_75t_R g3654 ( 
.A(n_3235),
.Y(n_3654)
);

BUFx6f_ASAP7_75t_L g3655 ( 
.A(n_3144),
.Y(n_3655)
);

BUFx3_ASAP7_75t_L g3656 ( 
.A(n_3261),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3225),
.B(n_1030),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_SL g3658 ( 
.A(n_3324),
.B(n_2751),
.Y(n_3658)
);

AOI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3230),
.A2(n_3231),
.B1(n_3365),
.B2(n_3353),
.Y(n_3659)
);

NOR2xp33_ASAP7_75t_L g3660 ( 
.A(n_3242),
.B(n_2857),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3306),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_SL g3662 ( 
.A(n_3587),
.B(n_3198),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3390),
.B(n_3230),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_SL g3664 ( 
.A(n_3587),
.B(n_3194),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3390),
.B(n_3231),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3410),
.B(n_3194),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_SL g3667 ( 
.A(n_3428),
.B(n_3202),
.Y(n_3667)
);

NAND2xp33_ASAP7_75t_SL g3668 ( 
.A(n_3473),
.B(n_3343),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3499),
.B(n_3481),
.Y(n_3669)
);

NAND2xp33_ASAP7_75t_SL g3670 ( 
.A(n_3496),
.B(n_3095),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_SL g3671 ( 
.A(n_3608),
.B(n_3202),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_SL g3672 ( 
.A(n_3608),
.B(n_3271),
.Y(n_3672)
);

AND2x2_ASAP7_75t_L g3673 ( 
.A(n_3389),
.B(n_3067),
.Y(n_3673)
);

AND2x4_ASAP7_75t_L g3674 ( 
.A(n_3462),
.B(n_3355),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_SL g3675 ( 
.A(n_3499),
.B(n_3271),
.Y(n_3675)
);

NAND2xp33_ASAP7_75t_SL g3676 ( 
.A(n_3528),
.B(n_3604),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_SL g3677 ( 
.A(n_3579),
.B(n_3274),
.Y(n_3677)
);

NAND2xp33_ASAP7_75t_SL g3678 ( 
.A(n_3567),
.B(n_3076),
.Y(n_3678)
);

NAND2xp33_ASAP7_75t_SL g3679 ( 
.A(n_3649),
.B(n_3406),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_3631),
.B(n_3210),
.Y(n_3680)
);

NAND2xp33_ASAP7_75t_SL g3681 ( 
.A(n_3591),
.B(n_3050),
.Y(n_3681)
);

NAND2xp33_ASAP7_75t_SL g3682 ( 
.A(n_3460),
.B(n_3106),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_SL g3683 ( 
.A(n_3391),
.B(n_3274),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_SL g3684 ( 
.A(n_3472),
.B(n_3272),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_SL g3685 ( 
.A(n_3426),
.B(n_3272),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_SL g3686 ( 
.A(n_3481),
.B(n_3313),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_SL g3687 ( 
.A(n_3447),
.B(n_3571),
.Y(n_3687)
);

AND2x4_ASAP7_75t_L g3688 ( 
.A(n_3462),
.B(n_3355),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_SL g3689 ( 
.A(n_3571),
.B(n_3350),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_SL g3690 ( 
.A(n_3392),
.B(n_3350),
.Y(n_3690)
);

NAND2xp33_ASAP7_75t_SL g3691 ( 
.A(n_3382),
.B(n_3421),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3485),
.B(n_3275),
.Y(n_3692)
);

NAND2xp33_ASAP7_75t_SL g3693 ( 
.A(n_3386),
.B(n_3181),
.Y(n_3693)
);

AND2x4_ASAP7_75t_L g3694 ( 
.A(n_3462),
.B(n_3156),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_SL g3695 ( 
.A(n_3545),
.B(n_3353),
.Y(n_3695)
);

NAND2xp33_ASAP7_75t_SL g3696 ( 
.A(n_3386),
.B(n_3263),
.Y(n_3696)
);

AND2x2_ASAP7_75t_L g3697 ( 
.A(n_3633),
.B(n_3279),
.Y(n_3697)
);

NAND2xp33_ASAP7_75t_SL g3698 ( 
.A(n_3408),
.B(n_3116),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_SL g3699 ( 
.A(n_3545),
.B(n_3365),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_SL g3700 ( 
.A(n_3659),
.B(n_3156),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3427),
.B(n_3237),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_SL g3702 ( 
.A(n_3640),
.B(n_3156),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_SL g3703 ( 
.A(n_3627),
.B(n_3156),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_SL g3704 ( 
.A(n_3627),
.B(n_3266),
.Y(n_3704)
);

AND2x4_ASAP7_75t_L g3705 ( 
.A(n_3462),
.B(n_3266),
.Y(n_3705)
);

AND2x4_ASAP7_75t_L g3706 ( 
.A(n_3488),
.B(n_3266),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_SL g3707 ( 
.A(n_3482),
.B(n_3266),
.Y(n_3707)
);

AND2x2_ASAP7_75t_L g3708 ( 
.A(n_3506),
.B(n_3279),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_SL g3709 ( 
.A(n_3603),
.B(n_3278),
.Y(n_3709)
);

NAND2xp33_ASAP7_75t_SL g3710 ( 
.A(n_3408),
.B(n_3126),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_SL g3711 ( 
.A(n_3603),
.B(n_3278),
.Y(n_3711)
);

NAND2xp33_ASAP7_75t_SL g3712 ( 
.A(n_3498),
.B(n_3589),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_SL g3713 ( 
.A(n_3444),
.B(n_3278),
.Y(n_3713)
);

AND2x4_ASAP7_75t_L g3714 ( 
.A(n_3488),
.B(n_3278),
.Y(n_3714)
);

NAND2xp33_ASAP7_75t_SL g3715 ( 
.A(n_3556),
.B(n_3147),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3531),
.B(n_3260),
.Y(n_3716)
);

NAND2xp33_ASAP7_75t_SL g3717 ( 
.A(n_3415),
.B(n_3079),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3497),
.B(n_3557),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_SL g3719 ( 
.A(n_3524),
.B(n_3351),
.Y(n_3719)
);

AND2x4_ASAP7_75t_L g3720 ( 
.A(n_3488),
.B(n_3351),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3550),
.B(n_3315),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_SL g3722 ( 
.A(n_3524),
.B(n_3351),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_SL g3723 ( 
.A(n_3384),
.B(n_3351),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3599),
.B(n_3255),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3497),
.B(n_3293),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_SL g3726 ( 
.A(n_3384),
.B(n_3354),
.Y(n_3726)
);

NAND2xp33_ASAP7_75t_SL g3727 ( 
.A(n_3415),
.B(n_3429),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_3657),
.B(n_3293),
.Y(n_3728)
);

NAND2xp33_ASAP7_75t_SL g3729 ( 
.A(n_3415),
.B(n_3112),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3557),
.B(n_3314),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_3615),
.B(n_3354),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3618),
.B(n_3314),
.Y(n_3732)
);

NAND2xp33_ASAP7_75t_SL g3733 ( 
.A(n_3463),
.B(n_3061),
.Y(n_3733)
);

NAND2xp33_ASAP7_75t_SL g3734 ( 
.A(n_3463),
.B(n_3239),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_SL g3735 ( 
.A(n_3411),
.B(n_3354),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3618),
.B(n_3317),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_SL g3737 ( 
.A(n_3420),
.B(n_3354),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_SL g3738 ( 
.A(n_3580),
.B(n_3038),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3413),
.B(n_3317),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_SL g3740 ( 
.A(n_3494),
.B(n_3281),
.Y(n_3740)
);

NAND2xp33_ASAP7_75t_SL g3741 ( 
.A(n_3505),
.B(n_3062),
.Y(n_3741)
);

NAND2xp33_ASAP7_75t_SL g3742 ( 
.A(n_3505),
.B(n_3074),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_SL g3743 ( 
.A(n_3494),
.B(n_3501),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3628),
.B(n_3113),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_SL g3745 ( 
.A(n_3494),
.B(n_3281),
.Y(n_3745)
);

AND2x4_ASAP7_75t_L g3746 ( 
.A(n_3488),
.B(n_3323),
.Y(n_3746)
);

NAND2xp33_ASAP7_75t_SL g3747 ( 
.A(n_3525),
.B(n_3135),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_SL g3748 ( 
.A(n_3501),
.B(n_3298),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3554),
.B(n_3286),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_SL g3750 ( 
.A(n_3501),
.B(n_3145),
.Y(n_3750)
);

NAND2xp33_ASAP7_75t_SL g3751 ( 
.A(n_3525),
.B(n_3093),
.Y(n_3751)
);

NOR2xp33_ASAP7_75t_L g3752 ( 
.A(n_3614),
.B(n_3053),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_SL g3753 ( 
.A(n_3570),
.B(n_3361),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_SL g3754 ( 
.A(n_3555),
.B(n_3364),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_SL g3755 ( 
.A(n_3555),
.B(n_3304),
.Y(n_3755)
);

NAND2xp33_ASAP7_75t_SL g3756 ( 
.A(n_3641),
.B(n_3212),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_SL g3757 ( 
.A(n_3493),
.B(n_3323),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3443),
.B(n_3286),
.Y(n_3758)
);

AND2x2_ASAP7_75t_SL g3759 ( 
.A(n_3441),
.B(n_3160),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_SL g3760 ( 
.A(n_3464),
.B(n_3325),
.Y(n_3760)
);

NAND2xp33_ASAP7_75t_SL g3761 ( 
.A(n_3402),
.B(n_2751),
.Y(n_3761)
);

NAND2xp33_ASAP7_75t_SL g3762 ( 
.A(n_3654),
.B(n_2781),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_3396),
.B(n_3204),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_SL g3764 ( 
.A(n_3464),
.B(n_3187),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3543),
.B(n_3173),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_SL g3766 ( 
.A(n_3465),
.B(n_3466),
.Y(n_3766)
);

NAND2xp33_ASAP7_75t_SL g3767 ( 
.A(n_3388),
.B(n_3400),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3443),
.B(n_3141),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3508),
.B(n_3334),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3508),
.B(n_3336),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_SL g3771 ( 
.A(n_3465),
.B(n_3348),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_3385),
.B(n_3339),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_SL g3773 ( 
.A(n_3466),
.B(n_3300),
.Y(n_3773)
);

NAND2x1_ASAP7_75t_L g3774 ( 
.A(n_3601),
.B(n_2983),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_SL g3775 ( 
.A(n_3470),
.B(n_3302),
.Y(n_3775)
);

NAND2xp33_ASAP7_75t_SL g3776 ( 
.A(n_3388),
.B(n_2781),
.Y(n_3776)
);

AND2x4_ASAP7_75t_L g3777 ( 
.A(n_3520),
.B(n_3322),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_SL g3778 ( 
.A(n_3470),
.B(n_3305),
.Y(n_3778)
);

NAND2xp33_ASAP7_75t_SL g3779 ( 
.A(n_3400),
.B(n_2781),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_SL g3780 ( 
.A(n_3479),
.B(n_3374),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3394),
.B(n_3345),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_SL g3782 ( 
.A(n_3522),
.B(n_3331),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3401),
.B(n_3352),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_SL g3784 ( 
.A(n_3522),
.B(n_3332),
.Y(n_3784)
);

NAND2xp33_ASAP7_75t_SL g3785 ( 
.A(n_3405),
.B(n_2781),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_SL g3786 ( 
.A(n_3452),
.B(n_3459),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_SL g3787 ( 
.A(n_3452),
.B(n_3342),
.Y(n_3787)
);

NAND2xp33_ASAP7_75t_SL g3788 ( 
.A(n_3405),
.B(n_2828),
.Y(n_3788)
);

AND2x2_ASAP7_75t_L g3789 ( 
.A(n_3457),
.B(n_1030),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_SL g3790 ( 
.A(n_3459),
.B(n_3346),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_SL g3791 ( 
.A(n_3475),
.B(n_3357),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_SL g3792 ( 
.A(n_3478),
.B(n_3521),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_SL g3793 ( 
.A(n_3581),
.B(n_3018),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_SL g3794 ( 
.A(n_3581),
.B(n_3018),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_SL g3795 ( 
.A(n_3584),
.B(n_3018),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_SL g3796 ( 
.A(n_3610),
.B(n_3018),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_SL g3797 ( 
.A(n_3611),
.B(n_3028),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3433),
.B(n_3569),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_SL g3799 ( 
.A(n_3527),
.B(n_3028),
.Y(n_3799)
);

NAND2xp33_ASAP7_75t_SL g3800 ( 
.A(n_3422),
.B(n_3597),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_SL g3801 ( 
.A(n_3616),
.B(n_3028),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_SL g3802 ( 
.A(n_3616),
.B(n_3028),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_SL g3803 ( 
.A(n_3622),
.B(n_2828),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3404),
.B(n_3372),
.Y(n_3804)
);

NAND2xp33_ASAP7_75t_SL g3805 ( 
.A(n_3423),
.B(n_2828),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3407),
.B(n_3377),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_SL g3807 ( 
.A(n_3622),
.B(n_2828),
.Y(n_3807)
);

NAND2xp33_ASAP7_75t_SL g3808 ( 
.A(n_3547),
.B(n_2830),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_SL g3809 ( 
.A(n_3566),
.B(n_2830),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_SL g3810 ( 
.A(n_3566),
.B(n_2830),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3416),
.B(n_3164),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_SL g3812 ( 
.A(n_3653),
.B(n_2830),
.Y(n_3812)
);

NAND2xp33_ASAP7_75t_SL g3813 ( 
.A(n_3547),
.B(n_3257),
.Y(n_3813)
);

AND2x2_ASAP7_75t_L g3814 ( 
.A(n_3484),
.B(n_1030),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_3445),
.B(n_3166),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_SL g3816 ( 
.A(n_3513),
.B(n_3217),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3453),
.B(n_3185),
.Y(n_3817)
);

NAND2xp33_ASAP7_75t_SL g3818 ( 
.A(n_3547),
.B(n_3259),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_SL g3819 ( 
.A(n_3513),
.B(n_2925),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_SL g3820 ( 
.A(n_3515),
.B(n_2925),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_SL g3821 ( 
.A(n_3515),
.B(n_2925),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_SL g3822 ( 
.A(n_3553),
.B(n_2979),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_SL g3823 ( 
.A(n_3553),
.B(n_2979),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_3558),
.B(n_2979),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_SL g3825 ( 
.A(n_3558),
.B(n_2979),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_SL g3826 ( 
.A(n_3539),
.B(n_3356),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3456),
.B(n_3229),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3480),
.B(n_3495),
.Y(n_3828)
);

NOR2xp33_ASAP7_75t_L g3829 ( 
.A(n_3442),
.B(n_3636),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_SL g3830 ( 
.A(n_3539),
.B(n_3370),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_SL g3831 ( 
.A(n_3551),
.B(n_3369),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_SL g3832 ( 
.A(n_3551),
.B(n_3559),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_SL g3833 ( 
.A(n_3559),
.B(n_3312),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_SL g3834 ( 
.A(n_3563),
.B(n_3316),
.Y(n_3834)
);

NAND2xp33_ASAP7_75t_SL g3835 ( 
.A(n_3561),
.B(n_3264),
.Y(n_3835)
);

NAND2xp33_ASAP7_75t_SL g3836 ( 
.A(n_3561),
.B(n_3282),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3458),
.B(n_3157),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_SL g3838 ( 
.A(n_3563),
.B(n_3318),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3467),
.B(n_3158),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_SL g3840 ( 
.A(n_3563),
.B(n_3573),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_SL g3841 ( 
.A(n_3563),
.B(n_3326),
.Y(n_3841)
);

NAND2xp33_ASAP7_75t_SL g3842 ( 
.A(n_3561),
.B(n_3046),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_SL g3843 ( 
.A(n_3573),
.B(n_3398),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_SL g3844 ( 
.A(n_3573),
.B(n_3347),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_SL g3845 ( 
.A(n_3573),
.B(n_3256),
.Y(n_3845)
);

NAND2xp33_ASAP7_75t_SL g3846 ( 
.A(n_3568),
.B(n_2993),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_SL g3847 ( 
.A(n_3412),
.B(n_3220),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3471),
.B(n_3115),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3474),
.B(n_3191),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_SL g3850 ( 
.A(n_3514),
.B(n_2600),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3476),
.B(n_3197),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_SL g3852 ( 
.A(n_3514),
.B(n_2600),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_SL g3853 ( 
.A(n_3568),
.B(n_2600),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_SL g3854 ( 
.A(n_3568),
.B(n_2637),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_SL g3855 ( 
.A(n_3655),
.B(n_2637),
.Y(n_3855)
);

NAND2xp33_ASAP7_75t_SL g3856 ( 
.A(n_3655),
.B(n_2993),
.Y(n_3856)
);

NAND2xp33_ASAP7_75t_SL g3857 ( 
.A(n_3655),
.B(n_3216),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_SL g3858 ( 
.A(n_3586),
.B(n_2637),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_SL g3859 ( 
.A(n_3586),
.B(n_2637),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_SL g3860 ( 
.A(n_3489),
.B(n_3283),
.Y(n_3860)
);

NAND2xp33_ASAP7_75t_SL g3861 ( 
.A(n_3446),
.B(n_2710),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3486),
.B(n_3333),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_SL g3863 ( 
.A(n_3430),
.B(n_3290),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_SL g3864 ( 
.A(n_3430),
.B(n_2861),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_SL g3865 ( 
.A(n_3438),
.B(n_2861),
.Y(n_3865)
);

NAND2xp33_ASAP7_75t_SL g3866 ( 
.A(n_3446),
.B(n_2710),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_SL g3867 ( 
.A(n_3438),
.B(n_3500),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_SL g3868 ( 
.A(n_3593),
.B(n_2944),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_SL g3869 ( 
.A(n_3509),
.B(n_3538),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_SL g3870 ( 
.A(n_3658),
.B(n_2944),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3594),
.B(n_2981),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_SL g3872 ( 
.A(n_3594),
.B(n_2981),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_SL g3873 ( 
.A(n_3519),
.B(n_3520),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_SL g3874 ( 
.A(n_3519),
.B(n_2992),
.Y(n_3874)
);

NAND2xp33_ASAP7_75t_SL g3875 ( 
.A(n_3455),
.B(n_2735),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_SL g3876 ( 
.A(n_3520),
.B(n_2992),
.Y(n_3876)
);

NAND2xp33_ASAP7_75t_SL g3877 ( 
.A(n_3455),
.B(n_2735),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_3490),
.B(n_3340),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_SL g3879 ( 
.A(n_3520),
.B(n_2996),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_SL g3880 ( 
.A(n_3483),
.B(n_2996),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_SL g3881 ( 
.A(n_3483),
.B(n_3013),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_SL g3882 ( 
.A(n_3507),
.B(n_3013),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3534),
.B(n_1030),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3516),
.B(n_3349),
.Y(n_3884)
);

NAND2xp33_ASAP7_75t_SL g3885 ( 
.A(n_3595),
.B(n_2758),
.Y(n_3885)
);

NAND2xp33_ASAP7_75t_SL g3886 ( 
.A(n_3601),
.B(n_2758),
.Y(n_3886)
);

NAND2xp33_ASAP7_75t_SL g3887 ( 
.A(n_3440),
.B(n_3373),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3517),
.B(n_3360),
.Y(n_3888)
);

AND2x2_ASAP7_75t_L g3889 ( 
.A(n_3523),
.B(n_1094),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_SL g3890 ( 
.A(n_3507),
.B(n_3269),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_SL g3891 ( 
.A(n_3511),
.B(n_3308),
.Y(n_3891)
);

AND2x4_ASAP7_75t_L g3892 ( 
.A(n_3511),
.B(n_3179),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_3552),
.B(n_3308),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_SL g3894 ( 
.A(n_3383),
.B(n_2980),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_SL g3895 ( 
.A(n_3383),
.B(n_2980),
.Y(n_3895)
);

NAND2xp33_ASAP7_75t_SL g3896 ( 
.A(n_3451),
.B(n_3395),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_SL g3897 ( 
.A(n_3600),
.B(n_3222),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3529),
.B(n_1094),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_SL g3899 ( 
.A(n_3600),
.B(n_3222),
.Y(n_3899)
);

NAND2xp33_ASAP7_75t_SL g3900 ( 
.A(n_3395),
.B(n_3288),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_SL g3901 ( 
.A(n_3432),
.B(n_3344),
.Y(n_3901)
);

NAND2xp33_ASAP7_75t_R g3902 ( 
.A(n_3399),
.B(n_2281),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3537),
.B(n_3541),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3549),
.B(n_3564),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_SL g3905 ( 
.A(n_3621),
.B(n_3358),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_SL g3906 ( 
.A(n_3560),
.B(n_3367),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_SL g3907 ( 
.A(n_3492),
.B(n_2860),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_SL g3908 ( 
.A(n_3562),
.B(n_2881),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_SL g3909 ( 
.A(n_3477),
.B(n_2881),
.Y(n_3909)
);

OAI22xp5_ASAP7_75t_L g3910 ( 
.A1(n_3667),
.A2(n_3414),
.B1(n_3454),
.B2(n_3632),
.Y(n_3910)
);

INVx1_ASAP7_75t_SL g3911 ( 
.A(n_3798),
.Y(n_3911)
);

OAI22xp5_ASAP7_75t_SL g3912 ( 
.A1(n_3829),
.A2(n_3442),
.B1(n_3436),
.B2(n_3397),
.Y(n_3912)
);

AND2x4_ASAP7_75t_L g3913 ( 
.A(n_3777),
.B(n_3632),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_SL g3914 ( 
.A(n_3756),
.B(n_3399),
.Y(n_3914)
);

AND2x2_ASAP7_75t_L g3915 ( 
.A(n_3739),
.B(n_3565),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3903),
.Y(n_3916)
);

BUFx6f_ASAP7_75t_L g3917 ( 
.A(n_3694),
.Y(n_3917)
);

AOI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_3893),
.A2(n_3764),
.B(n_3666),
.Y(n_3918)
);

AOI21xp5_ASAP7_75t_L g3919 ( 
.A1(n_3666),
.A2(n_3651),
.B(n_3439),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3904),
.Y(n_3920)
);

AOI21xp5_ASAP7_75t_L g3921 ( 
.A1(n_3693),
.A2(n_3901),
.B(n_3671),
.Y(n_3921)
);

OAI22xp5_ASAP7_75t_L g3922 ( 
.A1(n_3667),
.A2(n_3454),
.B1(n_3632),
.B2(n_3609),
.Y(n_3922)
);

INVx6_ASAP7_75t_L g3923 ( 
.A(n_3680),
.Y(n_3923)
);

INVxp67_ASAP7_75t_L g3924 ( 
.A(n_3718),
.Y(n_3924)
);

HB1xp67_ASAP7_75t_L g3925 ( 
.A(n_3736),
.Y(n_3925)
);

BUFx2_ASAP7_75t_L g3926 ( 
.A(n_3712),
.Y(n_3926)
);

OAI22xp5_ASAP7_75t_L g3927 ( 
.A1(n_3759),
.A2(n_3468),
.B1(n_3606),
.B2(n_3477),
.Y(n_3927)
);

AND2x4_ASAP7_75t_L g3928 ( 
.A(n_3777),
.B(n_3449),
.Y(n_3928)
);

AOI21xp5_ASAP7_75t_L g3929 ( 
.A1(n_3901),
.A2(n_3671),
.B(n_3886),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3669),
.B(n_3572),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3725),
.B(n_3576),
.Y(n_3931)
);

O2A1O1Ixp33_ASAP7_75t_L g3932 ( 
.A1(n_3683),
.A2(n_3686),
.B(n_3685),
.C(n_3675),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3772),
.Y(n_3933)
);

INVxp67_ASAP7_75t_SL g3934 ( 
.A(n_3867),
.Y(n_3934)
);

INVx4_ASAP7_75t_L g3935 ( 
.A(n_3763),
.Y(n_3935)
);

AND2x6_ASAP7_75t_L g3936 ( 
.A(n_3674),
.B(n_3546),
.Y(n_3936)
);

CKINVDCx20_ASAP7_75t_R g3937 ( 
.A(n_3676),
.Y(n_3937)
);

INVx2_ASAP7_75t_L g3938 ( 
.A(n_3781),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3783),
.Y(n_3939)
);

AND2x4_ASAP7_75t_L g3940 ( 
.A(n_3777),
.B(n_3450),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3663),
.B(n_3588),
.Y(n_3941)
);

BUFx3_ASAP7_75t_L g3942 ( 
.A(n_3828),
.Y(n_3942)
);

BUFx2_ASAP7_75t_L g3943 ( 
.A(n_3715),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3665),
.B(n_3612),
.Y(n_3944)
);

HB1xp67_ASAP7_75t_L g3945 ( 
.A(n_3749),
.Y(n_3945)
);

AOI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_3900),
.A2(n_3439),
.B(n_3626),
.Y(n_3946)
);

BUFx8_ASAP7_75t_SL g3947 ( 
.A(n_3716),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3804),
.Y(n_3948)
);

INVx2_ASAP7_75t_SL g3949 ( 
.A(n_3721),
.Y(n_3949)
);

NOR2xp33_ASAP7_75t_L g3950 ( 
.A(n_3713),
.B(n_3656),
.Y(n_3950)
);

AOI22xp33_ASAP7_75t_L g3951 ( 
.A1(n_3690),
.A2(n_3409),
.B1(n_3417),
.B2(n_3403),
.Y(n_3951)
);

BUFx6f_ASAP7_75t_L g3952 ( 
.A(n_3694),
.Y(n_3952)
);

BUFx2_ASAP7_75t_SL g3953 ( 
.A(n_3677),
.Y(n_3953)
);

NOR2xp33_ASAP7_75t_L g3954 ( 
.A(n_3752),
.B(n_3647),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_SL g3955 ( 
.A(n_3682),
.B(n_3629),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3758),
.B(n_3617),
.Y(n_3956)
);

BUFx2_ASAP7_75t_L g3957 ( 
.A(n_3691),
.Y(n_3957)
);

OR2x6_ASAP7_75t_L g3958 ( 
.A(n_3738),
.B(n_3418),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3806),
.Y(n_3959)
);

O2A1O1Ixp33_ASAP7_75t_L g3960 ( 
.A1(n_3675),
.A2(n_3548),
.B(n_921),
.C(n_937),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3730),
.B(n_3732),
.Y(n_3961)
);

BUFx6f_ASAP7_75t_L g3962 ( 
.A(n_3694),
.Y(n_3962)
);

INVx3_ASAP7_75t_L g3963 ( 
.A(n_3705),
.Y(n_3963)
);

BUFx5_ASAP7_75t_L g3964 ( 
.A(n_3705),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3862),
.Y(n_3965)
);

INVx1_ASAP7_75t_SL g3966 ( 
.A(n_3800),
.Y(n_3966)
);

CKINVDCx8_ASAP7_75t_R g3967 ( 
.A(n_3892),
.Y(n_3967)
);

CKINVDCx5p33_ASAP7_75t_R g3968 ( 
.A(n_3883),
.Y(n_3968)
);

BUFx6f_ASAP7_75t_L g3969 ( 
.A(n_3705),
.Y(n_3969)
);

INVx2_ASAP7_75t_L g3970 ( 
.A(n_3878),
.Y(n_3970)
);

BUFx12f_ASAP7_75t_L g3971 ( 
.A(n_3814),
.Y(n_3971)
);

BUFx6f_ASAP7_75t_L g3972 ( 
.A(n_3706),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3731),
.A2(n_3652),
.B(n_3598),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3813),
.A2(n_3598),
.B(n_3645),
.Y(n_3974)
);

CKINVDCx8_ASAP7_75t_R g3975 ( 
.A(n_3892),
.Y(n_3975)
);

AOI21x1_ASAP7_75t_L g3976 ( 
.A1(n_3860),
.A2(n_3899),
.B(n_3897),
.Y(n_3976)
);

NAND2x1p5_ASAP7_75t_L g3977 ( 
.A(n_3740),
.B(n_3469),
.Y(n_3977)
);

INVx4_ASAP7_75t_L g3978 ( 
.A(n_3706),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3744),
.B(n_3619),
.Y(n_3979)
);

INVx2_ASAP7_75t_SL g3980 ( 
.A(n_3708),
.Y(n_3980)
);

O2A1O1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_3664),
.A2(n_921),
.B(n_937),
.C(n_925),
.Y(n_3981)
);

INVx4_ASAP7_75t_L g3982 ( 
.A(n_3706),
.Y(n_3982)
);

OAI22xp33_ASAP7_75t_L g3983 ( 
.A1(n_3701),
.A2(n_3468),
.B1(n_3583),
.B2(n_3645),
.Y(n_3983)
);

CKINVDCx5p33_ASAP7_75t_R g3984 ( 
.A(n_3902),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3884),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3888),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3769),
.Y(n_3987)
);

OAI22x1_ASAP7_75t_L g3988 ( 
.A1(n_3692),
.A2(n_3624),
.B1(n_3634),
.B2(n_3623),
.Y(n_3988)
);

INVxp67_ASAP7_75t_SL g3989 ( 
.A(n_3672),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3770),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3703),
.Y(n_3991)
);

OAI22xp5_ASAP7_75t_L g3992 ( 
.A1(n_3759),
.A2(n_3605),
.B1(n_3660),
.B2(n_3620),
.Y(n_3992)
);

A2O1A1Ixp33_ASAP7_75t_L g3993 ( 
.A1(n_3789),
.A2(n_3638),
.B(n_3644),
.C(n_3639),
.Y(n_3993)
);

BUFx3_ASAP7_75t_L g3994 ( 
.A(n_3697),
.Y(n_3994)
);

O2A1O1Ixp33_ASAP7_75t_SL g3995 ( 
.A1(n_3702),
.A2(n_925),
.B(n_941),
.C(n_939),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3704),
.Y(n_3996)
);

AOI22xp33_ASAP7_75t_L g3997 ( 
.A1(n_3689),
.A2(n_3425),
.B1(n_3431),
.B2(n_3419),
.Y(n_3997)
);

BUFx3_ASAP7_75t_L g3998 ( 
.A(n_3714),
.Y(n_3998)
);

INVx4_ASAP7_75t_L g3999 ( 
.A(n_3714),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_SL g4000 ( 
.A(n_3734),
.B(n_3629),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_3849),
.Y(n_4001)
);

NOR2xp33_ASAP7_75t_L g4002 ( 
.A(n_3724),
.B(n_3613),
.Y(n_4002)
);

AND2x2_ASAP7_75t_SL g4003 ( 
.A(n_3848),
.B(n_3546),
.Y(n_4003)
);

AO21x2_ASAP7_75t_L g4004 ( 
.A1(n_3782),
.A2(n_3585),
.B(n_3583),
.Y(n_4004)
);

AOI21xp5_ASAP7_75t_L g4005 ( 
.A1(n_3818),
.A2(n_3643),
.B(n_3637),
.Y(n_4005)
);

A2O1A1Ixp33_ASAP7_75t_L g4006 ( 
.A1(n_3670),
.A2(n_3661),
.B(n_3650),
.C(n_3502),
.Y(n_4006)
);

OAI22xp5_ASAP7_75t_L g4007 ( 
.A1(n_3664),
.A2(n_3461),
.B1(n_3643),
.B2(n_3637),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3851),
.Y(n_4008)
);

INVx2_ASAP7_75t_L g4009 ( 
.A(n_3827),
.Y(n_4009)
);

OR2x2_ASAP7_75t_L g4010 ( 
.A(n_3728),
.B(n_3518),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3673),
.B(n_3544),
.Y(n_4011)
);

BUFx6f_ASAP7_75t_L g4012 ( 
.A(n_3714),
.Y(n_4012)
);

AND2x2_ASAP7_75t_L g4013 ( 
.A(n_3765),
.B(n_3630),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_SL g4014 ( 
.A(n_3762),
.B(n_3630),
.Y(n_4014)
);

NOR2x1_ASAP7_75t_L g4015 ( 
.A(n_3672),
.B(n_3424),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3709),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3695),
.B(n_3380),
.Y(n_4017)
);

INVx4_ASAP7_75t_L g4018 ( 
.A(n_3720),
.Y(n_4018)
);

O2A1O1Ixp33_ASAP7_75t_L g4019 ( 
.A1(n_3792),
.A2(n_939),
.B(n_942),
.C(n_941),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_L g4020 ( 
.A(n_3699),
.B(n_3381),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3711),
.Y(n_4021)
);

INVx1_ASAP7_75t_SL g4022 ( 
.A(n_3727),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3837),
.Y(n_4023)
);

INVx2_ASAP7_75t_L g4024 ( 
.A(n_3839),
.Y(n_4024)
);

BUFx4f_ASAP7_75t_SL g4025 ( 
.A(n_3745),
.Y(n_4025)
);

INVx1_ASAP7_75t_SL g4026 ( 
.A(n_3717),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3811),
.Y(n_4027)
);

O2A1O1Ixp33_ASAP7_75t_L g4028 ( 
.A1(n_3684),
.A2(n_942),
.B(n_951),
.C(n_950),
.Y(n_4028)
);

AOI21xp5_ASAP7_75t_L g4029 ( 
.A1(n_3835),
.A2(n_3022),
.B(n_3435),
.Y(n_4029)
);

BUFx4f_ASAP7_75t_L g4030 ( 
.A(n_3720),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3766),
.B(n_3387),
.Y(n_4031)
);

AOI22xp33_ASAP7_75t_L g4032 ( 
.A1(n_3687),
.A2(n_3434),
.B1(n_3448),
.B2(n_3437),
.Y(n_4032)
);

BUFx3_ASAP7_75t_L g4033 ( 
.A(n_3720),
.Y(n_4033)
);

INVx4_ASAP7_75t_L g4034 ( 
.A(n_3892),
.Y(n_4034)
);

INVxp67_ASAP7_75t_L g4035 ( 
.A(n_3889),
.Y(n_4035)
);

AND3x1_ASAP7_75t_SL g4036 ( 
.A(n_3668),
.B(n_950),
.C(n_912),
.Y(n_4036)
);

BUFx2_ASAP7_75t_L g4037 ( 
.A(n_3761),
.Y(n_4037)
);

NAND2x1p5_ASAP7_75t_L g4038 ( 
.A(n_3743),
.B(n_3469),
.Y(n_4038)
);

INVx4_ASAP7_75t_L g4039 ( 
.A(n_3674),
.Y(n_4039)
);

OR2x6_ASAP7_75t_SL g4040 ( 
.A(n_3768),
.B(n_3535),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3815),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3817),
.Y(n_4042)
);

BUFx2_ASAP7_75t_SL g4043 ( 
.A(n_3700),
.Y(n_4043)
);

AND2x6_ASAP7_75t_L g4044 ( 
.A(n_3674),
.B(n_3688),
.Y(n_4044)
);

INVx2_ASAP7_75t_L g4045 ( 
.A(n_3760),
.Y(n_4045)
);

AND2x2_ASAP7_75t_L g4046 ( 
.A(n_3898),
.B(n_951),
.Y(n_4046)
);

AND2x2_ASAP7_75t_L g4047 ( 
.A(n_3735),
.B(n_953),
.Y(n_4047)
);

A2O1A1Ixp33_ASAP7_75t_SL g4048 ( 
.A1(n_3733),
.A2(n_960),
.B(n_965),
.C(n_953),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3786),
.Y(n_4049)
);

AOI22xp5_ASAP7_75t_L g4050 ( 
.A1(n_3678),
.A2(n_3613),
.B1(n_3592),
.B2(n_3532),
.Y(n_4050)
);

A2O1A1Ixp33_ASAP7_75t_L g4051 ( 
.A1(n_3662),
.A2(n_3575),
.B(n_3592),
.C(n_3532),
.Y(n_4051)
);

A2O1A1Ixp33_ASAP7_75t_L g4052 ( 
.A1(n_3662),
.A2(n_965),
.B(n_973),
.C(n_960),
.Y(n_4052)
);

AOI21xp5_ASAP7_75t_L g4053 ( 
.A1(n_3836),
.A2(n_3022),
.B(n_3435),
.Y(n_4053)
);

A2O1A1Ixp33_ASAP7_75t_L g4054 ( 
.A1(n_3679),
.A2(n_974),
.B(n_976),
.C(n_973),
.Y(n_4054)
);

NOR2xp67_ASAP7_75t_L g4055 ( 
.A(n_3750),
.B(n_1505),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3832),
.Y(n_4056)
);

AOI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_3896),
.A2(n_3535),
.B1(n_1119),
.B2(n_1094),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3780),
.B(n_974),
.Y(n_4058)
);

INVx5_ASAP7_75t_L g4059 ( 
.A(n_3688),
.Y(n_4059)
);

AOI222xp33_ASAP7_75t_L g4060 ( 
.A1(n_3754),
.A2(n_988),
.B1(n_983),
.B2(n_992),
.C1(n_986),
.C2(n_976),
.Y(n_4060)
);

INVx5_ASAP7_75t_L g4061 ( 
.A(n_3688),
.Y(n_4061)
);

O2A1O1Ixp33_ASAP7_75t_L g4062 ( 
.A1(n_3831),
.A2(n_986),
.B(n_992),
.C(n_983),
.Y(n_4062)
);

BUFx6f_ASAP7_75t_L g4063 ( 
.A(n_3746),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3773),
.B(n_3393),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3833),
.Y(n_4065)
);

OAI22xp5_ASAP7_75t_L g4066 ( 
.A1(n_3909),
.A2(n_3574),
.B1(n_3578),
.B2(n_994),
.Y(n_4066)
);

BUFx6f_ASAP7_75t_L g4067 ( 
.A(n_3746),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_3830),
.Y(n_4068)
);

AOI21xp5_ASAP7_75t_L g4069 ( 
.A1(n_3808),
.A2(n_3036),
.B(n_2414),
.Y(n_4069)
);

A2O1A1Ixp33_ASAP7_75t_L g4070 ( 
.A1(n_3681),
.A2(n_994),
.B(n_995),
.C(n_988),
.Y(n_4070)
);

OAI22xp5_ASAP7_75t_L g4071 ( 
.A1(n_3909),
.A2(n_996),
.B1(n_1002),
.B2(n_995),
.Y(n_4071)
);

AOI22xp33_ASAP7_75t_L g4072 ( 
.A1(n_3908),
.A2(n_3491),
.B1(n_3503),
.B2(n_3487),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_3775),
.B(n_3504),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3787),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3778),
.B(n_3510),
.Y(n_4075)
);

XOR2x2_ASAP7_75t_L g4076 ( 
.A(n_3771),
.B(n_996),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_SL g4077 ( 
.A(n_3857),
.B(n_3625),
.Y(n_4077)
);

OAI21x1_ASAP7_75t_L g4078 ( 
.A1(n_3799),
.A2(n_2286),
.B(n_3642),
.Y(n_4078)
);

BUFx2_ASAP7_75t_L g4079 ( 
.A(n_3805),
.Y(n_4079)
);

A2O1A1Ixp33_ASAP7_75t_L g4080 ( 
.A1(n_3861),
.A2(n_3875),
.B(n_3877),
.C(n_3866),
.Y(n_4080)
);

INVxp67_ASAP7_75t_L g4081 ( 
.A(n_3801),
.Y(n_4081)
);

BUFx2_ASAP7_75t_SL g4082 ( 
.A(n_3891),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3790),
.Y(n_4083)
);

AOI22xp5_ASAP7_75t_L g4084 ( 
.A1(n_3737),
.A2(n_1119),
.B1(n_1094),
.B2(n_3625),
.Y(n_4084)
);

O2A1O1Ixp33_ASAP7_75t_L g4085 ( 
.A1(n_3890),
.A2(n_3847),
.B(n_1016),
.C(n_1025),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3784),
.Y(n_4086)
);

AOI21xp5_ASAP7_75t_L g4087 ( 
.A1(n_3897),
.A2(n_3036),
.B(n_2417),
.Y(n_4087)
);

A2O1A1Ixp33_ASAP7_75t_L g4088 ( 
.A1(n_3907),
.A2(n_1016),
.B(n_1025),
.C(n_1002),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_3894),
.B(n_1026),
.Y(n_4089)
);

AOI21xp5_ASAP7_75t_L g4090 ( 
.A1(n_3899),
.A2(n_2417),
.B(n_2391),
.Y(n_4090)
);

NAND2x1p5_ASAP7_75t_L g4091 ( 
.A(n_3748),
.B(n_3512),
.Y(n_4091)
);

INVx4_ASAP7_75t_L g4092 ( 
.A(n_3746),
.Y(n_4092)
);

AND2x2_ASAP7_75t_L g4093 ( 
.A(n_3895),
.B(n_1026),
.Y(n_4093)
);

AOI21xp5_ASAP7_75t_L g4094 ( 
.A1(n_3776),
.A2(n_2421),
.B(n_2417),
.Y(n_4094)
);

BUFx6f_ASAP7_75t_L g4095 ( 
.A(n_3774),
.Y(n_4095)
);

INVx2_ASAP7_75t_L g4096 ( 
.A(n_3874),
.Y(n_4096)
);

A2O1A1Ixp33_ASAP7_75t_L g4097 ( 
.A1(n_3907),
.A2(n_1043),
.B(n_1044),
.C(n_1031),
.Y(n_4097)
);

AOI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3908),
.A2(n_1119),
.B1(n_944),
.B2(n_947),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3753),
.B(n_3526),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_SL g4100 ( 
.A(n_3767),
.B(n_3741),
.Y(n_4100)
);

OAI22xp5_ASAP7_75t_L g4101 ( 
.A1(n_3871),
.A2(n_1043),
.B1(n_1044),
.B2(n_1031),
.Y(n_4101)
);

AND2x2_ASAP7_75t_SL g4102 ( 
.A(n_3840),
.B(n_3530),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_3826),
.B(n_3533),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_SL g4104 ( 
.A(n_3742),
.B(n_3536),
.Y(n_4104)
);

INVx2_ASAP7_75t_L g4105 ( 
.A(n_3864),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_3723),
.Y(n_4106)
);

INVx1_ASAP7_75t_SL g4107 ( 
.A(n_3729),
.Y(n_4107)
);

BUFx6f_ASAP7_75t_L g4108 ( 
.A(n_3803),
.Y(n_4108)
);

INVx2_ASAP7_75t_L g4109 ( 
.A(n_3865),
.Y(n_4109)
);

OAI22xp33_ASAP7_75t_L g4110 ( 
.A1(n_3707),
.A2(n_1125),
.B1(n_1083),
.B2(n_1052),
.Y(n_4110)
);

AOI22xp5_ASAP7_75t_L g4111 ( 
.A1(n_3696),
.A2(n_3872),
.B1(n_3751),
.B2(n_3842),
.Y(n_4111)
);

AOI21xp5_ASAP7_75t_L g4112 ( 
.A1(n_3779),
.A2(n_2443),
.B(n_2421),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_3863),
.Y(n_4113)
);

AND2x4_ASAP7_75t_SL g4114 ( 
.A(n_3698),
.B(n_3542),
.Y(n_4114)
);

INVx2_ASAP7_75t_L g4115 ( 
.A(n_3726),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3793),
.Y(n_4116)
);

INVx5_ASAP7_75t_L g4117 ( 
.A(n_3747),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3816),
.B(n_3540),
.Y(n_4118)
);

NOR2xp33_ASAP7_75t_L g4119 ( 
.A(n_3710),
.B(n_940),
.Y(n_4119)
);

CKINVDCx16_ASAP7_75t_R g4120 ( 
.A(n_3846),
.Y(n_4120)
);

A2O1A1Ixp33_ASAP7_75t_L g4121 ( 
.A1(n_3755),
.A2(n_1052),
.B(n_1055),
.C(n_1045),
.Y(n_4121)
);

INVx3_ASAP7_75t_L g4122 ( 
.A(n_3887),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3794),
.Y(n_4123)
);

INVx2_ASAP7_75t_SL g4124 ( 
.A(n_3802),
.Y(n_4124)
);

CKINVDCx8_ASAP7_75t_R g4125 ( 
.A(n_3856),
.Y(n_4125)
);

BUFx3_ASAP7_75t_L g4126 ( 
.A(n_3807),
.Y(n_4126)
);

BUFx6f_ASAP7_75t_L g4127 ( 
.A(n_3881),
.Y(n_4127)
);

INVx3_ASAP7_75t_L g4128 ( 
.A(n_3785),
.Y(n_4128)
);

INVx5_ASAP7_75t_L g4129 ( 
.A(n_3788),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3873),
.Y(n_4130)
);

AND2x2_ASAP7_75t_L g4131 ( 
.A(n_3868),
.B(n_1045),
.Y(n_4131)
);

INVx2_ASAP7_75t_L g4132 ( 
.A(n_3850),
.Y(n_4132)
);

AOI222xp33_ASAP7_75t_L g4133 ( 
.A1(n_3906),
.A2(n_1067),
.B1(n_1057),
.B2(n_1070),
.C1(n_1061),
.C2(n_1055),
.Y(n_4133)
);

INVx1_ASAP7_75t_SL g4134 ( 
.A(n_3882),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_3869),
.B(n_3577),
.Y(n_4135)
);

HB1xp67_ASAP7_75t_L g4136 ( 
.A(n_3906),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3852),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_3858),
.Y(n_4138)
);

BUFx4f_ASAP7_75t_L g4139 ( 
.A(n_3843),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_3859),
.Y(n_4140)
);

BUFx4_ASAP7_75t_SL g4141 ( 
.A(n_3757),
.Y(n_4141)
);

OR2x6_ASAP7_75t_L g4142 ( 
.A(n_3845),
.B(n_3582),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3791),
.B(n_3590),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4056),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_SL g4145 ( 
.A(n_4122),
.B(n_3719),
.Y(n_4145)
);

OA21x2_ASAP7_75t_L g4146 ( 
.A1(n_3921),
.A2(n_3905),
.B(n_3722),
.Y(n_4146)
);

BUFx12f_ASAP7_75t_L g4147 ( 
.A(n_3968),
.Y(n_4147)
);

A2O1A1Ixp33_ASAP7_75t_L g4148 ( 
.A1(n_3918),
.A2(n_1061),
.B(n_1067),
.C(n_1057),
.Y(n_4148)
);

AOI21xp33_ASAP7_75t_L g4149 ( 
.A1(n_4085),
.A2(n_3844),
.B(n_3838),
.Y(n_4149)
);

O2A1O1Ixp33_ASAP7_75t_L g4150 ( 
.A1(n_4070),
.A2(n_1080),
.B(n_1083),
.C(n_1070),
.Y(n_4150)
);

AND2x2_ASAP7_75t_SL g4151 ( 
.A(n_4120),
.B(n_1080),
.Y(n_4151)
);

OAI21x1_ASAP7_75t_L g4152 ( 
.A1(n_3976),
.A2(n_3810),
.B(n_3809),
.Y(n_4152)
);

AO31x2_ASAP7_75t_L g4153 ( 
.A1(n_3927),
.A2(n_3602),
.A3(n_3607),
.B(n_3596),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3945),
.B(n_3905),
.Y(n_4154)
);

AOI21xp5_ASAP7_75t_L g4155 ( 
.A1(n_4080),
.A2(n_3885),
.B(n_3812),
.Y(n_4155)
);

AOI22xp5_ASAP7_75t_L g4156 ( 
.A1(n_3910),
.A2(n_3796),
.B1(n_3797),
.B2(n_3795),
.Y(n_4156)
);

OAI21x1_ASAP7_75t_L g4157 ( 
.A1(n_3929),
.A2(n_3841),
.B(n_3834),
.Y(n_4157)
);

OAI22xp5_ASAP7_75t_L g4158 ( 
.A1(n_3957),
.A2(n_3819),
.B1(n_3821),
.B2(n_3820),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_3925),
.B(n_1084),
.Y(n_4159)
);

BUFx6f_ASAP7_75t_L g4160 ( 
.A(n_4125),
.Y(n_4160)
);

O2A1O1Ixp33_ASAP7_75t_L g4161 ( 
.A1(n_3932),
.A2(n_1086),
.B(n_1091),
.C(n_1084),
.Y(n_4161)
);

BUFx3_ASAP7_75t_L g4162 ( 
.A(n_3942),
.Y(n_4162)
);

OAI22xp33_ASAP7_75t_L g4163 ( 
.A1(n_3922),
.A2(n_3870),
.B1(n_3880),
.B2(n_1091),
.Y(n_4163)
);

OAI21x1_ASAP7_75t_L g4164 ( 
.A1(n_3973),
.A2(n_3823),
.B(n_3822),
.Y(n_4164)
);

A2O1A1Ixp33_ASAP7_75t_L g4165 ( 
.A1(n_4057),
.A2(n_1106),
.B(n_1110),
.C(n_1086),
.Y(n_4165)
);

AO21x2_ASAP7_75t_L g4166 ( 
.A1(n_4118),
.A2(n_3879),
.B(n_3876),
.Y(n_4166)
);

BUFx2_ASAP7_75t_L g4167 ( 
.A(n_3935),
.Y(n_4167)
);

AO31x2_ASAP7_75t_L g4168 ( 
.A1(n_3946),
.A2(n_3646),
.A3(n_3635),
.B(n_3366),
.Y(n_4168)
);

AOI221x1_ASAP7_75t_L g4169 ( 
.A1(n_3993),
.A2(n_1114),
.B1(n_1115),
.B2(n_1110),
.C(n_1106),
.Y(n_4169)
);

AOI21xp5_ASAP7_75t_L g4170 ( 
.A1(n_4100),
.A2(n_3854),
.B(n_3853),
.Y(n_4170)
);

INVxp67_ASAP7_75t_L g4171 ( 
.A(n_3994),
.Y(n_4171)
);

OAI21x1_ASAP7_75t_L g4172 ( 
.A1(n_4078),
.A2(n_3919),
.B(n_4029),
.Y(n_4172)
);

INVx2_ASAP7_75t_L g4173 ( 
.A(n_4009),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4041),
.Y(n_4174)
);

AOI21xp5_ASAP7_75t_L g4175 ( 
.A1(n_3974),
.A2(n_3855),
.B(n_3825),
.Y(n_4175)
);

AOI22xp5_ASAP7_75t_L g4176 ( 
.A1(n_3992),
.A2(n_1115),
.B1(n_1120),
.B2(n_1114),
.Y(n_4176)
);

INVx4_ASAP7_75t_SL g4177 ( 
.A(n_3912),
.Y(n_4177)
);

A2O1A1Ixp33_ASAP7_75t_L g4178 ( 
.A1(n_4098),
.A2(n_1122),
.B(n_1126),
.C(n_1120),
.Y(n_4178)
);

AOI21x1_ASAP7_75t_L g4179 ( 
.A1(n_4077),
.A2(n_3824),
.B(n_1514),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4023),
.Y(n_4180)
);

NOR4xp25_ASAP7_75t_L g4181 ( 
.A(n_3981),
.B(n_1122),
.C(n_1126),
.D(n_1512),
.Y(n_4181)
);

NOR2x1_ASAP7_75t_SL g4182 ( 
.A(n_4117),
.B(n_879),
.Y(n_4182)
);

OAI22xp5_ASAP7_75t_L g4183 ( 
.A1(n_3953),
.A2(n_967),
.B1(n_1021),
.B2(n_879),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_4049),
.B(n_967),
.Y(n_4184)
);

OAI22xp5_ASAP7_75t_L g4185 ( 
.A1(n_3953),
.A2(n_1021),
.B1(n_1046),
.B2(n_967),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4024),
.Y(n_4186)
);

CKINVDCx20_ASAP7_75t_R g4187 ( 
.A(n_3947),
.Y(n_4187)
);

O2A1O1Ixp33_ASAP7_75t_L g4188 ( 
.A1(n_4054),
.A2(n_1515),
.B(n_1516),
.C(n_1888),
.Y(n_4188)
);

CKINVDCx5p33_ASAP7_75t_R g4189 ( 
.A(n_3971),
.Y(n_4189)
);

AOI221x1_ASAP7_75t_L g4190 ( 
.A1(n_3988),
.A2(n_1542),
.B1(n_1046),
.B2(n_1063),
.C(n_1021),
.Y(n_4190)
);

OAI21x1_ASAP7_75t_L g4191 ( 
.A1(n_4053),
.A2(n_3648),
.B(n_2263),
.Y(n_4191)
);

OR2x2_ASAP7_75t_L g4192 ( 
.A(n_3980),
.B(n_1415),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4027),
.Y(n_4193)
);

AOI21xp5_ASAP7_75t_L g4194 ( 
.A1(n_4117),
.A2(n_2275),
.B(n_2257),
.Y(n_4194)
);

OAI21x1_ASAP7_75t_L g4195 ( 
.A1(n_4122),
.A2(n_2263),
.B(n_2281),
.Y(n_4195)
);

INVx3_ASAP7_75t_SL g4196 ( 
.A(n_3937),
.Y(n_4196)
);

A2O1A1Ixp33_ASAP7_75t_L g4197 ( 
.A1(n_3954),
.A2(n_957),
.B(n_958),
.C(n_948),
.Y(n_4197)
);

A2O1A1Ixp33_ASAP7_75t_L g4198 ( 
.A1(n_4084),
.A2(n_962),
.B(n_963),
.C(n_955),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_L g4199 ( 
.A(n_3941),
.B(n_967),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4042),
.Y(n_4200)
);

NAND3xp33_ASAP7_75t_L g4201 ( 
.A(n_4060),
.B(n_1021),
.C(n_967),
.Y(n_4201)
);

OAI21x1_ASAP7_75t_L g4202 ( 
.A1(n_4087),
.A2(n_2263),
.B(n_2281),
.Y(n_4202)
);

AO31x2_ASAP7_75t_L g4203 ( 
.A1(n_4007),
.A2(n_3368),
.A3(n_3362),
.B(n_2793),
.Y(n_4203)
);

O2A1O1Ixp33_ASAP7_75t_L g4204 ( 
.A1(n_4052),
.A2(n_4097),
.B(n_4088),
.C(n_4071),
.Y(n_4204)
);

AOI21xp5_ASAP7_75t_L g4205 ( 
.A1(n_4117),
.A2(n_2275),
.B(n_2257),
.Y(n_4205)
);

AND2x2_ASAP7_75t_L g4206 ( 
.A(n_3923),
.B(n_967),
.Y(n_4206)
);

A2O1A1Ixp33_ASAP7_75t_L g4207 ( 
.A1(n_4119),
.A2(n_969),
.B(n_970),
.C(n_959),
.Y(n_4207)
);

INVx3_ASAP7_75t_L g4208 ( 
.A(n_3923),
.Y(n_4208)
);

AO22x2_ASAP7_75t_L g4209 ( 
.A1(n_3916),
.A2(n_3002),
.B1(n_2989),
.B2(n_2795),
.Y(n_4209)
);

INVxp67_ASAP7_75t_SL g4210 ( 
.A(n_4136),
.Y(n_4210)
);

BUFx2_ASAP7_75t_SL g4211 ( 
.A(n_3966),
.Y(n_4211)
);

NAND3xp33_ASAP7_75t_L g4212 ( 
.A(n_4133),
.B(n_1046),
.C(n_1021),
.Y(n_4212)
);

A2O1A1Ixp33_ASAP7_75t_L g4213 ( 
.A1(n_3960),
.A2(n_978),
.B(n_979),
.C(n_966),
.Y(n_4213)
);

AOI21x1_ASAP7_75t_L g4214 ( 
.A1(n_3943),
.A2(n_1542),
.B(n_1421),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_3944),
.B(n_1021),
.Y(n_4215)
);

OAI21x1_ASAP7_75t_L g4216 ( 
.A1(n_4005),
.A2(n_2285),
.B(n_2283),
.Y(n_4216)
);

INVx2_ASAP7_75t_SL g4217 ( 
.A(n_4010),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_3956),
.B(n_1046),
.Y(n_4218)
);

AO21x1_ASAP7_75t_L g4219 ( 
.A1(n_3983),
.A2(n_1119),
.B(n_1418),
.Y(n_4219)
);

INVx2_ASAP7_75t_L g4220 ( 
.A(n_4001),
.Y(n_4220)
);

AO31x2_ASAP7_75t_L g4221 ( 
.A1(n_4116),
.A2(n_2796),
.A3(n_2824),
.B(n_2791),
.Y(n_4221)
);

AO31x2_ASAP7_75t_L g4222 ( 
.A1(n_4123),
.A2(n_2884),
.A3(n_2885),
.B(n_2826),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_3961),
.B(n_1046),
.Y(n_4223)
);

NOR2xp33_ASAP7_75t_SL g4224 ( 
.A(n_3984),
.B(n_4022),
.Y(n_4224)
);

NAND3x1_ASAP7_75t_L g4225 ( 
.A(n_4002),
.B(n_2443),
.C(n_2421),
.Y(n_4225)
);

AO31x2_ASAP7_75t_L g4226 ( 
.A1(n_4132),
.A2(n_2912),
.A3(n_2922),
.B(n_2905),
.Y(n_4226)
);

OAI21x1_ASAP7_75t_L g4227 ( 
.A1(n_4090),
.A2(n_4128),
.B(n_4015),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4008),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3920),
.Y(n_4229)
);

OAI21x1_ASAP7_75t_L g4230 ( 
.A1(n_4128),
.A2(n_2285),
.B(n_2283),
.Y(n_4230)
);

OAI21xp5_ASAP7_75t_L g4231 ( 
.A1(n_4121),
.A2(n_980),
.B(n_977),
.Y(n_4231)
);

OAI21x1_ASAP7_75t_L g4232 ( 
.A1(n_4000),
.A2(n_2285),
.B(n_2283),
.Y(n_4232)
);

AOI21xp5_ASAP7_75t_L g4233 ( 
.A1(n_4129),
.A2(n_2292),
.B(n_2443),
.Y(n_4233)
);

AOI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_4129),
.A2(n_2292),
.B(n_2447),
.Y(n_4234)
);

OR2x2_ASAP7_75t_L g4235 ( 
.A(n_3915),
.B(n_1418),
.Y(n_4235)
);

OAI21xp5_ASAP7_75t_SL g4236 ( 
.A1(n_3926),
.A2(n_1100),
.B(n_1063),
.Y(n_4236)
);

NOR4xp25_ASAP7_75t_L g4237 ( 
.A(n_4058),
.B(n_1422),
.C(n_1451),
.D(n_1421),
.Y(n_4237)
);

NOR2xp33_ASAP7_75t_L g4238 ( 
.A(n_4040),
.B(n_3),
.Y(n_4238)
);

CKINVDCx5p33_ASAP7_75t_R g4239 ( 
.A(n_3911),
.Y(n_4239)
);

OAI21x1_ASAP7_75t_L g4240 ( 
.A1(n_4069),
.A2(n_2539),
.B(n_2537),
.Y(n_4240)
);

CKINVDCx11_ASAP7_75t_R g4241 ( 
.A(n_3967),
.Y(n_4241)
);

OAI21x1_ASAP7_75t_L g4242 ( 
.A1(n_4104),
.A2(n_2549),
.B(n_2539),
.Y(n_4242)
);

A2O1A1Ixp33_ASAP7_75t_L g4243 ( 
.A1(n_4019),
.A2(n_985),
.B(n_987),
.C(n_981),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_4086),
.B(n_1046),
.Y(n_4244)
);

OAI21xp5_ASAP7_75t_L g4245 ( 
.A1(n_4006),
.A2(n_989),
.B(n_982),
.Y(n_4245)
);

CKINVDCx5p33_ASAP7_75t_R g4246 ( 
.A(n_3924),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_3933),
.Y(n_4247)
);

AO31x2_ASAP7_75t_L g4248 ( 
.A1(n_4138),
.A2(n_2935),
.A3(n_2945),
.B(n_2929),
.Y(n_4248)
);

AO21x2_ASAP7_75t_L g4249 ( 
.A1(n_4099),
.A2(n_1451),
.B(n_1422),
.Y(n_4249)
);

AOI21x1_ASAP7_75t_L g4250 ( 
.A1(n_4079),
.A2(n_1461),
.B(n_1459),
.Y(n_4250)
);

AO21x1_ASAP7_75t_L g4251 ( 
.A1(n_3979),
.A2(n_1461),
.B(n_1459),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_3938),
.Y(n_4252)
);

AOI21xp5_ASAP7_75t_L g4253 ( 
.A1(n_4129),
.A2(n_2459),
.B(n_2447),
.Y(n_4253)
);

A2O1A1Ixp33_ASAP7_75t_L g4254 ( 
.A1(n_4111),
.A2(n_999),
.B(n_1003),
.C(n_990),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_3939),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_3959),
.B(n_1063),
.Y(n_4256)
);

AOI21x1_ASAP7_75t_L g4257 ( 
.A1(n_4089),
.A2(n_1479),
.B(n_1473),
.Y(n_4257)
);

HB1xp67_ASAP7_75t_L g4258 ( 
.A(n_3989),
.Y(n_4258)
);

OR2x6_ASAP7_75t_L g4259 ( 
.A(n_4043),
.B(n_2549),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_4139),
.A2(n_2459),
.B(n_2447),
.Y(n_4260)
);

O2A1O1Ixp33_ASAP7_75t_L g4261 ( 
.A1(n_4048),
.A2(n_2135),
.B(n_1479),
.C(n_1481),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_3987),
.B(n_3990),
.Y(n_4262)
);

O2A1O1Ixp5_ASAP7_75t_SL g4263 ( 
.A1(n_4035),
.A2(n_2512),
.B(n_2528),
.C(n_2499),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_3930),
.B(n_1063),
.Y(n_4264)
);

AOI21xp5_ASAP7_75t_L g4265 ( 
.A1(n_4139),
.A2(n_2512),
.B(n_2499),
.Y(n_4265)
);

A2O1A1Ixp33_ASAP7_75t_L g4266 ( 
.A1(n_4028),
.A2(n_1006),
.B(n_1008),
.C(n_997),
.Y(n_4266)
);

AOI21xp5_ASAP7_75t_SL g4267 ( 
.A1(n_3914),
.A2(n_2555),
.B(n_2553),
.Y(n_4267)
);

AOI22xp33_ASAP7_75t_L g4268 ( 
.A1(n_3951),
.A2(n_2976),
.B1(n_2985),
.B2(n_2947),
.Y(n_4268)
);

OAI21xp5_ASAP7_75t_L g4269 ( 
.A1(n_4055),
.A2(n_1010),
.B(n_1005),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_4074),
.B(n_1063),
.Y(n_4270)
);

OAI21x1_ASAP7_75t_L g4271 ( 
.A1(n_4140),
.A2(n_2555),
.B(n_2553),
.Y(n_4271)
);

OAI21x1_ASAP7_75t_L g4272 ( 
.A1(n_3955),
.A2(n_2561),
.B(n_2560),
.Y(n_4272)
);

O2A1O1Ixp33_ASAP7_75t_SL g4273 ( 
.A1(n_4026),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_3970),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_4083),
.B(n_1063),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_SL g4276 ( 
.A(n_4037),
.B(n_1473),
.Y(n_4276)
);

AOI21xp5_ASAP7_75t_L g4277 ( 
.A1(n_4014),
.A2(n_2512),
.B(n_2499),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_SL g4278 ( 
.A(n_4107),
.B(n_1481),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_3949),
.B(n_1100),
.Y(n_4279)
);

INVx2_ASAP7_75t_SL g4280 ( 
.A(n_4011),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_3948),
.Y(n_4281)
);

BUFx2_ASAP7_75t_L g4282 ( 
.A(n_3935),
.Y(n_4282)
);

NOR2xp33_ASAP7_75t_L g4283 ( 
.A(n_3950),
.B(n_6),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3965),
.Y(n_4284)
);

INVx4_ASAP7_75t_L g4285 ( 
.A(n_4095),
.Y(n_4285)
);

AO22x2_ASAP7_75t_L g4286 ( 
.A1(n_3985),
.A2(n_3986),
.B1(n_4130),
.B2(n_4045),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_3934),
.Y(n_4287)
);

OR2x2_ASAP7_75t_L g4288 ( 
.A(n_3931),
.B(n_1483),
.Y(n_4288)
);

AOI221xp5_ASAP7_75t_L g4289 ( 
.A1(n_4062),
.A2(n_1020),
.B1(n_1022),
.B2(n_1013),
.C(n_1011),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_4065),
.B(n_4013),
.Y(n_4290)
);

OAI21xp5_ASAP7_75t_L g4291 ( 
.A1(n_4076),
.A2(n_4101),
.B(n_4137),
.Y(n_4291)
);

AOI21xp5_ASAP7_75t_L g4292 ( 
.A1(n_4094),
.A2(n_2540),
.B(n_2528),
.Y(n_4292)
);

INVx1_ASAP7_75t_SL g4293 ( 
.A(n_4003),
.Y(n_4293)
);

NOR4xp25_ASAP7_75t_L g4294 ( 
.A(n_4046),
.B(n_4047),
.C(n_4093),
.D(n_4131),
.Y(n_4294)
);

AO21x2_ASAP7_75t_L g4295 ( 
.A1(n_4103),
.A2(n_1501),
.B(n_1483),
.Y(n_4295)
);

AOI22xp5_ASAP7_75t_L g4296 ( 
.A1(n_4036),
.A2(n_4066),
.B1(n_4082),
.B2(n_3958),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4068),
.B(n_1100),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4113),
.B(n_1100),
.Y(n_4298)
);

OAI21x1_ASAP7_75t_L g4299 ( 
.A1(n_4135),
.A2(n_2561),
.B(n_2560),
.Y(n_4299)
);

O2A1O1Ixp33_ASAP7_75t_L g4300 ( 
.A1(n_3995),
.A2(n_1502),
.B(n_1530),
.C(n_1501),
.Y(n_4300)
);

NOR2xp33_ASAP7_75t_SL g4301 ( 
.A(n_3975),
.B(n_2567),
.Y(n_4301)
);

INVx4_ASAP7_75t_L g4302 ( 
.A(n_4095),
.Y(n_4302)
);

INVx1_ASAP7_75t_SL g4303 ( 
.A(n_4025),
.Y(n_4303)
);

OR2x6_ASAP7_75t_L g4304 ( 
.A(n_4043),
.B(n_2567),
.Y(n_4304)
);

AOI21xp5_ASAP7_75t_L g4305 ( 
.A1(n_4112),
.A2(n_2540),
.B(n_2528),
.Y(n_4305)
);

A2O1A1Ixp33_ASAP7_75t_L g4306 ( 
.A1(n_4051),
.A2(n_4082),
.B(n_4050),
.C(n_4114),
.Y(n_4306)
);

OA21x2_ASAP7_75t_L g4307 ( 
.A1(n_4016),
.A2(n_1530),
.B(n_1502),
.Y(n_4307)
);

NOR2xp67_ASAP7_75t_L g4308 ( 
.A(n_4059),
.B(n_6),
.Y(n_4308)
);

AO21x2_ASAP7_75t_L g4309 ( 
.A1(n_4073),
.A2(n_2569),
.B(n_2568),
.Y(n_4309)
);

OAI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_4081),
.A2(n_1027),
.B(n_1023),
.Y(n_4310)
);

AOI21xp5_ASAP7_75t_L g4311 ( 
.A1(n_3958),
.A2(n_2540),
.B(n_2551),
.Y(n_4311)
);

NAND3x1_ASAP7_75t_L g4312 ( 
.A(n_3991),
.B(n_2597),
.C(n_2551),
.Y(n_4312)
);

AO21x1_ASAP7_75t_L g4313 ( 
.A1(n_3996),
.A2(n_9),
.B(n_10),
.Y(n_4313)
);

OR2x2_ASAP7_75t_L g4314 ( 
.A(n_4021),
.B(n_4034),
.Y(n_4314)
);

OAI21x1_ASAP7_75t_L g4315 ( 
.A1(n_4143),
.A2(n_2569),
.B(n_2568),
.Y(n_4315)
);

AO31x2_ASAP7_75t_L g4316 ( 
.A1(n_4115),
.A2(n_2573),
.A3(n_2579),
.B(n_2574),
.Y(n_4316)
);

OAI21x1_ASAP7_75t_L g4317 ( 
.A1(n_4091),
.A2(n_2574),
.B(n_2573),
.Y(n_4317)
);

AOI21xp5_ASAP7_75t_L g4318 ( 
.A1(n_4030),
.A2(n_2551),
.B(n_2597),
.Y(n_4318)
);

INVx4_ASAP7_75t_SL g4319 ( 
.A(n_4044),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4031),
.Y(n_4320)
);

INVx4_ASAP7_75t_SL g4321 ( 
.A(n_4044),
.Y(n_4321)
);

HB1xp67_ASAP7_75t_L g4322 ( 
.A(n_4106),
.Y(n_4322)
);

AOI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_4030),
.A2(n_2597),
.B(n_2582),
.Y(n_4323)
);

AO31x2_ASAP7_75t_L g4324 ( 
.A1(n_4096),
.A2(n_2579),
.A3(n_2583),
.B(n_2582),
.Y(n_4324)
);

AOI22xp5_ASAP7_75t_L g4325 ( 
.A1(n_4110),
.A2(n_1029),
.B1(n_1034),
.B2(n_1032),
.Y(n_4325)
);

OAI221xp5_ASAP7_75t_L g4326 ( 
.A1(n_4134),
.A2(n_1037),
.B1(n_1038),
.B2(n_1036),
.C(n_1035),
.Y(n_4326)
);

OAI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_4105),
.A2(n_1041),
.B(n_1039),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4064),
.Y(n_4328)
);

AO21x2_ASAP7_75t_L g4329 ( 
.A1(n_4075),
.A2(n_2587),
.B(n_2583),
.Y(n_4329)
);

OR2x2_ASAP7_75t_L g4330 ( 
.A(n_4034),
.B(n_1100),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_4004),
.B(n_1100),
.Y(n_4331)
);

A2O1A1Ixp33_ASAP7_75t_L g4332 ( 
.A1(n_4102),
.A2(n_1050),
.B(n_1051),
.C(n_1049),
.Y(n_4332)
);

OA21x2_ASAP7_75t_L g4333 ( 
.A1(n_4072),
.A2(n_2593),
.B(n_2587),
.Y(n_4333)
);

AOI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_4109),
.A2(n_4061),
.B(n_4059),
.Y(n_4334)
);

BUFx3_ASAP7_75t_L g4335 ( 
.A(n_3928),
.Y(n_4335)
);

AOI22xp33_ASAP7_75t_L g4336 ( 
.A1(n_3997),
.A2(n_2594),
.B1(n_2626),
.B2(n_2593),
.Y(n_4336)
);

BUFx12f_ASAP7_75t_L g4337 ( 
.A(n_4095),
.Y(n_4337)
);

CKINVDCx11_ASAP7_75t_R g4338 ( 
.A(n_3917),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_4059),
.A2(n_2626),
.B(n_2594),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_4126),
.B(n_9),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_4124),
.B(n_10),
.Y(n_4341)
);

AOI21xp5_ASAP7_75t_L g4342 ( 
.A1(n_4061),
.A2(n_2640),
.B(n_2636),
.Y(n_4342)
);

OAI21x1_ASAP7_75t_L g4343 ( 
.A1(n_4017),
.A2(n_2640),
.B(n_2636),
.Y(n_4343)
);

AOI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_4061),
.A2(n_2416),
.B(n_2334),
.Y(n_4344)
);

HB1xp67_ASAP7_75t_L g4345 ( 
.A(n_4108),
.Y(n_4345)
);

A2O1A1Ixp33_ASAP7_75t_L g4346 ( 
.A1(n_3913),
.A2(n_1059),
.B(n_1062),
.C(n_1058),
.Y(n_4346)
);

OAI21x1_ASAP7_75t_L g4347 ( 
.A1(n_4020),
.A2(n_2334),
.B(n_2316),
.Y(n_4347)
);

AND2x4_ASAP7_75t_L g4348 ( 
.A(n_4039),
.B(n_11),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_4039),
.B(n_11),
.Y(n_4349)
);

OR2x2_ASAP7_75t_L g4350 ( 
.A(n_3963),
.B(n_12),
.Y(n_4350)
);

AND2x4_ASAP7_75t_L g4351 ( 
.A(n_4092),
.B(n_13),
.Y(n_4351)
);

OAI21xp5_ASAP7_75t_L g4352 ( 
.A1(n_3977),
.A2(n_1065),
.B(n_1064),
.Y(n_4352)
);

OR2x2_ASAP7_75t_L g4353 ( 
.A(n_3963),
.B(n_14),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4092),
.B(n_14),
.Y(n_4354)
);

AO21x2_ASAP7_75t_L g4355 ( 
.A1(n_3913),
.A2(n_2327),
.B(n_2416),
.Y(n_4355)
);

NOR2xp33_ASAP7_75t_SL g4356 ( 
.A(n_3978),
.B(n_727),
.Y(n_4356)
);

OAI21x1_ASAP7_75t_L g4357 ( 
.A1(n_4032),
.A2(n_2334),
.B(n_2316),
.Y(n_4357)
);

O2A1O1Ixp33_ASAP7_75t_L g4358 ( 
.A1(n_4038),
.A2(n_1192),
.B(n_1244),
.C(n_1177),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4142),
.Y(n_4359)
);

OAI21x1_ASAP7_75t_L g4360 ( 
.A1(n_4141),
.A2(n_2316),
.B(n_1916),
.Y(n_4360)
);

AO32x2_ASAP7_75t_L g4361 ( 
.A1(n_3978),
.A2(n_3999),
.A3(n_4018),
.B1(n_3982),
.B2(n_3964),
.Y(n_4361)
);

OAI21x1_ASAP7_75t_L g4362 ( 
.A1(n_3964),
.A2(n_1916),
.B(n_1192),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_3982),
.B(n_3999),
.Y(n_4363)
);

NOR2xp33_ASAP7_75t_L g4364 ( 
.A(n_4018),
.B(n_15),
.Y(n_4364)
);

AOI22xp33_ASAP7_75t_L g4365 ( 
.A1(n_4127),
.A2(n_727),
.B1(n_1916),
.B2(n_1068),
.Y(n_4365)
);

OAI21x1_ASAP7_75t_L g4366 ( 
.A1(n_3964),
.A2(n_1244),
.B(n_1177),
.Y(n_4366)
);

NOR2xp67_ASAP7_75t_L g4367 ( 
.A(n_3928),
.B(n_15),
.Y(n_4367)
);

AOI22xp5_ASAP7_75t_L g4368 ( 
.A1(n_3936),
.A2(n_4127),
.B1(n_4142),
.B2(n_3940),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_3940),
.B(n_16),
.Y(n_4369)
);

INVx2_ASAP7_75t_L g4370 ( 
.A(n_4108),
.Y(n_4370)
);

AOI22xp5_ASAP7_75t_L g4371 ( 
.A1(n_3936),
.A2(n_1066),
.B1(n_1075),
.B2(n_1073),
.Y(n_4371)
);

AOI21xp5_ASAP7_75t_L g4372 ( 
.A1(n_4127),
.A2(n_4108),
.B(n_4067),
.Y(n_4372)
);

BUFx10_ASAP7_75t_L g4373 ( 
.A(n_3917),
.Y(n_4373)
);

O2A1O1Ixp5_ASAP7_75t_L g4374 ( 
.A1(n_3964),
.A2(n_1263),
.B(n_1280),
.C(n_1247),
.Y(n_4374)
);

AO31x2_ASAP7_75t_L g4375 ( 
.A1(n_3917),
.A2(n_1247),
.A3(n_1280),
.B(n_1263),
.Y(n_4375)
);

AOI21xp5_ASAP7_75t_L g4376 ( 
.A1(n_4067),
.A2(n_1077),
.B(n_1076),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_3936),
.A2(n_727),
.B1(n_1079),
.B2(n_1078),
.Y(n_4377)
);

AOI21xp5_ASAP7_75t_L g4378 ( 
.A1(n_4067),
.A2(n_1085),
.B(n_1082),
.Y(n_4378)
);

AOI21xp5_ASAP7_75t_L g4379 ( 
.A1(n_4063),
.A2(n_4033),
.B(n_3998),
.Y(n_4379)
);

OAI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_4063),
.A2(n_1089),
.B1(n_1090),
.B2(n_1087),
.Y(n_4380)
);

AOI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_4063),
.A2(n_1093),
.B(n_1092),
.Y(n_4381)
);

AOI22xp33_ASAP7_75t_L g4382 ( 
.A1(n_4151),
.A2(n_3962),
.B1(n_3969),
.B2(n_3952),
.Y(n_4382)
);

A2O1A1Ixp33_ASAP7_75t_SL g4383 ( 
.A1(n_4364),
.A2(n_1303),
.B(n_1310),
.C(n_1292),
.Y(n_4383)
);

OAI22xp33_ASAP7_75t_L g4384 ( 
.A1(n_4176),
.A2(n_3972),
.B1(n_3952),
.B2(n_3969),
.Y(n_4384)
);

AOI21x1_ASAP7_75t_L g4385 ( 
.A1(n_4331),
.A2(n_1303),
.B(n_1292),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4287),
.Y(n_4386)
);

CKINVDCx20_ASAP7_75t_R g4387 ( 
.A(n_4187),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_4162),
.B(n_4044),
.Y(n_4388)
);

OAI21x1_ASAP7_75t_L g4389 ( 
.A1(n_4172),
.A2(n_4044),
.B(n_3962),
.Y(n_4389)
);

OAI21x1_ASAP7_75t_L g4390 ( 
.A1(n_4227),
.A2(n_3962),
.B(n_3952),
.Y(n_4390)
);

BUFx6f_ASAP7_75t_L g4391 ( 
.A(n_4337),
.Y(n_4391)
);

HB1xp67_ASAP7_75t_L g4392 ( 
.A(n_4258),
.Y(n_4392)
);

OR2x2_ASAP7_75t_L g4393 ( 
.A(n_4290),
.B(n_3969),
.Y(n_4393)
);

AOI22xp5_ASAP7_75t_SL g4394 ( 
.A1(n_4211),
.A2(n_3936),
.B1(n_4012),
.B2(n_3972),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4144),
.Y(n_4395)
);

OAI222xp33_ASAP7_75t_L g4396 ( 
.A1(n_4293),
.A2(n_1098),
.B1(n_1096),
.B2(n_1101),
.C1(n_1097),
.C2(n_1095),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4174),
.Y(n_4397)
);

OAI21x1_ASAP7_75t_L g4398 ( 
.A1(n_4152),
.A2(n_4012),
.B(n_3972),
.Y(n_4398)
);

A2O1A1Ixp33_ASAP7_75t_L g4399 ( 
.A1(n_4332),
.A2(n_1130),
.B(n_1116),
.C(n_1103),
.Y(n_4399)
);

INVx3_ASAP7_75t_L g4400 ( 
.A(n_4285),
.Y(n_4400)
);

OA21x2_ASAP7_75t_L g4401 ( 
.A1(n_4372),
.A2(n_1105),
.B(n_1102),
.Y(n_4401)
);

OAI21xp5_ASAP7_75t_L g4402 ( 
.A1(n_4236),
.A2(n_1117),
.B(n_1112),
.Y(n_4402)
);

BUFx2_ASAP7_75t_L g4403 ( 
.A(n_4361),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_4210),
.B(n_4012),
.Y(n_4404)
);

OA21x2_ASAP7_75t_L g4405 ( 
.A1(n_4157),
.A2(n_1123),
.B(n_1121),
.Y(n_4405)
);

OAI21x1_ASAP7_75t_L g4406 ( 
.A1(n_4312),
.A2(n_1330),
.B(n_1310),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_4280),
.B(n_16),
.Y(n_4407)
);

AND2x2_ASAP7_75t_L g4408 ( 
.A(n_4217),
.B(n_17),
.Y(n_4408)
);

OAI21x1_ASAP7_75t_L g4409 ( 
.A1(n_4250),
.A2(n_4175),
.B(n_4164),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4322),
.Y(n_4410)
);

INVx4_ASAP7_75t_SL g4411 ( 
.A(n_4160),
.Y(n_4411)
);

NAND2xp33_ASAP7_75t_L g4412 ( 
.A(n_4160),
.B(n_4303),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4229),
.Y(n_4413)
);

OAI21x1_ASAP7_75t_L g4414 ( 
.A1(n_4216),
.A2(n_1351),
.B(n_1330),
.Y(n_4414)
);

INVx1_ASAP7_75t_SL g4415 ( 
.A(n_4167),
.Y(n_4415)
);

INVx2_ASAP7_75t_L g4416 ( 
.A(n_4286),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_4286),
.Y(n_4417)
);

OAI21x1_ASAP7_75t_L g4418 ( 
.A1(n_4214),
.A2(n_1364),
.B(n_1351),
.Y(n_4418)
);

AND2x4_ASAP7_75t_L g4419 ( 
.A(n_4319),
.B(n_18),
.Y(n_4419)
);

OA21x2_ASAP7_75t_L g4420 ( 
.A1(n_4145),
.A2(n_1127),
.B(n_1124),
.Y(n_4420)
);

CKINVDCx5p33_ASAP7_75t_R g4421 ( 
.A(n_4147),
.Y(n_4421)
);

AOI221xp5_ASAP7_75t_L g4422 ( 
.A1(n_4161),
.A2(n_1129),
.B1(n_1128),
.B2(n_1372),
.C(n_1364),
.Y(n_4422)
);

OR2x6_ASAP7_75t_L g4423 ( 
.A(n_4334),
.B(n_1298),
.Y(n_4423)
);

INVx2_ASAP7_75t_L g4424 ( 
.A(n_4173),
.Y(n_4424)
);

AOI21xp33_ASAP7_75t_L g4425 ( 
.A1(n_4313),
.A2(n_19),
.B(n_20),
.Y(n_4425)
);

NOR2xp33_ASAP7_75t_SL g4426 ( 
.A(n_4306),
.B(n_4285),
.Y(n_4426)
);

A2O1A1Ixp33_ASAP7_75t_L g4427 ( 
.A1(n_4283),
.A2(n_23),
.B(n_20),
.C(n_22),
.Y(n_4427)
);

AND2x4_ASAP7_75t_L g4428 ( 
.A(n_4319),
.B(n_22),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_4154),
.B(n_23),
.Y(n_4429)
);

OAI21x1_ASAP7_75t_L g4430 ( 
.A1(n_4263),
.A2(n_1399),
.B(n_1372),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4220),
.Y(n_4431)
);

OAI21x1_ASAP7_75t_L g4432 ( 
.A1(n_4195),
.A2(n_1399),
.B(n_727),
.Y(n_4432)
);

AND2x4_ASAP7_75t_L g4433 ( 
.A(n_4321),
.B(n_4282),
.Y(n_4433)
);

NAND2xp33_ASAP7_75t_L g4434 ( 
.A(n_4160),
.B(n_727),
.Y(n_4434)
);

OAI21x1_ASAP7_75t_L g4435 ( 
.A1(n_4155),
.A2(n_4225),
.B(n_4347),
.Y(n_4435)
);

AOI22xp33_ASAP7_75t_L g4436 ( 
.A1(n_4201),
.A2(n_727),
.B1(n_1304),
.B2(n_1298),
.Y(n_4436)
);

OAI22xp5_ASAP7_75t_L g4437 ( 
.A1(n_4296),
.A2(n_28),
.B1(n_25),
.B2(n_26),
.Y(n_4437)
);

AO31x2_ASAP7_75t_L g4438 ( 
.A1(n_4251),
.A2(n_4190),
.A3(n_4219),
.B(n_4169),
.Y(n_4438)
);

OAI21x1_ASAP7_75t_SL g4439 ( 
.A1(n_4182),
.A2(n_25),
.B(n_26),
.Y(n_4439)
);

OAI21x1_ASAP7_75t_L g4440 ( 
.A1(n_4232),
.A2(n_28),
.B(n_29),
.Y(n_4440)
);

BUFx3_ASAP7_75t_L g4441 ( 
.A(n_4189),
.Y(n_4441)
);

CKINVDCx8_ASAP7_75t_R g4442 ( 
.A(n_4177),
.Y(n_4442)
);

AND2x2_ASAP7_75t_L g4443 ( 
.A(n_4171),
.B(n_30),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_4180),
.Y(n_4444)
);

INVx2_ASAP7_75t_SL g4445 ( 
.A(n_4208),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4284),
.Y(n_4446)
);

NAND2xp33_ASAP7_75t_SL g4447 ( 
.A(n_4196),
.B(n_30),
.Y(n_4447)
);

AND2x4_ASAP7_75t_L g4448 ( 
.A(n_4321),
.B(n_32),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_4320),
.Y(n_4449)
);

BUFx12f_ASAP7_75t_L g4450 ( 
.A(n_4241),
.Y(n_4450)
);

OAI21x1_ASAP7_75t_L g4451 ( 
.A1(n_4299),
.A2(n_32),
.B(n_34),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4159),
.B(n_35),
.Y(n_4452)
);

OAI21xp5_ASAP7_75t_L g4453 ( 
.A1(n_4183),
.A2(n_37),
.B(n_39),
.Y(n_4453)
);

OA21x2_ASAP7_75t_L g4454 ( 
.A1(n_4264),
.A2(n_37),
.B(n_40),
.Y(n_4454)
);

BUFx6f_ASAP7_75t_L g4455 ( 
.A(n_4259),
.Y(n_4455)
);

OAI21x1_ASAP7_75t_L g4456 ( 
.A1(n_4343),
.A2(n_41),
.B(n_42),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_4328),
.B(n_4262),
.Y(n_4457)
);

CKINVDCx5p33_ASAP7_75t_R g4458 ( 
.A(n_4239),
.Y(n_4458)
);

INVx3_ASAP7_75t_L g4459 ( 
.A(n_4302),
.Y(n_4459)
);

OAI22xp5_ASAP7_75t_L g4460 ( 
.A1(n_4156),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_4460)
);

OAI21x1_ASAP7_75t_L g4461 ( 
.A1(n_4315),
.A2(n_4360),
.B(n_4230),
.Y(n_4461)
);

NOR2xp33_ASAP7_75t_L g4462 ( 
.A(n_4224),
.B(n_43),
.Y(n_4462)
);

AO21x2_ASAP7_75t_L g4463 ( 
.A1(n_4256),
.A2(n_46),
.B(n_47),
.Y(n_4463)
);

OAI22xp5_ASAP7_75t_L g4464 ( 
.A1(n_4212),
.A2(n_4291),
.B1(n_4246),
.B2(n_4340),
.Y(n_4464)
);

O2A1O1Ixp33_ASAP7_75t_SL g4465 ( 
.A1(n_4254),
.A2(n_51),
.B(n_48),
.C(n_49),
.Y(n_4465)
);

AND2x2_ASAP7_75t_L g4466 ( 
.A(n_4363),
.B(n_48),
.Y(n_4466)
);

OR2x2_ASAP7_75t_L g4467 ( 
.A(n_4235),
.B(n_53),
.Y(n_4467)
);

INVx1_ASAP7_75t_SL g4468 ( 
.A(n_4206),
.Y(n_4468)
);

OAI21x1_ASAP7_75t_L g4469 ( 
.A1(n_4244),
.A2(n_54),
.B(n_55),
.Y(n_4469)
);

BUFx2_ASAP7_75t_L g4470 ( 
.A(n_4361),
.Y(n_4470)
);

OAI21x1_ASAP7_75t_L g4471 ( 
.A1(n_4270),
.A2(n_55),
.B(n_56),
.Y(n_4471)
);

INVx6_ASAP7_75t_L g4472 ( 
.A(n_4373),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4186),
.Y(n_4473)
);

BUFx12f_ASAP7_75t_L g4474 ( 
.A(n_4338),
.Y(n_4474)
);

INVx5_ASAP7_75t_L g4475 ( 
.A(n_4259),
.Y(n_4475)
);

OAI21x1_ASAP7_75t_L g4476 ( 
.A1(n_4275),
.A2(n_56),
.B(n_58),
.Y(n_4476)
);

OAI21x1_ASAP7_75t_L g4477 ( 
.A1(n_4297),
.A2(n_59),
.B(n_60),
.Y(n_4477)
);

OAI21x1_ASAP7_75t_L g4478 ( 
.A1(n_4298),
.A2(n_59),
.B(n_61),
.Y(n_4478)
);

AO21x2_ASAP7_75t_L g4479 ( 
.A1(n_4184),
.A2(n_61),
.B(n_62),
.Y(n_4479)
);

OAI21xp5_ASAP7_75t_L g4480 ( 
.A1(n_4185),
.A2(n_62),
.B(n_63),
.Y(n_4480)
);

OAI21x1_ASAP7_75t_L g4481 ( 
.A1(n_4271),
.A2(n_63),
.B(n_64),
.Y(n_4481)
);

INVx1_ASAP7_75t_SL g4482 ( 
.A(n_4192),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4146),
.B(n_64),
.Y(n_4483)
);

AND2x2_ASAP7_75t_L g4484 ( 
.A(n_4361),
.B(n_65),
.Y(n_4484)
);

CKINVDCx11_ASAP7_75t_R g4485 ( 
.A(n_4177),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4193),
.Y(n_4486)
);

OA21x2_ASAP7_75t_L g4487 ( 
.A1(n_4199),
.A2(n_66),
.B(n_69),
.Y(n_4487)
);

OAI21x1_ASAP7_75t_L g4488 ( 
.A1(n_4170),
.A2(n_70),
.B(n_71),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_4223),
.B(n_71),
.Y(n_4489)
);

BUFx2_ASAP7_75t_L g4490 ( 
.A(n_4302),
.Y(n_4490)
);

AOI21xp5_ASAP7_75t_L g4491 ( 
.A1(n_4267),
.A2(n_1304),
.B(n_1298),
.Y(n_4491)
);

INVx2_ASAP7_75t_L g4492 ( 
.A(n_4200),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4146),
.B(n_72),
.Y(n_4493)
);

INVx2_ASAP7_75t_L g4494 ( 
.A(n_4228),
.Y(n_4494)
);

OAI21x1_ASAP7_75t_L g4495 ( 
.A1(n_4242),
.A2(n_73),
.B(n_74),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_4247),
.Y(n_4496)
);

OAI21x1_ASAP7_75t_L g4497 ( 
.A1(n_4272),
.A2(n_73),
.B(n_74),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_4215),
.B(n_75),
.Y(n_4498)
);

OAI21x1_ASAP7_75t_SL g4499 ( 
.A1(n_4349),
.A2(n_75),
.B(n_76),
.Y(n_4499)
);

BUFx3_ASAP7_75t_L g4500 ( 
.A(n_4335),
.Y(n_4500)
);

AND2x4_ASAP7_75t_L g4501 ( 
.A(n_4359),
.B(n_76),
.Y(n_4501)
);

OAI21x1_ASAP7_75t_SL g4502 ( 
.A1(n_4354),
.A2(n_4341),
.B(n_4158),
.Y(n_4502)
);

AO31x2_ASAP7_75t_L g4503 ( 
.A1(n_4370),
.A2(n_80),
.A3(n_77),
.B(n_78),
.Y(n_4503)
);

OAI21x1_ASAP7_75t_L g4504 ( 
.A1(n_4179),
.A2(n_78),
.B(n_80),
.Y(n_4504)
);

OAI21xp33_ASAP7_75t_SL g4505 ( 
.A1(n_4238),
.A2(n_82),
.B(n_84),
.Y(n_4505)
);

AOI21xp5_ASAP7_75t_L g4506 ( 
.A1(n_4276),
.A2(n_1304),
.B(n_1298),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4252),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4255),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4281),
.Y(n_4509)
);

AOI222xp33_ASAP7_75t_L g4510 ( 
.A1(n_4178),
.A2(n_88),
.B1(n_90),
.B2(n_85),
.C1(n_87),
.C2(n_89),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4288),
.Y(n_4511)
);

NOR2xp33_ASAP7_75t_L g4512 ( 
.A(n_4369),
.B(n_85),
.Y(n_4512)
);

AOI21xp5_ASAP7_75t_L g4513 ( 
.A1(n_4374),
.A2(n_1304),
.B(n_1298),
.Y(n_4513)
);

AND2x2_ASAP7_75t_L g4514 ( 
.A(n_4314),
.B(n_90),
.Y(n_4514)
);

CKINVDCx5p33_ASAP7_75t_R g4515 ( 
.A(n_4345),
.Y(n_4515)
);

OAI21x1_ASAP7_75t_L g4516 ( 
.A1(n_4257),
.A2(n_91),
.B(n_92),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_4274),
.Y(n_4517)
);

INVx4_ASAP7_75t_L g4518 ( 
.A(n_4348),
.Y(n_4518)
);

NOR2xp33_ASAP7_75t_L g4519 ( 
.A(n_4348),
.B(n_91),
.Y(n_4519)
);

INVx2_ASAP7_75t_L g4520 ( 
.A(n_4209),
.Y(n_4520)
);

NAND2xp33_ASAP7_75t_R g4521 ( 
.A(n_4351),
.B(n_92),
.Y(n_4521)
);

OAI21xp5_ASAP7_75t_L g4522 ( 
.A1(n_4148),
.A2(n_93),
.B(n_94),
.Y(n_4522)
);

AO21x2_ASAP7_75t_L g4523 ( 
.A1(n_4309),
.A2(n_93),
.B(n_94),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4221),
.Y(n_4524)
);

OAI21x1_ASAP7_75t_L g4525 ( 
.A1(n_4307),
.A2(n_95),
.B(n_96),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4221),
.Y(n_4526)
);

INVx5_ASAP7_75t_L g4527 ( 
.A(n_4304),
.Y(n_4527)
);

OAI21x1_ASAP7_75t_L g4528 ( 
.A1(n_4307),
.A2(n_95),
.B(n_98),
.Y(n_4528)
);

INVx6_ASAP7_75t_L g4529 ( 
.A(n_4373),
.Y(n_4529)
);

OAI22xp5_ASAP7_75t_L g4530 ( 
.A1(n_4371),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_4530)
);

OR2x2_ASAP7_75t_L g4531 ( 
.A(n_4294),
.B(n_101),
.Y(n_4531)
);

OR2x2_ASAP7_75t_L g4532 ( 
.A(n_4218),
.B(n_101),
.Y(n_4532)
);

HB1xp67_ASAP7_75t_L g4533 ( 
.A(n_4279),
.Y(n_4533)
);

AO21x2_ASAP7_75t_L g4534 ( 
.A1(n_4329),
.A2(n_102),
.B(n_103),
.Y(n_4534)
);

INVx2_ASAP7_75t_SL g4535 ( 
.A(n_4351),
.Y(n_4535)
);

O2A1O1Ixp33_ASAP7_75t_SL g4536 ( 
.A1(n_4197),
.A2(n_105),
.B(n_102),
.C(n_103),
.Y(n_4536)
);

OAI21x1_ASAP7_75t_L g4537 ( 
.A1(n_4191),
.A2(n_4357),
.B(n_4362),
.Y(n_4537)
);

INVx1_ASAP7_75t_SL g4538 ( 
.A(n_4330),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4209),
.Y(n_4539)
);

OAI21x1_ASAP7_75t_L g4540 ( 
.A1(n_4240),
.A2(n_105),
.B(n_107),
.Y(n_4540)
);

O2A1O1Ixp33_ASAP7_75t_SL g4541 ( 
.A1(n_4346),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_4541)
);

A2O1A1Ixp33_ASAP7_75t_L g4542 ( 
.A1(n_4367),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_4542)
);

OAI21x1_ASAP7_75t_L g4543 ( 
.A1(n_4202),
.A2(n_111),
.B(n_113),
.Y(n_4543)
);

OAI22xp5_ASAP7_75t_L g4544 ( 
.A1(n_4163),
.A2(n_116),
.B1(n_111),
.B2(n_115),
.Y(n_4544)
);

AND2x4_ASAP7_75t_L g4545 ( 
.A(n_4379),
.B(n_116),
.Y(n_4545)
);

OR2x6_ASAP7_75t_L g4546 ( 
.A(n_4304),
.B(n_1304),
.Y(n_4546)
);

BUFx2_ASAP7_75t_L g4547 ( 
.A(n_4350),
.Y(n_4547)
);

OAI22xp5_ASAP7_75t_L g4548 ( 
.A1(n_4377),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_4548)
);

INVxp67_ASAP7_75t_SL g4549 ( 
.A(n_4333),
.Y(n_4549)
);

CKINVDCx5p33_ASAP7_75t_R g4550 ( 
.A(n_4368),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4221),
.Y(n_4551)
);

OAI22xp5_ASAP7_75t_L g4552 ( 
.A1(n_4353),
.A2(n_121),
.B1(n_117),
.B2(n_120),
.Y(n_4552)
);

OAI21x1_ASAP7_75t_L g4553 ( 
.A1(n_4278),
.A2(n_121),
.B(n_122),
.Y(n_4553)
);

OAI21x1_ASAP7_75t_L g4554 ( 
.A1(n_4317),
.A2(n_122),
.B(n_123),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_4166),
.B(n_4153),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4222),
.Y(n_4556)
);

INVx2_ASAP7_75t_SL g4557 ( 
.A(n_4355),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4222),
.Y(n_4558)
);

OAI21x1_ASAP7_75t_L g4559 ( 
.A1(n_4333),
.A2(n_123),
.B(n_124),
.Y(n_4559)
);

AOI22xp33_ASAP7_75t_SL g4560 ( 
.A1(n_4356),
.A2(n_1393),
.B1(n_1420),
.B2(n_1367),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_4222),
.Y(n_4561)
);

AOI22xp33_ASAP7_75t_L g4562 ( 
.A1(n_4336),
.A2(n_1393),
.B1(n_1420),
.B2(n_1367),
.Y(n_4562)
);

AOI21xp5_ASAP7_75t_L g4563 ( 
.A1(n_4292),
.A2(n_1393),
.B(n_1367),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4153),
.Y(n_4564)
);

OAI21x1_ASAP7_75t_SL g4565 ( 
.A1(n_4310),
.A2(n_4327),
.B(n_4245),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4153),
.Y(n_4566)
);

AOI21xp5_ASAP7_75t_L g4567 ( 
.A1(n_4305),
.A2(n_1393),
.B(n_1367),
.Y(n_4567)
);

INVx3_ASAP7_75t_L g4568 ( 
.A(n_4324),
.Y(n_4568)
);

CKINVDCx20_ASAP7_75t_R g4569 ( 
.A(n_4380),
.Y(n_4569)
);

AOI22xp33_ASAP7_75t_L g4570 ( 
.A1(n_4464),
.A2(n_4268),
.B1(n_4149),
.B2(n_4295),
.Y(n_4570)
);

BUFx3_ASAP7_75t_L g4571 ( 
.A(n_4387),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4386),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4395),
.Y(n_4573)
);

OA21x2_ASAP7_75t_L g4574 ( 
.A1(n_4403),
.A2(n_4308),
.B(n_4366),
.Y(n_4574)
);

NOR2xp33_ASAP7_75t_L g4575 ( 
.A(n_4442),
.B(n_4273),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4449),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4392),
.Y(n_4577)
);

AOI22xp5_ASAP7_75t_L g4578 ( 
.A1(n_4464),
.A2(n_4181),
.B1(n_4165),
.B2(n_4352),
.Y(n_4578)
);

CKINVDCx12_ASAP7_75t_R g4579 ( 
.A(n_4394),
.Y(n_4579)
);

AND2x2_ASAP7_75t_L g4580 ( 
.A(n_4415),
.B(n_4203),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4415),
.B(n_4203),
.Y(n_4581)
);

OAI22xp33_ASAP7_75t_L g4582 ( 
.A1(n_4531),
.A2(n_4301),
.B1(n_4311),
.B2(n_4325),
.Y(n_4582)
);

BUFx2_ASAP7_75t_L g4583 ( 
.A(n_4474),
.Y(n_4583)
);

BUFx3_ASAP7_75t_L g4584 ( 
.A(n_4450),
.Y(n_4584)
);

BUFx3_ASAP7_75t_L g4585 ( 
.A(n_4441),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4457),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4410),
.B(n_4457),
.Y(n_4587)
);

INVx6_ASAP7_75t_L g4588 ( 
.A(n_4411),
.Y(n_4588)
);

INVx2_ASAP7_75t_SL g4589 ( 
.A(n_4515),
.Y(n_4589)
);

AND2x2_ASAP7_75t_L g4590 ( 
.A(n_4547),
.B(n_4203),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4444),
.Y(n_4591)
);

INVx2_ASAP7_75t_L g4592 ( 
.A(n_4473),
.Y(n_4592)
);

BUFx6f_ASAP7_75t_L g4593 ( 
.A(n_4546),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4500),
.B(n_4168),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4397),
.Y(n_4595)
);

BUFx10_ASAP7_75t_L g4596 ( 
.A(n_4462),
.Y(n_4596)
);

AND2x4_ASAP7_75t_L g4597 ( 
.A(n_4433),
.B(n_4324),
.Y(n_4597)
);

NAND2xp33_ASAP7_75t_R g4598 ( 
.A(n_4458),
.B(n_4269),
.Y(n_4598)
);

AND2x2_ASAP7_75t_L g4599 ( 
.A(n_4388),
.B(n_4168),
.Y(n_4599)
);

CKINVDCx5p33_ASAP7_75t_R g4600 ( 
.A(n_4421),
.Y(n_4600)
);

NOR2xp33_ASAP7_75t_L g4601 ( 
.A(n_4485),
.B(n_4326),
.Y(n_4601)
);

AOI22xp33_ASAP7_75t_L g4602 ( 
.A1(n_4425),
.A2(n_4249),
.B1(n_4365),
.B2(n_4231),
.Y(n_4602)
);

AOI22xp33_ASAP7_75t_L g4603 ( 
.A1(n_4425),
.A2(n_4289),
.B1(n_4381),
.B2(n_4378),
.Y(n_4603)
);

OR2x2_ASAP7_75t_L g4604 ( 
.A(n_4538),
.B(n_4168),
.Y(n_4604)
);

INVxp67_ASAP7_75t_L g4605 ( 
.A(n_4502),
.Y(n_4605)
);

OAI22xp33_ASAP7_75t_L g4606 ( 
.A1(n_4521),
.A2(n_4194),
.B1(n_4205),
.B2(n_4260),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4413),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4446),
.Y(n_4608)
);

AOI22xp33_ASAP7_75t_L g4609 ( 
.A1(n_4401),
.A2(n_4376),
.B1(n_4339),
.B2(n_4342),
.Y(n_4609)
);

OAI22xp5_ASAP7_75t_L g4610 ( 
.A1(n_4427),
.A2(n_4460),
.B1(n_4437),
.B2(n_4484),
.Y(n_4610)
);

NAND3xp33_ASAP7_75t_L g4611 ( 
.A(n_4505),
.B(n_4207),
.C(n_4150),
.Y(n_4611)
);

AOI222xp33_ASAP7_75t_L g4612 ( 
.A1(n_4505),
.A2(n_4460),
.B1(n_4530),
.B2(n_4522),
.C1(n_4437),
.C2(n_4565),
.Y(n_4612)
);

AND2x4_ASAP7_75t_L g4613 ( 
.A(n_4433),
.B(n_4324),
.Y(n_4613)
);

NAND3xp33_ASAP7_75t_L g4614 ( 
.A(n_4510),
.B(n_4204),
.C(n_4266),
.Y(n_4614)
);

INVx1_ASAP7_75t_SL g4615 ( 
.A(n_4490),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_SL g4616 ( 
.A(n_4394),
.B(n_4237),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4538),
.B(n_4316),
.Y(n_4617)
);

OR2x2_ASAP7_75t_L g4618 ( 
.A(n_4404),
.B(n_4316),
.Y(n_4618)
);

AOI21xp33_ASAP7_75t_L g4619 ( 
.A1(n_4405),
.A2(n_4261),
.B(n_4300),
.Y(n_4619)
);

OAI22xp5_ASAP7_75t_L g4620 ( 
.A1(n_4518),
.A2(n_4198),
.B1(n_4213),
.B2(n_4243),
.Y(n_4620)
);

OR2x2_ASAP7_75t_L g4621 ( 
.A(n_4404),
.B(n_4316),
.Y(n_4621)
);

AND2x2_ASAP7_75t_L g4622 ( 
.A(n_4470),
.B(n_4375),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4535),
.B(n_4375),
.Y(n_4623)
);

OR2x2_ASAP7_75t_L g4624 ( 
.A(n_4393),
.B(n_4533),
.Y(n_4624)
);

AND2x2_ASAP7_75t_L g4625 ( 
.A(n_4445),
.B(n_4375),
.Y(n_4625)
);

AOI22xp33_ASAP7_75t_L g4626 ( 
.A1(n_4401),
.A2(n_4417),
.B1(n_4416),
.B2(n_4405),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4483),
.B(n_4226),
.Y(n_4627)
);

OAI22xp33_ASAP7_75t_L g4628 ( 
.A1(n_4426),
.A2(n_4483),
.B1(n_4493),
.B2(n_4402),
.Y(n_4628)
);

AOI222xp33_ASAP7_75t_L g4629 ( 
.A1(n_4522),
.A2(n_4530),
.B1(n_4402),
.B2(n_4447),
.C1(n_4480),
.C2(n_4453),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4518),
.B(n_4226),
.Y(n_4630)
);

NOR2xp33_ASAP7_75t_L g4631 ( 
.A(n_4391),
.B(n_124),
.Y(n_4631)
);

AND2x4_ASAP7_75t_L g4632 ( 
.A(n_4411),
.B(n_4226),
.Y(n_4632)
);

AOI22xp33_ASAP7_75t_L g4633 ( 
.A1(n_4520),
.A2(n_4277),
.B1(n_4323),
.B2(n_4234),
.Y(n_4633)
);

OR2x2_ASAP7_75t_L g4634 ( 
.A(n_4511),
.B(n_4248),
.Y(n_4634)
);

AOI22xp33_ASAP7_75t_SL g4635 ( 
.A1(n_4426),
.A2(n_4233),
.B1(n_4344),
.B2(n_4318),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4486),
.Y(n_4636)
);

OR2x2_ASAP7_75t_L g4637 ( 
.A(n_4482),
.B(n_4248),
.Y(n_4637)
);

OAI22xp33_ASAP7_75t_L g4638 ( 
.A1(n_4493),
.A2(n_4265),
.B1(n_4253),
.B2(n_4358),
.Y(n_4638)
);

AOI22xp33_ASAP7_75t_L g4639 ( 
.A1(n_4539),
.A2(n_1393),
.B1(n_1420),
.B2(n_1367),
.Y(n_4639)
);

AND2x4_ASAP7_75t_L g4640 ( 
.A(n_4400),
.B(n_4248),
.Y(n_4640)
);

CKINVDCx20_ASAP7_75t_R g4641 ( 
.A(n_4569),
.Y(n_4641)
);

AOI22xp33_ASAP7_75t_SL g4642 ( 
.A1(n_4420),
.A2(n_1543),
.B1(n_1420),
.B2(n_127),
.Y(n_4642)
);

AND2x4_ASAP7_75t_L g4643 ( 
.A(n_4400),
.B(n_125),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4459),
.B(n_125),
.Y(n_4644)
);

A2O1A1Ixp33_ASAP7_75t_L g4645 ( 
.A1(n_4512),
.A2(n_4188),
.B(n_128),
.C(n_126),
.Y(n_4645)
);

AOI22xp33_ASAP7_75t_L g4646 ( 
.A1(n_4510),
.A2(n_1543),
.B1(n_1420),
.B2(n_130),
.Y(n_4646)
);

OR2x2_ASAP7_75t_L g4647 ( 
.A(n_4482),
.B(n_127),
.Y(n_4647)
);

AOI22xp33_ASAP7_75t_L g4648 ( 
.A1(n_4454),
.A2(n_1543),
.B1(n_132),
.B2(n_128),
.Y(n_4648)
);

OAI22xp5_ASAP7_75t_L g4649 ( 
.A1(n_4552),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4429),
.B(n_133),
.Y(n_4650)
);

NOR2xp33_ASAP7_75t_L g4651 ( 
.A(n_4391),
.B(n_134),
.Y(n_4651)
);

OR2x6_ASAP7_75t_L g4652 ( 
.A(n_4389),
.B(n_1543),
.Y(n_4652)
);

AOI22xp33_ASAP7_75t_L g4653 ( 
.A1(n_4454),
.A2(n_1543),
.B1(n_137),
.B2(n_135),
.Y(n_4653)
);

AOI22xp33_ASAP7_75t_L g4654 ( 
.A1(n_4487),
.A2(n_4420),
.B1(n_4480),
.B2(n_4453),
.Y(n_4654)
);

NOR2xp33_ASAP7_75t_L g4655 ( 
.A(n_4391),
.B(n_4412),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4459),
.B(n_136),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4496),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4507),
.Y(n_4658)
);

OAI22xp5_ASAP7_75t_L g4659 ( 
.A1(n_4552),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_4659)
);

NOR2xp33_ASAP7_75t_L g4660 ( 
.A(n_4396),
.B(n_138),
.Y(n_4660)
);

OAI221xp5_ASAP7_75t_L g4661 ( 
.A1(n_4542),
.A2(n_4399),
.B1(n_4382),
.B2(n_4536),
.C(n_4548),
.Y(n_4661)
);

CKINVDCx5p33_ASAP7_75t_R g4662 ( 
.A(n_4550),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4508),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4492),
.Y(n_4664)
);

AOI22xp33_ASAP7_75t_SL g4665 ( 
.A1(n_4487),
.A2(n_143),
.B1(n_140),
.B2(n_142),
.Y(n_4665)
);

HB1xp67_ASAP7_75t_L g4666 ( 
.A(n_4514),
.Y(n_4666)
);

NOR3xp33_ASAP7_75t_SL g4667 ( 
.A(n_4519),
.B(n_142),
.C(n_144),
.Y(n_4667)
);

BUFx3_ASAP7_75t_L g4668 ( 
.A(n_4501),
.Y(n_4668)
);

AOI22xp33_ASAP7_75t_L g4669 ( 
.A1(n_4479),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4509),
.Y(n_4670)
);

OR2x2_ASAP7_75t_L g4671 ( 
.A(n_4468),
.B(n_4494),
.Y(n_4671)
);

INVx4_ASAP7_75t_SL g4672 ( 
.A(n_4419),
.Y(n_4672)
);

OAI22xp5_ASAP7_75t_L g4673 ( 
.A1(n_4419),
.A2(n_153),
.B1(n_148),
.B2(n_151),
.Y(n_4673)
);

BUFx2_ASAP7_75t_L g4674 ( 
.A(n_4472),
.Y(n_4674)
);

OAI22xp5_ASAP7_75t_L g4675 ( 
.A1(n_4428),
.A2(n_156),
.B1(n_151),
.B2(n_155),
.Y(n_4675)
);

NOR2xp33_ASAP7_75t_R g4676 ( 
.A(n_4428),
.B(n_155),
.Y(n_4676)
);

OAI22xp5_ASAP7_75t_L g4677 ( 
.A1(n_4448),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_4677)
);

AO21x2_ASAP7_75t_L g4678 ( 
.A1(n_4555),
.A2(n_157),
.B(n_159),
.Y(n_4678)
);

A2O1A1Ixp33_ASAP7_75t_L g4679 ( 
.A1(n_4448),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_4679)
);

OAI221xp5_ASAP7_75t_L g4680 ( 
.A1(n_4548),
.A2(n_166),
.B1(n_160),
.B2(n_165),
.C(n_167),
.Y(n_4680)
);

INVx2_ASAP7_75t_L g4681 ( 
.A(n_4424),
.Y(n_4681)
);

BUFx4f_ASAP7_75t_L g4682 ( 
.A(n_4501),
.Y(n_4682)
);

OAI22xp5_ASAP7_75t_L g4683 ( 
.A1(n_4498),
.A2(n_168),
.B1(n_165),
.B2(n_167),
.Y(n_4683)
);

BUFx2_ASAP7_75t_L g4684 ( 
.A(n_4472),
.Y(n_4684)
);

AND2x2_ASAP7_75t_L g4685 ( 
.A(n_4466),
.B(n_168),
.Y(n_4685)
);

CKINVDCx11_ASAP7_75t_R g4686 ( 
.A(n_4545),
.Y(n_4686)
);

AO31x2_ASAP7_75t_L g4687 ( 
.A1(n_4564),
.A2(n_171),
.A3(n_169),
.B(n_170),
.Y(n_4687)
);

CKINVDCx5p33_ASAP7_75t_R g4688 ( 
.A(n_4529),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4517),
.Y(n_4689)
);

AND2x4_ASAP7_75t_L g4690 ( 
.A(n_4390),
.B(n_4468),
.Y(n_4690)
);

AOI22xp33_ASAP7_75t_L g4691 ( 
.A1(n_4479),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_4691)
);

NAND2xp33_ASAP7_75t_SL g4692 ( 
.A(n_4407),
.B(n_173),
.Y(n_4692)
);

INVx2_ASAP7_75t_L g4693 ( 
.A(n_4431),
.Y(n_4693)
);

BUFx6f_ASAP7_75t_L g4694 ( 
.A(n_4546),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4557),
.Y(n_4695)
);

OAI22xp33_ASAP7_75t_L g4696 ( 
.A1(n_4475),
.A2(n_177),
.B1(n_174),
.B2(n_175),
.Y(n_4696)
);

BUFx3_ASAP7_75t_L g4697 ( 
.A(n_4443),
.Y(n_4697)
);

CKINVDCx5p33_ASAP7_75t_R g4698 ( 
.A(n_4529),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4566),
.Y(n_4699)
);

INVx8_ASAP7_75t_L g4700 ( 
.A(n_4546),
.Y(n_4700)
);

NAND2xp33_ASAP7_75t_R g4701 ( 
.A(n_4545),
.B(n_175),
.Y(n_4701)
);

CKINVDCx5p33_ASAP7_75t_R g4702 ( 
.A(n_4408),
.Y(n_4702)
);

OAI21xp5_ASAP7_75t_L g4703 ( 
.A1(n_4488),
.A2(n_179),
.B(n_180),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4524),
.Y(n_4704)
);

OR2x2_ASAP7_75t_L g4705 ( 
.A(n_4467),
.B(n_181),
.Y(n_4705)
);

BUFx2_ASAP7_75t_L g4706 ( 
.A(n_4435),
.Y(n_4706)
);

NAND2x1_ASAP7_75t_L g4707 ( 
.A(n_4423),
.B(n_181),
.Y(n_4707)
);

AOI221xp5_ASAP7_75t_L g4708 ( 
.A1(n_4541),
.A2(n_186),
.B1(n_183),
.B2(n_185),
.C(n_187),
.Y(n_4708)
);

NAND2xp33_ASAP7_75t_R g4709 ( 
.A(n_4452),
.B(n_183),
.Y(n_4709)
);

AND2x2_ASAP7_75t_L g4710 ( 
.A(n_4455),
.B(n_185),
.Y(n_4710)
);

NAND2x1p5_ASAP7_75t_L g4711 ( 
.A(n_4475),
.B(n_187),
.Y(n_4711)
);

BUFx8_ASAP7_75t_SL g4712 ( 
.A(n_4489),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4398),
.Y(n_4713)
);

AOI22xp5_ASAP7_75t_L g4714 ( 
.A1(n_4544),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_4714)
);

CKINVDCx6p67_ASAP7_75t_R g4715 ( 
.A(n_4498),
.Y(n_4715)
);

INVx2_ASAP7_75t_SL g4716 ( 
.A(n_4532),
.Y(n_4716)
);

BUFx2_ASAP7_75t_L g4717 ( 
.A(n_4503),
.Y(n_4717)
);

AOI22xp33_ASAP7_75t_L g4718 ( 
.A1(n_4614),
.A2(n_4523),
.B1(n_4534),
.B2(n_4463),
.Y(n_4718)
);

AOI22xp33_ASAP7_75t_L g4719 ( 
.A1(n_4614),
.A2(n_4523),
.B1(n_4534),
.B2(n_4463),
.Y(n_4719)
);

AOI22xp33_ASAP7_75t_L g4720 ( 
.A1(n_4612),
.A2(n_4499),
.B1(n_4544),
.B2(n_4384),
.Y(n_4720)
);

AOI21xp5_ASAP7_75t_L g4721 ( 
.A1(n_4628),
.A2(n_4423),
.B(n_4383),
.Y(n_4721)
);

OAI22xp33_ASAP7_75t_L g4722 ( 
.A1(n_4610),
.A2(n_4423),
.B1(n_4527),
.B2(n_4475),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_4576),
.Y(n_4723)
);

A2O1A1Ixp33_ASAP7_75t_L g4724 ( 
.A1(n_4654),
.A2(n_4434),
.B(n_4549),
.C(n_4471),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4573),
.Y(n_4725)
);

AND2x4_ASAP7_75t_L g4726 ( 
.A(n_4672),
.B(n_4716),
.Y(n_4726)
);

OAI211xp5_ASAP7_75t_L g4727 ( 
.A1(n_4629),
.A2(n_4465),
.B(n_4422),
.C(n_4409),
.Y(n_4727)
);

AOI21xp5_ASAP7_75t_L g4728 ( 
.A1(n_4606),
.A2(n_4491),
.B(n_4563),
.Y(n_4728)
);

OAI21x1_ASAP7_75t_L g4729 ( 
.A1(n_4713),
.A2(n_4568),
.B(n_4461),
.Y(n_4729)
);

BUFx2_ASAP7_75t_L g4730 ( 
.A(n_4588),
.Y(n_4730)
);

AND2x4_ASAP7_75t_L g4731 ( 
.A(n_4672),
.B(n_4455),
.Y(n_4731)
);

AOI21xp5_ASAP7_75t_L g4732 ( 
.A1(n_4616),
.A2(n_4567),
.B(n_4439),
.Y(n_4732)
);

OAI221xp5_ASAP7_75t_L g4733 ( 
.A1(n_4626),
.A2(n_4436),
.B1(n_4556),
.B2(n_4551),
.C(n_4526),
.Y(n_4733)
);

OAI22xp33_ASAP7_75t_L g4734 ( 
.A1(n_4701),
.A2(n_4578),
.B1(n_4709),
.B2(n_4582),
.Y(n_4734)
);

OAI21xp5_ASAP7_75t_L g4735 ( 
.A1(n_4605),
.A2(n_4476),
.B(n_4469),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4634),
.Y(n_4736)
);

AND2x2_ASAP7_75t_L g4737 ( 
.A(n_4666),
.B(n_4674),
.Y(n_4737)
);

AOI222xp33_ASAP7_75t_L g4738 ( 
.A1(n_4611),
.A2(n_4478),
.B1(n_4477),
.B2(n_4559),
.C1(n_4504),
.C2(n_4553),
.Y(n_4738)
);

AOI22xp33_ASAP7_75t_L g4739 ( 
.A1(n_4629),
.A2(n_4558),
.B1(n_4561),
.B2(n_4455),
.Y(n_4739)
);

AOI21xp5_ASAP7_75t_L g4740 ( 
.A1(n_4707),
.A2(n_4527),
.B(n_4506),
.Y(n_4740)
);

AOI22xp33_ASAP7_75t_L g4741 ( 
.A1(n_4611),
.A2(n_4527),
.B1(n_4528),
.B2(n_4525),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_4684),
.B(n_4543),
.Y(n_4742)
);

OR2x2_ASAP7_75t_L g4743 ( 
.A(n_4587),
.B(n_4503),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4615),
.B(n_4697),
.Y(n_4744)
);

OA21x2_ASAP7_75t_L g4745 ( 
.A1(n_4695),
.A2(n_4706),
.B(n_4699),
.Y(n_4745)
);

AOI22xp33_ASAP7_75t_L g4746 ( 
.A1(n_4678),
.A2(n_4568),
.B1(n_4516),
.B2(n_4451),
.Y(n_4746)
);

BUFx2_ASAP7_75t_L g4747 ( 
.A(n_4588),
.Y(n_4747)
);

AOI221xp5_ASAP7_75t_L g4748 ( 
.A1(n_4660),
.A2(n_4503),
.B1(n_4513),
.B2(n_4562),
.C(n_191),
.Y(n_4748)
);

AOI221xp5_ASAP7_75t_L g4749 ( 
.A1(n_4683),
.A2(n_192),
.B1(n_188),
.B2(n_190),
.C(n_193),
.Y(n_4749)
);

OAI222xp33_ASAP7_75t_L g4750 ( 
.A1(n_4717),
.A2(n_4385),
.B1(n_4560),
.B2(n_4438),
.C1(n_4537),
.C2(n_4456),
.Y(n_4750)
);

OAI21xp5_ASAP7_75t_L g4751 ( 
.A1(n_4665),
.A2(n_4440),
.B(n_4554),
.Y(n_4751)
);

A2O1A1Ixp33_ASAP7_75t_L g4752 ( 
.A1(n_4575),
.A2(n_4481),
.B(n_4540),
.C(n_4497),
.Y(n_4752)
);

OAI221xp5_ASAP7_75t_L g4753 ( 
.A1(n_4578),
.A2(n_4438),
.B1(n_4495),
.B2(n_4406),
.C(n_197),
.Y(n_4753)
);

AOI22xp33_ASAP7_75t_L g4754 ( 
.A1(n_4678),
.A2(n_4432),
.B1(n_4418),
.B2(n_4430),
.Y(n_4754)
);

AND2x6_ASAP7_75t_SL g4755 ( 
.A(n_4601),
.B(n_194),
.Y(n_4755)
);

AOI22xp33_ASAP7_75t_L g4756 ( 
.A1(n_4646),
.A2(n_4414),
.B1(n_4438),
.B2(n_198),
.Y(n_4756)
);

INVx2_ASAP7_75t_L g4757 ( 
.A(n_4618),
.Y(n_4757)
);

NAND2x1p5_ASAP7_75t_L g4758 ( 
.A(n_4682),
.B(n_194),
.Y(n_4758)
);

AO21x2_ASAP7_75t_L g4759 ( 
.A1(n_4627),
.A2(n_196),
.B(n_198),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4586),
.B(n_200),
.Y(n_4760)
);

NAND2x1_ASAP7_75t_L g4761 ( 
.A(n_4577),
.B(n_4690),
.Y(n_4761)
);

OAI21x1_ASAP7_75t_L g4762 ( 
.A1(n_4617),
.A2(n_201),
.B(n_202),
.Y(n_4762)
);

NAND2xp33_ASAP7_75t_R g4763 ( 
.A(n_4676),
.B(n_202),
.Y(n_4763)
);

NAND4xp25_ASAP7_75t_L g4764 ( 
.A(n_4708),
.B(n_205),
.C(n_203),
.D(n_204),
.Y(n_4764)
);

AOI21xp5_ASAP7_75t_L g4765 ( 
.A1(n_4635),
.A2(n_204),
.B(n_206),
.Y(n_4765)
);

AOI22xp33_ASAP7_75t_L g4766 ( 
.A1(n_4661),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4595),
.Y(n_4767)
);

OAI22x1_ASAP7_75t_L g4768 ( 
.A1(n_4702),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_4768)
);

AOI21xp5_ASAP7_75t_L g4769 ( 
.A1(n_4638),
.A2(n_210),
.B(n_213),
.Y(n_4769)
);

INVx2_ASAP7_75t_SL g4770 ( 
.A(n_4583),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_L g4771 ( 
.A(n_4615),
.B(n_216),
.Y(n_4771)
);

NOR2xp67_ASAP7_75t_L g4772 ( 
.A(n_4580),
.B(n_216),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4607),
.B(n_218),
.Y(n_4773)
);

AOI22xp33_ASAP7_75t_L g4774 ( 
.A1(n_4599),
.A2(n_222),
.B1(n_219),
.B2(n_221),
.Y(n_4774)
);

OAI22xp5_ASAP7_75t_SL g4775 ( 
.A1(n_4579),
.A2(n_222),
.B1(n_219),
.B2(n_221),
.Y(n_4775)
);

OAI322xp33_ASAP7_75t_L g4776 ( 
.A1(n_4714),
.A2(n_223),
.A3(n_224),
.B1(n_225),
.B2(n_226),
.C1(n_227),
.C2(n_228),
.Y(n_4776)
);

AOI22xp33_ASAP7_75t_L g4777 ( 
.A1(n_4570),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4608),
.Y(n_4778)
);

AO21x2_ASAP7_75t_L g4779 ( 
.A1(n_4704),
.A2(n_4650),
.B(n_4581),
.Y(n_4779)
);

AOI22xp33_ASAP7_75t_L g4780 ( 
.A1(n_4619),
.A2(n_230),
.B1(n_227),
.B2(n_229),
.Y(n_4780)
);

AOI22xp5_ASAP7_75t_L g4781 ( 
.A1(n_4714),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_4781)
);

BUFx3_ASAP7_75t_L g4782 ( 
.A(n_4571),
.Y(n_4782)
);

INVx3_ASAP7_75t_L g4783 ( 
.A(n_4640),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4636),
.B(n_231),
.Y(n_4784)
);

OA21x2_ASAP7_75t_L g4785 ( 
.A1(n_4690),
.A2(n_4590),
.B(n_4622),
.Y(n_4785)
);

BUFx2_ASAP7_75t_L g4786 ( 
.A(n_4688),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4715),
.B(n_232),
.Y(n_4787)
);

OAI22xp5_ASAP7_75t_L g4788 ( 
.A1(n_4682),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_4788)
);

INVx3_ASAP7_75t_L g4789 ( 
.A(n_4640),
.Y(n_4789)
);

INVx3_ASAP7_75t_L g4790 ( 
.A(n_4584),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4657),
.B(n_233),
.Y(n_4791)
);

INVx2_ASAP7_75t_L g4792 ( 
.A(n_4621),
.Y(n_4792)
);

AOI22xp33_ASAP7_75t_L g4793 ( 
.A1(n_4596),
.A2(n_239),
.B1(n_236),
.B2(n_238),
.Y(n_4793)
);

OAI221xp5_ASAP7_75t_L g4794 ( 
.A1(n_4642),
.A2(n_4669),
.B1(n_4691),
.B2(n_4653),
.C(n_4648),
.Y(n_4794)
);

BUFx6f_ASAP7_75t_L g4795 ( 
.A(n_4593),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4658),
.B(n_238),
.Y(n_4796)
);

OAI22xp5_ASAP7_75t_L g4797 ( 
.A1(n_4668),
.A2(n_4667),
.B1(n_4679),
.B2(n_4633),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_L g4798 ( 
.A(n_4663),
.B(n_4670),
.Y(n_4798)
);

AOI21xp33_ASAP7_75t_L g4799 ( 
.A1(n_4652),
.A2(n_239),
.B(n_240),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4689),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4572),
.Y(n_4801)
);

AOI22xp33_ASAP7_75t_L g4802 ( 
.A1(n_4596),
.A2(n_246),
.B1(n_241),
.B2(n_243),
.Y(n_4802)
);

OA21x2_ASAP7_75t_L g4803 ( 
.A1(n_4604),
.A2(n_243),
.B(n_246),
.Y(n_4803)
);

AO21x2_ASAP7_75t_L g4804 ( 
.A1(n_4594),
.A2(n_249),
.B(n_252),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_SL g4805 ( 
.A(n_4698),
.B(n_249),
.Y(n_4805)
);

OAI211xp5_ASAP7_75t_L g4806 ( 
.A1(n_4680),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_4806)
);

AOI21xp5_ASAP7_75t_L g4807 ( 
.A1(n_4645),
.A2(n_253),
.B(n_254),
.Y(n_4807)
);

INVx2_ASAP7_75t_L g4808 ( 
.A(n_4623),
.Y(n_4808)
);

INVx3_ASAP7_75t_L g4809 ( 
.A(n_4643),
.Y(n_4809)
);

AND2x2_ASAP7_75t_L g4810 ( 
.A(n_4589),
.B(n_255),
.Y(n_4810)
);

AO31x2_ASAP7_75t_L g4811 ( 
.A1(n_4655),
.A2(n_4659),
.A3(n_4649),
.B(n_4591),
.Y(n_4811)
);

AOI222xp33_ASAP7_75t_L g4812 ( 
.A1(n_4692),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.C1(n_259),
.C2(n_260),
.Y(n_4812)
);

OR2x2_ASAP7_75t_L g4813 ( 
.A(n_4624),
.B(n_257),
.Y(n_4813)
);

AOI22xp33_ASAP7_75t_L g4814 ( 
.A1(n_4602),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_4814)
);

AOI22xp33_ASAP7_75t_L g4815 ( 
.A1(n_4609),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_4815)
);

OAI22xp5_ASAP7_75t_L g4816 ( 
.A1(n_4643),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4637),
.Y(n_4817)
);

OAI211xp5_ASAP7_75t_L g4818 ( 
.A1(n_4703),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_4818)
);

OA21x2_ASAP7_75t_L g4819 ( 
.A1(n_4597),
.A2(n_266),
.B(n_267),
.Y(n_4819)
);

OAI22xp33_ASAP7_75t_L g4820 ( 
.A1(n_4647),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4671),
.Y(n_4821)
);

A2O1A1Ixp33_ASAP7_75t_L g4822 ( 
.A1(n_4631),
.A2(n_271),
.B(n_269),
.C(n_270),
.Y(n_4822)
);

AOI22xp33_ASAP7_75t_L g4823 ( 
.A1(n_4630),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_4823)
);

AOI221xp5_ASAP7_75t_L g4824 ( 
.A1(n_4673),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.C(n_278),
.Y(n_4824)
);

AOI21xp5_ASAP7_75t_L g4825 ( 
.A1(n_4696),
.A2(n_276),
.B(n_278),
.Y(n_4825)
);

OAI211xp5_ASAP7_75t_SL g4826 ( 
.A1(n_4603),
.A2(n_282),
.B(n_279),
.C(n_281),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4625),
.B(n_279),
.Y(n_4827)
);

A2O1A1Ixp33_ASAP7_75t_L g4828 ( 
.A1(n_4651),
.A2(n_283),
.B(n_281),
.C(n_282),
.Y(n_4828)
);

NAND2xp5_ASAP7_75t_L g4829 ( 
.A(n_4644),
.B(n_4656),
.Y(n_4829)
);

AOI22xp33_ASAP7_75t_L g4830 ( 
.A1(n_4641),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_4830)
);

OAI221xp5_ASAP7_75t_SL g4831 ( 
.A1(n_4705),
.A2(n_288),
.B1(n_284),
.B2(n_286),
.C(n_289),
.Y(n_4831)
);

AND2x4_ASAP7_75t_L g4832 ( 
.A(n_4597),
.B(n_288),
.Y(n_4832)
);

NOR2x1_ASAP7_75t_SL g4833 ( 
.A(n_4652),
.B(n_290),
.Y(n_4833)
);

AOI21xp5_ASAP7_75t_L g4834 ( 
.A1(n_4700),
.A2(n_291),
.B(n_292),
.Y(n_4834)
);

AOI22xp33_ASAP7_75t_L g4835 ( 
.A1(n_4574),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_4835)
);

OAI22xp5_ASAP7_75t_L g4836 ( 
.A1(n_4711),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_4836)
);

AOI21xp5_ASAP7_75t_L g4837 ( 
.A1(n_4700),
.A2(n_294),
.B(n_296),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_L g4838 ( 
.A(n_4687),
.B(n_296),
.Y(n_4838)
);

OR2x2_ASAP7_75t_L g4839 ( 
.A(n_4592),
.B(n_298),
.Y(n_4839)
);

AOI22xp33_ASAP7_75t_L g4840 ( 
.A1(n_4574),
.A2(n_302),
.B1(n_298),
.B2(n_300),
.Y(n_4840)
);

OAI21x1_ASAP7_75t_L g4841 ( 
.A1(n_4664),
.A2(n_302),
.B(n_304),
.Y(n_4841)
);

AO21x2_ASAP7_75t_L g4842 ( 
.A1(n_4632),
.A2(n_305),
.B(n_306),
.Y(n_4842)
);

AOI221xp5_ASAP7_75t_L g4843 ( 
.A1(n_4675),
.A2(n_308),
.B1(n_305),
.B2(n_307),
.C(n_309),
.Y(n_4843)
);

OAI21x1_ASAP7_75t_L g4844 ( 
.A1(n_4681),
.A2(n_307),
.B(n_308),
.Y(n_4844)
);

OAI22xp5_ASAP7_75t_L g4845 ( 
.A1(n_4677),
.A2(n_315),
.B1(n_311),
.B2(n_312),
.Y(n_4845)
);

NAND2xp5_ASAP7_75t_L g4846 ( 
.A(n_4687),
.B(n_312),
.Y(n_4846)
);

NAND2x1p5_ASAP7_75t_L g4847 ( 
.A(n_4585),
.B(n_315),
.Y(n_4847)
);

AOI211xp5_ASAP7_75t_SL g4848 ( 
.A1(n_4620),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_L g4849 ( 
.A(n_4687),
.B(n_316),
.Y(n_4849)
);

BUFx3_ASAP7_75t_L g4850 ( 
.A(n_4600),
.Y(n_4850)
);

AND2x4_ASAP7_75t_L g4851 ( 
.A(n_4613),
.B(n_318),
.Y(n_4851)
);

AOI22xp33_ASAP7_75t_L g4852 ( 
.A1(n_4693),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4613),
.Y(n_4853)
);

AOI22xp33_ASAP7_75t_SL g4854 ( 
.A1(n_4700),
.A2(n_325),
.B1(n_322),
.B2(n_323),
.Y(n_4854)
);

AOI221xp5_ASAP7_75t_L g4855 ( 
.A1(n_4685),
.A2(n_328),
.B1(n_323),
.B2(n_327),
.C(n_329),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4593),
.Y(n_4856)
);

NOR2xp33_ASAP7_75t_R g4857 ( 
.A(n_4790),
.B(n_4598),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4798),
.Y(n_4858)
);

AND2x4_ASAP7_75t_L g4859 ( 
.A(n_4726),
.B(n_4730),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4759),
.B(n_4710),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4759),
.B(n_4686),
.Y(n_4861)
);

XNOR2xp5_ASAP7_75t_L g4862 ( 
.A(n_4734),
.B(n_4662),
.Y(n_4862)
);

NAND2xp33_ASAP7_75t_SL g4863 ( 
.A(n_4744),
.B(n_4593),
.Y(n_4863)
);

NAND2xp33_ASAP7_75t_R g4864 ( 
.A(n_4819),
.B(n_4652),
.Y(n_4864)
);

NOR2xp33_ASAP7_75t_R g4865 ( 
.A(n_4790),
.B(n_4712),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4725),
.Y(n_4866)
);

AND2x4_ASAP7_75t_L g4867 ( 
.A(n_4726),
.B(n_4747),
.Y(n_4867)
);

AND2x2_ASAP7_75t_L g4868 ( 
.A(n_4737),
.B(n_4632),
.Y(n_4868)
);

NAND2xp33_ASAP7_75t_R g4869 ( 
.A(n_4819),
.B(n_327),
.Y(n_4869)
);

INVx2_ASAP7_75t_L g4870 ( 
.A(n_4842),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_SL g4871 ( 
.A(n_4731),
.B(n_4694),
.Y(n_4871)
);

NAND2xp33_ASAP7_75t_R g4872 ( 
.A(n_4803),
.B(n_328),
.Y(n_4872)
);

NAND2xp33_ASAP7_75t_SL g4873 ( 
.A(n_4809),
.B(n_4694),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_SL g4874 ( 
.A(n_4731),
.B(n_4694),
.Y(n_4874)
);

INVxp67_ASAP7_75t_L g4875 ( 
.A(n_4763),
.Y(n_4875)
);

INVxp67_ASAP7_75t_L g4876 ( 
.A(n_4770),
.Y(n_4876)
);

NAND2xp33_ASAP7_75t_R g4877 ( 
.A(n_4803),
.B(n_330),
.Y(n_4877)
);

INVxp33_ASAP7_75t_L g4878 ( 
.A(n_4786),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4718),
.B(n_4639),
.Y(n_4879)
);

NOR2xp33_ASAP7_75t_R g4880 ( 
.A(n_4850),
.B(n_331),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4809),
.B(n_331),
.Y(n_4881)
);

AND2x4_ASAP7_75t_L g4882 ( 
.A(n_4832),
.B(n_4851),
.Y(n_4882)
);

HB1xp67_ASAP7_75t_L g4883 ( 
.A(n_4800),
.Y(n_4883)
);

INVx2_ASAP7_75t_SL g4884 ( 
.A(n_4782),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_L g4885 ( 
.A(n_4719),
.B(n_4767),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4778),
.Y(n_4886)
);

AND2x4_ASAP7_75t_L g4887 ( 
.A(n_4832),
.B(n_332),
.Y(n_4887)
);

OR2x6_ASAP7_75t_L g4888 ( 
.A(n_4758),
.B(n_332),
.Y(n_4888)
);

INVxp67_ASAP7_75t_L g4889 ( 
.A(n_4742),
.Y(n_4889)
);

BUFx12f_ASAP7_75t_L g4890 ( 
.A(n_4755),
.Y(n_4890)
);

OR2x2_ASAP7_75t_L g4891 ( 
.A(n_4821),
.B(n_333),
.Y(n_4891)
);

CKINVDCx5p33_ASAP7_75t_R g4892 ( 
.A(n_4755),
.Y(n_4892)
);

BUFx3_ASAP7_75t_L g4893 ( 
.A(n_4787),
.Y(n_4893)
);

INVxp67_ASAP7_75t_L g4894 ( 
.A(n_4833),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_L g4895 ( 
.A(n_4762),
.B(n_333),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_L g4896 ( 
.A(n_4724),
.B(n_334),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_L g4897 ( 
.A(n_4827),
.B(n_335),
.Y(n_4897)
);

NAND2x1p5_ASAP7_75t_L g4898 ( 
.A(n_4851),
.B(n_335),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4760),
.B(n_336),
.Y(n_4899)
);

NAND2xp33_ASAP7_75t_R g4900 ( 
.A(n_4785),
.B(n_337),
.Y(n_4900)
);

BUFx3_ASAP7_75t_L g4901 ( 
.A(n_4810),
.Y(n_4901)
);

OR2x2_ASAP7_75t_L g4902 ( 
.A(n_4813),
.B(n_337),
.Y(n_4902)
);

AND2x4_ASAP7_75t_L g4903 ( 
.A(n_4735),
.B(n_338),
.Y(n_4903)
);

INVxp67_ASAP7_75t_L g4904 ( 
.A(n_4804),
.Y(n_4904)
);

OR2x6_ASAP7_75t_L g4905 ( 
.A(n_4834),
.B(n_338),
.Y(n_4905)
);

AND2x2_ASAP7_75t_L g4906 ( 
.A(n_4829),
.B(n_340),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_L g4907 ( 
.A(n_4804),
.B(n_340),
.Y(n_4907)
);

INVxp67_ASAP7_75t_L g4908 ( 
.A(n_4797),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4723),
.B(n_341),
.Y(n_4909)
);

NAND2xp33_ASAP7_75t_R g4910 ( 
.A(n_4785),
.B(n_342),
.Y(n_4910)
);

BUFx10_ASAP7_75t_L g4911 ( 
.A(n_4847),
.Y(n_4911)
);

AND2x4_ASAP7_75t_L g4912 ( 
.A(n_4853),
.B(n_343),
.Y(n_4912)
);

NAND2xp33_ASAP7_75t_SL g4913 ( 
.A(n_4761),
.B(n_343),
.Y(n_4913)
);

AND2x4_ASAP7_75t_L g4914 ( 
.A(n_4783),
.B(n_4789),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4838),
.Y(n_4915)
);

CKINVDCx5p33_ASAP7_75t_R g4916 ( 
.A(n_4795),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4846),
.Y(n_4917)
);

AND2x2_ASAP7_75t_L g4918 ( 
.A(n_4811),
.B(n_344),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_L g4919 ( 
.A(n_4779),
.B(n_345),
.Y(n_4919)
);

NOR2xp33_ASAP7_75t_R g4920 ( 
.A(n_4771),
.B(n_345),
.Y(n_4920)
);

INVxp67_ASAP7_75t_L g4921 ( 
.A(n_4856),
.Y(n_4921)
);

INVxp67_ASAP7_75t_L g4922 ( 
.A(n_4842),
.Y(n_4922)
);

NOR2xp33_ASAP7_75t_L g4923 ( 
.A(n_4805),
.B(n_346),
.Y(n_4923)
);

NAND2xp33_ASAP7_75t_R g4924 ( 
.A(n_4765),
.B(n_346),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4849),
.Y(n_4925)
);

AND2x4_ASAP7_75t_L g4926 ( 
.A(n_4811),
.B(n_351),
.Y(n_4926)
);

INVxp67_ASAP7_75t_SL g4927 ( 
.A(n_4745),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_4773),
.Y(n_4928)
);

NOR2xp33_ASAP7_75t_L g4929 ( 
.A(n_4784),
.B(n_351),
.Y(n_4929)
);

INVxp67_ASAP7_75t_L g4930 ( 
.A(n_4779),
.Y(n_4930)
);

AND2x4_ASAP7_75t_L g4931 ( 
.A(n_4783),
.B(n_4789),
.Y(n_4931)
);

INVxp67_ASAP7_75t_L g4932 ( 
.A(n_4839),
.Y(n_4932)
);

OR2x6_ASAP7_75t_L g4933 ( 
.A(n_4837),
.B(n_352),
.Y(n_4933)
);

AND2x2_ASAP7_75t_L g4934 ( 
.A(n_4811),
.B(n_352),
.Y(n_4934)
);

INVxp67_ASAP7_75t_L g4935 ( 
.A(n_4791),
.Y(n_4935)
);

AND2x4_ASAP7_75t_L g4936 ( 
.A(n_4752),
.B(n_354),
.Y(n_4936)
);

AND2x2_ASAP7_75t_L g4937 ( 
.A(n_4796),
.B(n_355),
.Y(n_4937)
);

NOR2xp33_ASAP7_75t_R g4938 ( 
.A(n_4766),
.B(n_356),
.Y(n_4938)
);

INVx2_ASAP7_75t_L g4939 ( 
.A(n_4795),
.Y(n_4939)
);

INVxp67_ASAP7_75t_L g4940 ( 
.A(n_4768),
.Y(n_4940)
);

CKINVDCx5p33_ASAP7_75t_R g4941 ( 
.A(n_4795),
.Y(n_4941)
);

NAND2xp33_ASAP7_75t_R g4942 ( 
.A(n_4745),
.B(n_356),
.Y(n_4942)
);

NAND2xp33_ASAP7_75t_R g4943 ( 
.A(n_4769),
.B(n_357),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4743),
.B(n_4720),
.Y(n_4944)
);

NOR2xp33_ASAP7_75t_L g4945 ( 
.A(n_4831),
.B(n_357),
.Y(n_4945)
);

BUFx10_ASAP7_75t_L g4946 ( 
.A(n_4775),
.Y(n_4946)
);

BUFx3_ASAP7_75t_L g4947 ( 
.A(n_4775),
.Y(n_4947)
);

AND2x2_ASAP7_75t_L g4948 ( 
.A(n_4739),
.B(n_359),
.Y(n_4948)
);

NOR2xp33_ASAP7_75t_R g4949 ( 
.A(n_4793),
.B(n_359),
.Y(n_4949)
);

BUFx10_ASAP7_75t_L g4950 ( 
.A(n_4788),
.Y(n_4950)
);

NAND2xp33_ASAP7_75t_SL g4951 ( 
.A(n_4816),
.B(n_360),
.Y(n_4951)
);

INVxp33_ASAP7_75t_L g4952 ( 
.A(n_4772),
.Y(n_4952)
);

NOR2xp33_ASAP7_75t_SL g4953 ( 
.A(n_4764),
.B(n_361),
.Y(n_4953)
);

AND2x2_ASAP7_75t_L g4954 ( 
.A(n_4808),
.B(n_361),
.Y(n_4954)
);

INVx2_ASAP7_75t_L g4955 ( 
.A(n_4729),
.Y(n_4955)
);

CKINVDCx8_ASAP7_75t_R g4956 ( 
.A(n_4848),
.Y(n_4956)
);

OR2x2_ASAP7_75t_L g4957 ( 
.A(n_4757),
.B(n_362),
.Y(n_4957)
);

AND2x4_ASAP7_75t_L g4958 ( 
.A(n_4746),
.B(n_362),
.Y(n_4958)
);

NAND2xp33_ASAP7_75t_R g4959 ( 
.A(n_4732),
.B(n_363),
.Y(n_4959)
);

NAND2xp5_ASAP7_75t_SL g4960 ( 
.A(n_4722),
.B(n_363),
.Y(n_4960)
);

INVxp67_ASAP7_75t_L g4961 ( 
.A(n_4772),
.Y(n_4961)
);

BUFx10_ASAP7_75t_L g4962 ( 
.A(n_4854),
.Y(n_4962)
);

INVx3_ASAP7_75t_L g4963 ( 
.A(n_4859),
.Y(n_4963)
);

AND2x2_ASAP7_75t_L g4964 ( 
.A(n_4859),
.B(n_4792),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4883),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4866),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4886),
.Y(n_4967)
);

AOI22xp33_ASAP7_75t_SL g4968 ( 
.A1(n_4936),
.A2(n_4890),
.B1(n_4944),
.B2(n_4926),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4919),
.Y(n_4969)
);

AND2x2_ASAP7_75t_L g4970 ( 
.A(n_4867),
.B(n_4868),
.Y(n_4970)
);

AND2x2_ASAP7_75t_L g4971 ( 
.A(n_4867),
.B(n_4736),
.Y(n_4971)
);

INVx2_ASAP7_75t_L g4972 ( 
.A(n_4946),
.Y(n_4972)
);

AND2x4_ASAP7_75t_L g4973 ( 
.A(n_4914),
.B(n_4721),
.Y(n_4973)
);

AND2x2_ASAP7_75t_L g4974 ( 
.A(n_4914),
.B(n_4741),
.Y(n_4974)
);

INVx2_ASAP7_75t_L g4975 ( 
.A(n_4918),
.Y(n_4975)
);

INVx2_ASAP7_75t_L g4976 ( 
.A(n_4934),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4935),
.B(n_4727),
.Y(n_4977)
);

INVx2_ASAP7_75t_L g4978 ( 
.A(n_4962),
.Y(n_4978)
);

AND2x4_ASAP7_75t_L g4979 ( 
.A(n_4931),
.B(n_4751),
.Y(n_4979)
);

INVx2_ASAP7_75t_L g4980 ( 
.A(n_4947),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4858),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_4936),
.B(n_4820),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_4907),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_4870),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4915),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4917),
.Y(n_4986)
);

AND2x2_ASAP7_75t_L g4987 ( 
.A(n_4931),
.B(n_4817),
.Y(n_4987)
);

BUFx2_ASAP7_75t_L g4988 ( 
.A(n_4865),
.Y(n_4988)
);

INVx2_ASAP7_75t_L g4989 ( 
.A(n_4957),
.Y(n_4989)
);

INVx1_ASAP7_75t_L g4990 ( 
.A(n_4925),
.Y(n_4990)
);

OR2x2_ASAP7_75t_L g4991 ( 
.A(n_4885),
.B(n_4928),
.Y(n_4991)
);

AND2x2_ASAP7_75t_L g4992 ( 
.A(n_4878),
.B(n_4801),
.Y(n_4992)
);

AND2x2_ASAP7_75t_L g4993 ( 
.A(n_4889),
.B(n_4738),
.Y(n_4993)
);

INVx2_ASAP7_75t_L g4994 ( 
.A(n_4901),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4922),
.Y(n_4995)
);

AND2x2_ASAP7_75t_L g4996 ( 
.A(n_4939),
.B(n_4738),
.Y(n_4996)
);

INVx2_ASAP7_75t_L g4997 ( 
.A(n_4896),
.Y(n_4997)
);

INVx2_ASAP7_75t_L g4998 ( 
.A(n_4893),
.Y(n_4998)
);

INVx2_ASAP7_75t_L g4999 ( 
.A(n_4961),
.Y(n_4999)
);

AOI22xp33_ASAP7_75t_SL g5000 ( 
.A1(n_4857),
.A2(n_4753),
.B1(n_4794),
.B2(n_4818),
.Y(n_5000)
);

INVx2_ASAP7_75t_L g5001 ( 
.A(n_4903),
.Y(n_5001)
);

OR2x2_ASAP7_75t_L g5002 ( 
.A(n_4921),
.B(n_4764),
.Y(n_5002)
);

INVx5_ASAP7_75t_L g5003 ( 
.A(n_4905),
.Y(n_5003)
);

INVx2_ASAP7_75t_L g5004 ( 
.A(n_4903),
.Y(n_5004)
);

INVxp67_ASAP7_75t_SL g5005 ( 
.A(n_4942),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4909),
.Y(n_5006)
);

AND2x4_ASAP7_75t_L g5007 ( 
.A(n_4927),
.B(n_4728),
.Y(n_5007)
);

AND2x2_ASAP7_75t_L g5008 ( 
.A(n_4876),
.B(n_4835),
.Y(n_5008)
);

INVx1_ASAP7_75t_SL g5009 ( 
.A(n_4880),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4891),
.Y(n_5010)
);

HB1xp67_ASAP7_75t_L g5011 ( 
.A(n_4940),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_4908),
.B(n_4774),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4904),
.Y(n_5013)
);

NOR2x1_ASAP7_75t_SL g5014 ( 
.A(n_4888),
.B(n_4836),
.Y(n_5014)
);

AND2x4_ASAP7_75t_L g5015 ( 
.A(n_4955),
.B(n_4840),
.Y(n_5015)
);

INVxp67_ASAP7_75t_R g5016 ( 
.A(n_4881),
.Y(n_5016)
);

BUFx6f_ASAP7_75t_L g5017 ( 
.A(n_4892),
.Y(n_5017)
);

OR2x2_ASAP7_75t_L g5018 ( 
.A(n_4930),
.B(n_4902),
.Y(n_5018)
);

AND2x2_ASAP7_75t_L g5019 ( 
.A(n_4894),
.B(n_4823),
.Y(n_5019)
);

INVx2_ASAP7_75t_L g5020 ( 
.A(n_4950),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_4895),
.Y(n_5021)
);

INVx2_ASAP7_75t_L g5022 ( 
.A(n_4875),
.Y(n_5022)
);

AND2x2_ASAP7_75t_L g5023 ( 
.A(n_4884),
.B(n_4802),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4932),
.Y(n_5024)
);

OAI22xp5_ASAP7_75t_L g5025 ( 
.A1(n_4956),
.A2(n_4781),
.B1(n_4828),
.B2(n_4822),
.Y(n_5025)
);

INVx2_ASAP7_75t_L g5026 ( 
.A(n_4860),
.Y(n_5026)
);

AOI22xp33_ASAP7_75t_L g5027 ( 
.A1(n_4879),
.A2(n_4748),
.B1(n_4807),
.B2(n_4826),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4954),
.Y(n_5028)
);

NOR2xp33_ASAP7_75t_L g5029 ( 
.A(n_4862),
.B(n_4806),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4899),
.Y(n_5030)
);

CKINVDCx6p67_ASAP7_75t_R g5031 ( 
.A(n_4888),
.Y(n_5031)
);

INVx2_ASAP7_75t_L g5032 ( 
.A(n_4958),
.Y(n_5032)
);

AND2x2_ASAP7_75t_L g5033 ( 
.A(n_4882),
.B(n_4781),
.Y(n_5033)
);

NOR2xp67_ASAP7_75t_L g5034 ( 
.A(n_4861),
.B(n_4825),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4906),
.Y(n_5035)
);

BUFx3_ASAP7_75t_L g5036 ( 
.A(n_4911),
.Y(n_5036)
);

INVx2_ASAP7_75t_L g5037 ( 
.A(n_4958),
.Y(n_5037)
);

AND2x2_ASAP7_75t_L g5038 ( 
.A(n_4882),
.B(n_4740),
.Y(n_5038)
);

AOI22xp33_ASAP7_75t_SL g5039 ( 
.A1(n_5005),
.A2(n_4953),
.B1(n_4920),
.B2(n_4948),
.Y(n_5039)
);

OAI211xp5_ASAP7_75t_L g5040 ( 
.A1(n_5000),
.A2(n_4951),
.B(n_4945),
.C(n_4913),
.Y(n_5040)
);

AND2x2_ASAP7_75t_L g5041 ( 
.A(n_4963),
.B(n_4916),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_5035),
.B(n_4937),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_5035),
.B(n_5028),
.Y(n_5043)
);

AND2x2_ASAP7_75t_L g5044 ( 
.A(n_4963),
.B(n_4941),
.Y(n_5044)
);

OAI22xp5_ASAP7_75t_L g5045 ( 
.A1(n_5002),
.A2(n_4960),
.B1(n_4952),
.B2(n_4933),
.Y(n_5045)
);

NAND2xp5_ASAP7_75t_L g5046 ( 
.A(n_5028),
.B(n_4929),
.Y(n_5046)
);

AND2x2_ASAP7_75t_L g5047 ( 
.A(n_4963),
.B(n_4912),
.Y(n_5047)
);

NAND2xp5_ASAP7_75t_L g5048 ( 
.A(n_5010),
.B(n_4912),
.Y(n_5048)
);

OR2x2_ASAP7_75t_SL g5049 ( 
.A(n_5020),
.B(n_4897),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_5010),
.B(n_4923),
.Y(n_5050)
);

AND2x2_ASAP7_75t_L g5051 ( 
.A(n_4970),
.B(n_4898),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_5011),
.Y(n_5052)
);

NOR2xp67_ASAP7_75t_L g5053 ( 
.A(n_5003),
.B(n_4871),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_5013),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_4997),
.B(n_4887),
.Y(n_5055)
);

AND2x2_ASAP7_75t_L g5056 ( 
.A(n_4970),
.B(n_4874),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_L g5057 ( 
.A(n_4997),
.B(n_4905),
.Y(n_5057)
);

AND2x2_ASAP7_75t_L g5058 ( 
.A(n_5036),
.B(n_4933),
.Y(n_5058)
);

OAI21xp5_ASAP7_75t_L g5059 ( 
.A1(n_5025),
.A2(n_4863),
.B(n_4812),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_5030),
.B(n_4855),
.Y(n_5060)
);

NAND2xp5_ASAP7_75t_L g5061 ( 
.A(n_5030),
.B(n_4780),
.Y(n_5061)
);

AND2x2_ASAP7_75t_L g5062 ( 
.A(n_4994),
.B(n_4749),
.Y(n_5062)
);

AOI22xp33_ASAP7_75t_L g5063 ( 
.A1(n_4978),
.A2(n_4949),
.B1(n_4938),
.B2(n_4777),
.Y(n_5063)
);

AOI221xp5_ASAP7_75t_L g5064 ( 
.A1(n_4996),
.A2(n_4776),
.B1(n_4814),
.B2(n_4845),
.C(n_4824),
.Y(n_5064)
);

NAND3xp33_ASAP7_75t_L g5065 ( 
.A(n_4977),
.B(n_4959),
.C(n_4924),
.Y(n_5065)
);

AND2x2_ASAP7_75t_L g5066 ( 
.A(n_5036),
.B(n_4830),
.Y(n_5066)
);

OAI221xp5_ASAP7_75t_SL g5067 ( 
.A1(n_4993),
.A2(n_4843),
.B1(n_4756),
.B2(n_4815),
.C(n_4900),
.Y(n_5067)
);

NAND3xp33_ASAP7_75t_L g5068 ( 
.A(n_5027),
.B(n_4910),
.C(n_4943),
.Y(n_5068)
);

OAI21xp5_ASAP7_75t_SL g5069 ( 
.A1(n_4993),
.A2(n_4750),
.B(n_4799),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_5022),
.B(n_4852),
.Y(n_5070)
);

AOI221xp5_ASAP7_75t_L g5071 ( 
.A1(n_4996),
.A2(n_4776),
.B1(n_4877),
.B2(n_4872),
.C(n_4869),
.Y(n_5071)
);

OAI221xp5_ASAP7_75t_L g5072 ( 
.A1(n_4968),
.A2(n_4864),
.B1(n_4873),
.B2(n_4733),
.C(n_4754),
.Y(n_5072)
);

NAND2xp5_ASAP7_75t_L g5073 ( 
.A(n_5022),
.B(n_4841),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_5013),
.Y(n_5074)
);

NAND4xp25_ASAP7_75t_L g5075 ( 
.A(n_4972),
.B(n_4988),
.C(n_5002),
.D(n_4965),
.Y(n_5075)
);

NAND2xp5_ASAP7_75t_L g5076 ( 
.A(n_5033),
.B(n_4844),
.Y(n_5076)
);

NAND4xp25_ASAP7_75t_L g5077 ( 
.A(n_4972),
.B(n_4988),
.C(n_4965),
.D(n_5034),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_L g5078 ( 
.A(n_5033),
.B(n_364),
.Y(n_5078)
);

AND2x2_ASAP7_75t_SL g5079 ( 
.A(n_4978),
.B(n_365),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_4969),
.B(n_366),
.Y(n_5080)
);

NAND3xp33_ASAP7_75t_L g5081 ( 
.A(n_5007),
.B(n_366),
.C(n_367),
.Y(n_5081)
);

AND2x2_ASAP7_75t_L g5082 ( 
.A(n_4994),
.B(n_368),
.Y(n_5082)
);

AND2x2_ASAP7_75t_L g5083 ( 
.A(n_5007),
.B(n_369),
.Y(n_5083)
);

NAND3xp33_ASAP7_75t_L g5084 ( 
.A(n_5007),
.B(n_369),
.C(n_370),
.Y(n_5084)
);

NAND2xp5_ASAP7_75t_L g5085 ( 
.A(n_4969),
.B(n_5021),
.Y(n_5085)
);

AND2x2_ASAP7_75t_L g5086 ( 
.A(n_5007),
.B(n_371),
.Y(n_5086)
);

OAI22xp5_ASAP7_75t_L g5087 ( 
.A1(n_5031),
.A2(n_375),
.B1(n_372),
.B2(n_373),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_5021),
.B(n_373),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_5052),
.Y(n_5089)
);

AND2x2_ASAP7_75t_L g5090 ( 
.A(n_5051),
.B(n_5017),
.Y(n_5090)
);

AND2x2_ASAP7_75t_L g5091 ( 
.A(n_5041),
.B(n_5017),
.Y(n_5091)
);

INVx2_ASAP7_75t_L g5092 ( 
.A(n_5079),
.Y(n_5092)
);

NOR3xp33_ASAP7_75t_L g5093 ( 
.A(n_5077),
.B(n_4999),
.C(n_4995),
.Y(n_5093)
);

AND2x2_ASAP7_75t_L g5094 ( 
.A(n_5041),
.B(n_5017),
.Y(n_5094)
);

AND2x2_ASAP7_75t_L g5095 ( 
.A(n_5044),
.B(n_5017),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_5043),
.Y(n_5096)
);

OAI33xp33_ASAP7_75t_L g5097 ( 
.A1(n_5075),
.A2(n_4995),
.A3(n_4991),
.B1(n_5018),
.B2(n_5024),
.B3(n_4999),
.Y(n_5097)
);

CKINVDCx16_ASAP7_75t_R g5098 ( 
.A(n_5058),
.Y(n_5098)
);

OAI221xp5_ASAP7_75t_SL g5099 ( 
.A1(n_5069),
.A2(n_5031),
.B1(n_4991),
.B2(n_5029),
.C(n_4982),
.Y(n_5099)
);

OAI321xp33_ASAP7_75t_L g5100 ( 
.A1(n_5068),
.A2(n_5071),
.A3(n_5072),
.B1(n_5065),
.B2(n_5059),
.C(n_5040),
.Y(n_5100)
);

INVx3_ASAP7_75t_L g5101 ( 
.A(n_5047),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_5085),
.Y(n_5102)
);

NOR3xp33_ASAP7_75t_SL g5103 ( 
.A(n_5054),
.B(n_5024),
.C(n_4981),
.Y(n_5103)
);

OR2x2_ASAP7_75t_L g5104 ( 
.A(n_5042),
.B(n_4980),
.Y(n_5104)
);

INVx4_ASAP7_75t_L g5105 ( 
.A(n_5083),
.Y(n_5105)
);

AOI31xp33_ASAP7_75t_L g5106 ( 
.A1(n_5044),
.A2(n_4980),
.A3(n_5020),
.B(n_4998),
.Y(n_5106)
);

AO21x2_ASAP7_75t_L g5107 ( 
.A1(n_5074),
.A2(n_4984),
.B(n_5026),
.Y(n_5107)
);

OR2x2_ASAP7_75t_L g5108 ( 
.A(n_5046),
.B(n_4998),
.Y(n_5108)
);

AO21x2_ASAP7_75t_L g5109 ( 
.A1(n_5083),
.A2(n_4984),
.B(n_5026),
.Y(n_5109)
);

NAND3xp33_ASAP7_75t_SL g5110 ( 
.A(n_5039),
.B(n_5009),
.C(n_5012),
.Y(n_5110)
);

AOI221xp5_ASAP7_75t_L g5111 ( 
.A1(n_5067),
.A2(n_4983),
.B1(n_5018),
.B2(n_5015),
.C(n_4976),
.Y(n_5111)
);

AND2x2_ASAP7_75t_L g5112 ( 
.A(n_5056),
.B(n_5017),
.Y(n_5112)
);

NAND2xp5_ASAP7_75t_SL g5113 ( 
.A(n_5053),
.B(n_5003),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_5086),
.B(n_5079),
.Y(n_5114)
);

NOR2xp33_ASAP7_75t_L g5115 ( 
.A(n_5082),
.B(n_5014),
.Y(n_5115)
);

NAND2xp5_ASAP7_75t_L g5116 ( 
.A(n_5086),
.B(n_5014),
.Y(n_5116)
);

AND2x2_ASAP7_75t_L g5117 ( 
.A(n_5047),
.B(n_4992),
.Y(n_5117)
);

INVx3_ASAP7_75t_L g5118 ( 
.A(n_5082),
.Y(n_5118)
);

AND2x4_ASAP7_75t_SL g5119 ( 
.A(n_5066),
.B(n_5023),
.Y(n_5119)
);

OAI21xp5_ASAP7_75t_L g5120 ( 
.A1(n_5081),
.A2(n_5003),
.B(n_5019),
.Y(n_5120)
);

OR2x2_ASAP7_75t_L g5121 ( 
.A(n_5049),
.B(n_5006),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_5078),
.Y(n_5122)
);

AND2x4_ASAP7_75t_L g5123 ( 
.A(n_5048),
.B(n_5038),
.Y(n_5123)
);

NAND2xp5_ASAP7_75t_L g5124 ( 
.A(n_5118),
.B(n_5062),
.Y(n_5124)
);

AND2x4_ASAP7_75t_SL g5125 ( 
.A(n_5091),
.B(n_5094),
.Y(n_5125)
);

NOR2xp33_ASAP7_75t_L g5126 ( 
.A(n_5098),
.B(n_5055),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_5118),
.Y(n_5127)
);

OR2x2_ASAP7_75t_L g5128 ( 
.A(n_5101),
.B(n_5050),
.Y(n_5128)
);

NAND2xp5_ASAP7_75t_L g5129 ( 
.A(n_5118),
.B(n_5062),
.Y(n_5129)
);

INVx1_ASAP7_75t_L g5130 ( 
.A(n_5119),
.Y(n_5130)
);

INVx2_ASAP7_75t_L g5131 ( 
.A(n_5107),
.Y(n_5131)
);

OR2x2_ASAP7_75t_L g5132 ( 
.A(n_5101),
.B(n_5080),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_5119),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_5101),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_SL g5135 ( 
.A(n_5103),
.B(n_5003),
.Y(n_5135)
);

AND2x2_ASAP7_75t_L g5136 ( 
.A(n_5112),
.B(n_4992),
.Y(n_5136)
);

AND2x2_ASAP7_75t_L g5137 ( 
.A(n_5091),
.B(n_5094),
.Y(n_5137)
);

AND2x2_ASAP7_75t_L g5138 ( 
.A(n_5095),
.B(n_4964),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_5107),
.Y(n_5139)
);

OR2x2_ASAP7_75t_L g5140 ( 
.A(n_5104),
.B(n_5088),
.Y(n_5140)
);

AND2x4_ASAP7_75t_L g5141 ( 
.A(n_5090),
.B(n_5038),
.Y(n_5141)
);

AND2x2_ASAP7_75t_L g5142 ( 
.A(n_5117),
.B(n_4964),
.Y(n_5142)
);

NAND2xp5_ASAP7_75t_L g5143 ( 
.A(n_5105),
.B(n_5019),
.Y(n_5143)
);

AND2x2_ASAP7_75t_L g5144 ( 
.A(n_5117),
.B(n_4979),
.Y(n_5144)
);

OR2x2_ASAP7_75t_L g5145 ( 
.A(n_5105),
.B(n_5108),
.Y(n_5145)
);

NAND2x1p5_ASAP7_75t_L g5146 ( 
.A(n_5113),
.B(n_5003),
.Y(n_5146)
);

BUFx3_ASAP7_75t_L g5147 ( 
.A(n_5105),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_5109),
.Y(n_5148)
);

AND2x2_ASAP7_75t_L g5149 ( 
.A(n_5103),
.B(n_4979),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_5131),
.Y(n_5150)
);

INVx2_ASAP7_75t_L g5151 ( 
.A(n_5137),
.Y(n_5151)
);

NAND4xp25_ASAP7_75t_SL g5152 ( 
.A(n_5149),
.B(n_5093),
.C(n_5116),
.D(n_5111),
.Y(n_5152)
);

AND2x2_ASAP7_75t_L g5153 ( 
.A(n_5137),
.B(n_5142),
.Y(n_5153)
);

AND2x2_ASAP7_75t_L g5154 ( 
.A(n_5142),
.B(n_5123),
.Y(n_5154)
);

NAND2xp5_ASAP7_75t_L g5155 ( 
.A(n_5144),
.B(n_5115),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_L g5156 ( 
.A(n_5144),
.B(n_5136),
.Y(n_5156)
);

INVx1_ASAP7_75t_SL g5157 ( 
.A(n_5125),
.Y(n_5157)
);

AND2x2_ASAP7_75t_L g5158 ( 
.A(n_5125),
.B(n_5123),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_5136),
.B(n_5115),
.Y(n_5159)
);

OR2x2_ASAP7_75t_L g5160 ( 
.A(n_5143),
.B(n_5096),
.Y(n_5160)
);

OR2x2_ASAP7_75t_L g5161 ( 
.A(n_5128),
.B(n_5089),
.Y(n_5161)
);

OR2x2_ASAP7_75t_L g5162 ( 
.A(n_5145),
.B(n_5121),
.Y(n_5162)
);

OR2x2_ASAP7_75t_L g5163 ( 
.A(n_5124),
.B(n_5102),
.Y(n_5163)
);

NAND2xp5_ASAP7_75t_L g5164 ( 
.A(n_5138),
.B(n_5092),
.Y(n_5164)
);

AND2x2_ASAP7_75t_L g5165 ( 
.A(n_5138),
.B(n_5123),
.Y(n_5165)
);

AOI21xp33_ASAP7_75t_SL g5166 ( 
.A1(n_5135),
.A2(n_5106),
.B(n_5113),
.Y(n_5166)
);

NAND2xp5_ASAP7_75t_L g5167 ( 
.A(n_5130),
.B(n_5092),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_5141),
.B(n_5016),
.Y(n_5168)
);

OR2x6_ASAP7_75t_L g5169 ( 
.A(n_5147),
.B(n_5133),
.Y(n_5169)
);

AND2x4_ASAP7_75t_L g5170 ( 
.A(n_5141),
.B(n_5147),
.Y(n_5170)
);

NOR4xp25_ASAP7_75t_SL g5171 ( 
.A(n_5166),
.B(n_5135),
.C(n_5099),
.D(n_5100),
.Y(n_5171)
);

NAND2xp5_ASAP7_75t_L g5172 ( 
.A(n_5153),
.B(n_5149),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_5154),
.B(n_5126),
.Y(n_5173)
);

NOR2x1_ASAP7_75t_L g5174 ( 
.A(n_5170),
.B(n_5131),
.Y(n_5174)
);

NAND2xp5_ASAP7_75t_L g5175 ( 
.A(n_5165),
.B(n_5126),
.Y(n_5175)
);

NOR4xp25_ASAP7_75t_SL g5176 ( 
.A(n_5166),
.B(n_5148),
.C(n_5127),
.D(n_5134),
.Y(n_5176)
);

AOI22xp5_ASAP7_75t_L g5177 ( 
.A1(n_5152),
.A2(n_5139),
.B1(n_5110),
.B2(n_5114),
.Y(n_5177)
);

NOR2xp33_ASAP7_75t_L g5178 ( 
.A(n_5156),
.B(n_5141),
.Y(n_5178)
);

OAI221xp5_ASAP7_75t_L g5179 ( 
.A1(n_5164),
.A2(n_5120),
.B1(n_5139),
.B2(n_5039),
.C(n_5129),
.Y(n_5179)
);

NOR2xp33_ASAP7_75t_R g5180 ( 
.A(n_5157),
.B(n_5132),
.Y(n_5180)
);

INVx2_ASAP7_75t_L g5181 ( 
.A(n_5151),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_5157),
.B(n_5122),
.Y(n_5182)
);

NOR2xp33_ASAP7_75t_L g5183 ( 
.A(n_5170),
.B(n_5097),
.Y(n_5183)
);

INVx3_ASAP7_75t_L g5184 ( 
.A(n_5169),
.Y(n_5184)
);

NOR2x1_ASAP7_75t_L g5185 ( 
.A(n_5174),
.B(n_5169),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_5184),
.B(n_5158),
.Y(n_5186)
);

INVx2_ASAP7_75t_L g5187 ( 
.A(n_5175),
.Y(n_5187)
);

AND2x2_ASAP7_75t_L g5188 ( 
.A(n_5178),
.B(n_5168),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_L g5189 ( 
.A(n_5173),
.B(n_5155),
.Y(n_5189)
);

NAND2xp5_ASAP7_75t_L g5190 ( 
.A(n_5177),
.B(n_5159),
.Y(n_5190)
);

AND3x2_ASAP7_75t_L g5191 ( 
.A(n_5181),
.B(n_5150),
.C(n_5167),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_5182),
.Y(n_5192)
);

OR2x2_ASAP7_75t_L g5193 ( 
.A(n_5172),
.B(n_5162),
.Y(n_5193)
);

AND2x2_ASAP7_75t_L g5194 ( 
.A(n_5180),
.B(n_5146),
.Y(n_5194)
);

AOI22xp33_ASAP7_75t_L g5195 ( 
.A1(n_5183),
.A2(n_5109),
.B1(n_5150),
.B2(n_5015),
.Y(n_5195)
);

NAND2xp5_ASAP7_75t_L g5196 ( 
.A(n_5176),
.B(n_5140),
.Y(n_5196)
);

OR2x6_ASAP7_75t_L g5197 ( 
.A(n_5171),
.B(n_5161),
.Y(n_5197)
);

NOR2xp33_ASAP7_75t_L g5198 ( 
.A(n_5179),
.B(n_5146),
.Y(n_5198)
);

AND2x4_ASAP7_75t_L g5199 ( 
.A(n_5184),
.B(n_5163),
.Y(n_5199)
);

INVx1_ASAP7_75t_L g5200 ( 
.A(n_5174),
.Y(n_5200)
);

HB1xp67_ASAP7_75t_L g5201 ( 
.A(n_5197),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_5193),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5199),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_5187),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_5191),
.Y(n_5205)
);

AOI22xp33_ASAP7_75t_L g5206 ( 
.A1(n_5195),
.A2(n_5084),
.B1(n_5070),
.B2(n_5073),
.Y(n_5206)
);

AND2x2_ASAP7_75t_L g5207 ( 
.A(n_5197),
.B(n_5160),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_5189),
.Y(n_5208)
);

NAND2xp5_ASAP7_75t_L g5209 ( 
.A(n_5185),
.B(n_5006),
.Y(n_5209)
);

AND2x2_ASAP7_75t_L g5210 ( 
.A(n_5188),
.B(n_4979),
.Y(n_5210)
);

AO22x1_ASAP7_75t_L g5211 ( 
.A1(n_5194),
.A2(n_5087),
.B1(n_5045),
.B2(n_5003),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5200),
.Y(n_5212)
);

AOI22xp33_ASAP7_75t_L g5213 ( 
.A1(n_5201),
.A2(n_5196),
.B1(n_5192),
.B2(n_5190),
.Y(n_5213)
);

AOI22xp5_ASAP7_75t_L g5214 ( 
.A1(n_5201),
.A2(n_5198),
.B1(n_5186),
.B2(n_4973),
.Y(n_5214)
);

OAI21xp5_ASAP7_75t_L g5215 ( 
.A1(n_5207),
.A2(n_5210),
.B(n_5202),
.Y(n_5215)
);

OAI221xp5_ASAP7_75t_L g5216 ( 
.A1(n_5206),
.A2(n_5064),
.B1(n_5063),
.B2(n_5057),
.C(n_4983),
.Y(n_5216)
);

AND2x2_ASAP7_75t_L g5217 ( 
.A(n_5203),
.B(n_4979),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_5208),
.Y(n_5218)
);

AOI21xp33_ASAP7_75t_SL g5219 ( 
.A1(n_5205),
.A2(n_4986),
.B(n_4985),
.Y(n_5219)
);

AOI22xp5_ASAP7_75t_L g5220 ( 
.A1(n_5204),
.A2(n_4973),
.B1(n_4976),
.B2(n_4975),
.Y(n_5220)
);

OAI21xp5_ASAP7_75t_L g5221 ( 
.A1(n_5209),
.A2(n_4973),
.B(n_5060),
.Y(n_5221)
);

OR2x2_ASAP7_75t_L g5222 ( 
.A(n_5215),
.B(n_5212),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_5217),
.Y(n_5223)
);

AOI21xp5_ASAP7_75t_L g5224 ( 
.A1(n_5213),
.A2(n_5211),
.B(n_5206),
.Y(n_5224)
);

OAI21xp33_ASAP7_75t_L g5225 ( 
.A1(n_5214),
.A2(n_4973),
.B(n_5061),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_5220),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_5218),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_5221),
.Y(n_5228)
);

INVx1_ASAP7_75t_SL g5229 ( 
.A(n_5219),
.Y(n_5229)
);

AOI322xp5_ASAP7_75t_L g5230 ( 
.A1(n_5229),
.A2(n_5225),
.A3(n_5223),
.B1(n_5227),
.B2(n_5226),
.C1(n_5228),
.C2(n_5216),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_5224),
.B(n_4985),
.Y(n_5231)
);

AOI32xp33_ASAP7_75t_L g5232 ( 
.A1(n_5222),
.A2(n_5063),
.A3(n_4990),
.B1(n_4986),
.B2(n_5008),
.Y(n_5232)
);

NAND2xp5_ASAP7_75t_L g5233 ( 
.A(n_5223),
.B(n_4990),
.Y(n_5233)
);

XNOR2x1_ASAP7_75t_L g5234 ( 
.A(n_5222),
.B(n_4975),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_5222),
.Y(n_5235)
);

OAI21xp33_ASAP7_75t_SL g5236 ( 
.A1(n_5222),
.A2(n_4967),
.B(n_4966),
.Y(n_5236)
);

NAND3xp33_ASAP7_75t_L g5237 ( 
.A(n_5224),
.B(n_5076),
.C(n_5037),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_5223),
.B(n_5023),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5222),
.Y(n_5239)
);

AOI21xp33_ASAP7_75t_SL g5240 ( 
.A1(n_5222),
.A2(n_4981),
.B(n_5001),
.Y(n_5240)
);

OAI22xp5_ASAP7_75t_L g5241 ( 
.A1(n_5222),
.A2(n_4967),
.B1(n_4966),
.B2(n_4974),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_5222),
.Y(n_5242)
);

NAND2xp5_ASAP7_75t_L g5243 ( 
.A(n_5223),
.B(n_5008),
.Y(n_5243)
);

NAND2xp5_ASAP7_75t_L g5244 ( 
.A(n_5223),
.B(n_5001),
.Y(n_5244)
);

XNOR2xp5_ASAP7_75t_L g5245 ( 
.A(n_5223),
.B(n_5032),
.Y(n_5245)
);

NAND2xp5_ASAP7_75t_L g5246 ( 
.A(n_5223),
.B(n_5004),
.Y(n_5246)
);

NAND2xp5_ASAP7_75t_SL g5247 ( 
.A(n_5224),
.B(n_4974),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5243),
.Y(n_5248)
);

INVxp33_ASAP7_75t_SL g5249 ( 
.A(n_5245),
.Y(n_5249)
);

CKINVDCx6p67_ASAP7_75t_R g5250 ( 
.A(n_5235),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_5238),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_5234),
.Y(n_5252)
);

INVx2_ASAP7_75t_L g5253 ( 
.A(n_5239),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_5242),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_5244),
.Y(n_5255)
);

INVx1_ASAP7_75t_SL g5256 ( 
.A(n_5246),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_5241),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5247),
.Y(n_5258)
);

NOR2xp33_ASAP7_75t_L g5259 ( 
.A(n_5240),
.B(n_5004),
.Y(n_5259)
);

HB1xp67_ASAP7_75t_L g5260 ( 
.A(n_5231),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_5233),
.Y(n_5261)
);

INVxp67_ASAP7_75t_L g5262 ( 
.A(n_5237),
.Y(n_5262)
);

INVx1_ASAP7_75t_SL g5263 ( 
.A(n_5230),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_5236),
.Y(n_5264)
);

INVx2_ASAP7_75t_L g5265 ( 
.A(n_5232),
.Y(n_5265)
);

HB1xp67_ASAP7_75t_L g5266 ( 
.A(n_5245),
.Y(n_5266)
);

HB1xp67_ASAP7_75t_L g5267 ( 
.A(n_5235),
.Y(n_5267)
);

INVx1_ASAP7_75t_SL g5268 ( 
.A(n_5234),
.Y(n_5268)
);

INVx1_ASAP7_75t_SL g5269 ( 
.A(n_5234),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_5243),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_5243),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_5243),
.Y(n_5272)
);

INVx1_ASAP7_75t_L g5273 ( 
.A(n_5243),
.Y(n_5273)
);

AOI221xp5_ASAP7_75t_L g5274 ( 
.A1(n_5267),
.A2(n_5015),
.B1(n_5032),
.B2(n_5037),
.C(n_4989),
.Y(n_5274)
);

OAI21xp5_ASAP7_75t_SL g5275 ( 
.A1(n_5267),
.A2(n_4971),
.B(n_5015),
.Y(n_5275)
);

XNOR2x1_ASAP7_75t_L g5276 ( 
.A(n_5263),
.B(n_4989),
.Y(n_5276)
);

OR2x2_ASAP7_75t_L g5277 ( 
.A(n_5250),
.B(n_5256),
.Y(n_5277)
);

AOI21xp5_ASAP7_75t_L g5278 ( 
.A1(n_5258),
.A2(n_5016),
.B(n_4971),
.Y(n_5278)
);

INVx2_ASAP7_75t_L g5279 ( 
.A(n_5253),
.Y(n_5279)
);

OAI22xp33_ASAP7_75t_L g5280 ( 
.A1(n_5254),
.A2(n_4987),
.B1(n_379),
.B2(n_376),
.Y(n_5280)
);

OAI21xp5_ASAP7_75t_L g5281 ( 
.A1(n_5262),
.A2(n_4987),
.B(n_376),
.Y(n_5281)
);

OAI221xp5_ASAP7_75t_L g5282 ( 
.A1(n_5262),
.A2(n_5259),
.B1(n_5264),
.B2(n_5268),
.C(n_5269),
.Y(n_5282)
);

NAND5xp2_ASAP7_75t_L g5283 ( 
.A(n_5249),
.B(n_378),
.C(n_381),
.D(n_382),
.E(n_383),
.Y(n_5283)
);

AOI21xp33_ASAP7_75t_L g5284 ( 
.A1(n_5260),
.A2(n_378),
.B(n_381),
.Y(n_5284)
);

AOI22xp5_ASAP7_75t_L g5285 ( 
.A1(n_5252),
.A2(n_387),
.B1(n_384),
.B2(n_385),
.Y(n_5285)
);

INVx1_ASAP7_75t_L g5286 ( 
.A(n_5260),
.Y(n_5286)
);

OAI21xp33_ASAP7_75t_L g5287 ( 
.A1(n_5248),
.A2(n_387),
.B(n_388),
.Y(n_5287)
);

OAI22xp5_ASAP7_75t_L g5288 ( 
.A1(n_5261),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_5266),
.Y(n_5289)
);

OAI31xp33_ASAP7_75t_L g5290 ( 
.A1(n_5270),
.A2(n_392),
.A3(n_389),
.B(n_391),
.Y(n_5290)
);

OAI21xp33_ASAP7_75t_L g5291 ( 
.A1(n_5271),
.A2(n_391),
.B(n_392),
.Y(n_5291)
);

OAI211xp5_ASAP7_75t_SL g5292 ( 
.A1(n_5272),
.A2(n_397),
.B(n_394),
.C(n_396),
.Y(n_5292)
);

NAND2xp5_ASAP7_75t_L g5293 ( 
.A(n_5273),
.B(n_397),
.Y(n_5293)
);

OAI211xp5_ASAP7_75t_SL g5294 ( 
.A1(n_5251),
.A2(n_400),
.B(n_398),
.C(n_399),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_5255),
.B(n_399),
.Y(n_5295)
);

AOI22xp5_ASAP7_75t_L g5296 ( 
.A1(n_5265),
.A2(n_404),
.B1(n_401),
.B2(n_403),
.Y(n_5296)
);

AOI22xp5_ASAP7_75t_L g5297 ( 
.A1(n_5257),
.A2(n_404),
.B1(n_401),
.B2(n_403),
.Y(n_5297)
);

INVx2_ASAP7_75t_L g5298 ( 
.A(n_5267),
.Y(n_5298)
);

AOI321xp33_ASAP7_75t_L g5299 ( 
.A1(n_5259),
.A2(n_405),
.A3(n_407),
.B1(n_408),
.B2(n_409),
.C(n_410),
.Y(n_5299)
);

NAND2xp33_ASAP7_75t_SL g5300 ( 
.A(n_5258),
.B(n_407),
.Y(n_5300)
);

AOI221xp5_ASAP7_75t_L g5301 ( 
.A1(n_5298),
.A2(n_408),
.B1(n_409),
.B2(n_410),
.C(n_411),
.Y(n_5301)
);

AOI31xp33_ASAP7_75t_L g5302 ( 
.A1(n_5277),
.A2(n_411),
.A3(n_412),
.B(n_413),
.Y(n_5302)
);

OAI211xp5_ASAP7_75t_SL g5303 ( 
.A1(n_5282),
.A2(n_412),
.B(n_415),
.C(n_416),
.Y(n_5303)
);

AOI21xp5_ASAP7_75t_L g5304 ( 
.A1(n_5286),
.A2(n_415),
.B(n_417),
.Y(n_5304)
);

NAND2xp5_ASAP7_75t_L g5305 ( 
.A(n_5275),
.B(n_418),
.Y(n_5305)
);

OAI211xp5_ASAP7_75t_L g5306 ( 
.A1(n_5296),
.A2(n_419),
.B(n_420),
.C(n_421),
.Y(n_5306)
);

AOI22xp5_ASAP7_75t_L g5307 ( 
.A1(n_5279),
.A2(n_422),
.B1(n_423),
.B2(n_425),
.Y(n_5307)
);

OAI221xp5_ASAP7_75t_L g5308 ( 
.A1(n_5278),
.A2(n_5289),
.B1(n_5290),
.B2(n_5287),
.C(n_5291),
.Y(n_5308)
);

AOI211x1_ASAP7_75t_SL g5309 ( 
.A1(n_5281),
.A2(n_426),
.B(n_427),
.C(n_430),
.Y(n_5309)
);

AOI21xp5_ASAP7_75t_L g5310 ( 
.A1(n_5293),
.A2(n_427),
.B(n_430),
.Y(n_5310)
);

INVx2_ASAP7_75t_L g5311 ( 
.A(n_5276),
.Y(n_5311)
);

INVx1_ASAP7_75t_SL g5312 ( 
.A(n_5300),
.Y(n_5312)
);

AOI331xp33_ASAP7_75t_L g5313 ( 
.A1(n_5299),
.A2(n_431),
.A3(n_432),
.B1(n_434),
.B2(n_436),
.B3(n_437),
.C1(n_438),
.Y(n_5313)
);

AOI22xp5_ASAP7_75t_L g5314 ( 
.A1(n_5285),
.A2(n_431),
.B1(n_432),
.B2(n_436),
.Y(n_5314)
);

NOR2xp33_ASAP7_75t_SL g5315 ( 
.A(n_5284),
.B(n_5295),
.Y(n_5315)
);

OAI221xp5_ASAP7_75t_L g5316 ( 
.A1(n_5297),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.C(n_441),
.Y(n_5316)
);

OAI21xp5_ASAP7_75t_L g5317 ( 
.A1(n_5280),
.A2(n_441),
.B(n_442),
.Y(n_5317)
);

CKINVDCx5p33_ASAP7_75t_R g5318 ( 
.A(n_5288),
.Y(n_5318)
);

O2A1O1Ixp33_ASAP7_75t_L g5319 ( 
.A1(n_5292),
.A2(n_442),
.B(n_443),
.C(n_446),
.Y(n_5319)
);

O2A1O1Ixp33_ASAP7_75t_L g5320 ( 
.A1(n_5294),
.A2(n_443),
.B(n_447),
.C(n_448),
.Y(n_5320)
);

AOI221x1_ASAP7_75t_SL g5321 ( 
.A1(n_5283),
.A2(n_447),
.B1(n_448),
.B2(n_449),
.C(n_450),
.Y(n_5321)
);

OAI21xp5_ASAP7_75t_SL g5322 ( 
.A1(n_5274),
.A2(n_449),
.B(n_450),
.Y(n_5322)
);

OAI22xp5_ASAP7_75t_L g5323 ( 
.A1(n_5277),
.A2(n_451),
.B1(n_452),
.B2(n_455),
.Y(n_5323)
);

OAI211xp5_ASAP7_75t_SL g5324 ( 
.A1(n_5282),
.A2(n_451),
.B(n_452),
.C(n_456),
.Y(n_5324)
);

OA22x2_ASAP7_75t_L g5325 ( 
.A1(n_5322),
.A2(n_456),
.B1(n_458),
.B2(n_459),
.Y(n_5325)
);

OR2x2_ASAP7_75t_L g5326 ( 
.A(n_5312),
.B(n_459),
.Y(n_5326)
);

OAI211xp5_ASAP7_75t_SL g5327 ( 
.A1(n_5311),
.A2(n_5305),
.B(n_5308),
.C(n_5309),
.Y(n_5327)
);

OAI211xp5_ASAP7_75t_L g5328 ( 
.A1(n_5304),
.A2(n_5324),
.B(n_5303),
.C(n_5314),
.Y(n_5328)
);

NOR2xp67_ASAP7_75t_L g5329 ( 
.A(n_5306),
.B(n_460),
.Y(n_5329)
);

OAI221xp5_ASAP7_75t_SL g5330 ( 
.A1(n_5319),
.A2(n_5320),
.B1(n_5310),
.B2(n_5316),
.C(n_5307),
.Y(n_5330)
);

OAI22xp33_ASAP7_75t_L g5331 ( 
.A1(n_5302),
.A2(n_460),
.B1(n_461),
.B2(n_462),
.Y(n_5331)
);

AOI222xp33_ASAP7_75t_L g5332 ( 
.A1(n_5317),
.A2(n_461),
.B1(n_463),
.B2(n_465),
.C1(n_466),
.C2(n_467),
.Y(n_5332)
);

AOI31xp33_ASAP7_75t_L g5333 ( 
.A1(n_5318),
.A2(n_463),
.A3(n_465),
.B(n_466),
.Y(n_5333)
);

INVx1_ASAP7_75t_SL g5334 ( 
.A(n_5315),
.Y(n_5334)
);

NOR2x1_ASAP7_75t_L g5335 ( 
.A(n_5323),
.B(n_5313),
.Y(n_5335)
);

XOR2xp5_ASAP7_75t_L g5336 ( 
.A(n_5321),
.B(n_467),
.Y(n_5336)
);

O2A1O1Ixp5_ASAP7_75t_SL g5337 ( 
.A1(n_5301),
.A2(n_468),
.B(n_470),
.C(n_471),
.Y(n_5337)
);

OAI21xp33_ASAP7_75t_SL g5338 ( 
.A1(n_5305),
.A2(n_471),
.B(n_472),
.Y(n_5338)
);

INVxp33_ASAP7_75t_L g5339 ( 
.A(n_5311),
.Y(n_5339)
);

AOI221x1_ASAP7_75t_L g5340 ( 
.A1(n_5305),
.A2(n_472),
.B1(n_473),
.B2(n_474),
.C(n_475),
.Y(n_5340)
);

OAI211xp5_ASAP7_75t_L g5341 ( 
.A1(n_5305),
.A2(n_474),
.B(n_475),
.C(n_477),
.Y(n_5341)
);

AOI211xp5_ASAP7_75t_L g5342 ( 
.A1(n_5308),
.A2(n_477),
.B(n_478),
.C(n_479),
.Y(n_5342)
);

INVxp67_ASAP7_75t_SL g5343 ( 
.A(n_5326),
.Y(n_5343)
);

AO22x2_ASAP7_75t_L g5344 ( 
.A1(n_5334),
.A2(n_478),
.B1(n_479),
.B2(n_480),
.Y(n_5344)
);

HB1xp67_ASAP7_75t_L g5345 ( 
.A(n_5336),
.Y(n_5345)
);

NAND2xp5_ASAP7_75t_L g5346 ( 
.A(n_5339),
.B(n_480),
.Y(n_5346)
);

AND2x2_ASAP7_75t_L g5347 ( 
.A(n_5335),
.B(n_5329),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_5333),
.Y(n_5348)
);

NOR2x1_ASAP7_75t_L g5349 ( 
.A(n_5327),
.B(n_481),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5325),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_5340),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5338),
.Y(n_5352)
);

INVx1_ASAP7_75t_L g5353 ( 
.A(n_5341),
.Y(n_5353)
);

NAND2xp5_ASAP7_75t_L g5354 ( 
.A(n_5331),
.B(n_482),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_5328),
.Y(n_5355)
);

AOI22xp5_ASAP7_75t_L g5356 ( 
.A1(n_5332),
.A2(n_482),
.B1(n_483),
.B2(n_484),
.Y(n_5356)
);

OAI22xp33_ASAP7_75t_L g5357 ( 
.A1(n_5342),
.A2(n_5337),
.B1(n_5330),
.B2(n_485),
.Y(n_5357)
);

NOR3xp33_ASAP7_75t_L g5358 ( 
.A(n_5343),
.B(n_483),
.C(n_484),
.Y(n_5358)
);

INVxp33_ASAP7_75t_L g5359 ( 
.A(n_5349),
.Y(n_5359)
);

AND2x4_ASAP7_75t_L g5360 ( 
.A(n_5347),
.B(n_486),
.Y(n_5360)
);

OR2x2_ASAP7_75t_L g5361 ( 
.A(n_5352),
.B(n_486),
.Y(n_5361)
);

INVx2_ASAP7_75t_SL g5362 ( 
.A(n_5351),
.Y(n_5362)
);

OR2x2_ASAP7_75t_L g5363 ( 
.A(n_5355),
.B(n_487),
.Y(n_5363)
);

AOI222xp33_ASAP7_75t_L g5364 ( 
.A1(n_5350),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.C1(n_490),
.C2(n_491),
.Y(n_5364)
);

INVx2_ASAP7_75t_L g5365 ( 
.A(n_5344),
.Y(n_5365)
);

BUFx6f_ASAP7_75t_L g5366 ( 
.A(n_5346),
.Y(n_5366)
);

OAI211xp5_ASAP7_75t_SL g5367 ( 
.A1(n_5348),
.A2(n_488),
.B(n_490),
.C(n_491),
.Y(n_5367)
);

INVx1_ASAP7_75t_SL g5368 ( 
.A(n_5344),
.Y(n_5368)
);

OAI211xp5_ASAP7_75t_L g5369 ( 
.A1(n_5345),
.A2(n_492),
.B(n_493),
.C(n_494),
.Y(n_5369)
);

NOR2xp67_ASAP7_75t_SL g5370 ( 
.A(n_5353),
.B(n_492),
.Y(n_5370)
);

NOR2xp33_ASAP7_75t_R g5371 ( 
.A(n_5362),
.B(n_5354),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_L g5372 ( 
.A(n_5368),
.B(n_5365),
.Y(n_5372)
);

NOR2xp33_ASAP7_75t_R g5373 ( 
.A(n_5363),
.B(n_5357),
.Y(n_5373)
);

NAND2xp5_ASAP7_75t_SL g5374 ( 
.A(n_5359),
.B(n_5366),
.Y(n_5374)
);

NAND2xp5_ASAP7_75t_SL g5375 ( 
.A(n_5366),
.B(n_5356),
.Y(n_5375)
);

NAND3xp33_ASAP7_75t_L g5376 ( 
.A(n_5361),
.B(n_493),
.C(n_494),
.Y(n_5376)
);

NOR3xp33_ASAP7_75t_SL g5377 ( 
.A(n_5367),
.B(n_495),
.C(n_496),
.Y(n_5377)
);

NAND2xp33_ASAP7_75t_SL g5378 ( 
.A(n_5370),
.B(n_497),
.Y(n_5378)
);

NAND3xp33_ASAP7_75t_SL g5379 ( 
.A(n_5358),
.B(n_498),
.C(n_500),
.Y(n_5379)
);

NAND3xp33_ASAP7_75t_SL g5380 ( 
.A(n_5369),
.B(n_500),
.C(n_501),
.Y(n_5380)
);

AOI221xp5_ASAP7_75t_L g5381 ( 
.A1(n_5374),
.A2(n_5360),
.B1(n_5364),
.B2(n_503),
.C(n_505),
.Y(n_5381)
);

NAND4xp25_ASAP7_75t_SL g5382 ( 
.A(n_5372),
.B(n_501),
.C(n_502),
.D(n_506),
.Y(n_5382)
);

A2O1A1Ixp33_ASAP7_75t_L g5383 ( 
.A1(n_5376),
.A2(n_508),
.B(n_509),
.C(n_510),
.Y(n_5383)
);

AOI211xp5_ASAP7_75t_L g5384 ( 
.A1(n_5375),
.A2(n_509),
.B(n_510),
.C(n_511),
.Y(n_5384)
);

AOI22xp5_ASAP7_75t_SL g5385 ( 
.A1(n_5378),
.A2(n_511),
.B1(n_513),
.B2(n_515),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_5373),
.Y(n_5386)
);

OA22x2_ASAP7_75t_L g5387 ( 
.A1(n_5371),
.A2(n_515),
.B1(n_516),
.B2(n_517),
.Y(n_5387)
);

INVx1_ASAP7_75t_SL g5388 ( 
.A(n_5386),
.Y(n_5388)
);

AOI21xp5_ASAP7_75t_L g5389 ( 
.A1(n_5385),
.A2(n_5379),
.B(n_5380),
.Y(n_5389)
);

XNOR2xp5_ASAP7_75t_L g5390 ( 
.A(n_5381),
.B(n_5377),
.Y(n_5390)
);

OAI21xp5_ASAP7_75t_L g5391 ( 
.A1(n_5388),
.A2(n_5383),
.B(n_5382),
.Y(n_5391)
);

AO21x1_ASAP7_75t_L g5392 ( 
.A1(n_5389),
.A2(n_5384),
.B(n_5387),
.Y(n_5392)
);

XNOR2xp5_ASAP7_75t_L g5393 ( 
.A(n_5391),
.B(n_5390),
.Y(n_5393)
);

INVx1_ASAP7_75t_L g5394 ( 
.A(n_5392),
.Y(n_5394)
);

AOI22xp5_ASAP7_75t_L g5395 ( 
.A1(n_5394),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.Y(n_5395)
);

OAI22xp5_ASAP7_75t_L g5396 ( 
.A1(n_5393),
.A2(n_519),
.B1(n_520),
.B2(n_521),
.Y(n_5396)
);

OAI22xp5_ASAP7_75t_L g5397 ( 
.A1(n_5394),
.A2(n_522),
.B1(n_523),
.B2(n_524),
.Y(n_5397)
);

AOI31xp33_ASAP7_75t_L g5398 ( 
.A1(n_5396),
.A2(n_522),
.A3(n_525),
.B(n_526),
.Y(n_5398)
);

AOI31xp33_ASAP7_75t_L g5399 ( 
.A1(n_5397),
.A2(n_526),
.A3(n_527),
.B(n_528),
.Y(n_5399)
);

AOI22xp33_ASAP7_75t_L g5400 ( 
.A1(n_5395),
.A2(n_527),
.B1(n_529),
.B2(n_533),
.Y(n_5400)
);

AOI31xp33_ASAP7_75t_L g5401 ( 
.A1(n_5396),
.A2(n_529),
.A3(n_534),
.B(n_535),
.Y(n_5401)
);

OAI21xp5_ASAP7_75t_L g5402 ( 
.A1(n_5398),
.A2(n_534),
.B(n_537),
.Y(n_5402)
);

INVx1_ASAP7_75t_L g5403 ( 
.A(n_5401),
.Y(n_5403)
);

OA22x2_ASAP7_75t_L g5404 ( 
.A1(n_5399),
.A2(n_537),
.B1(n_538),
.B2(n_539),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5400),
.Y(n_5405)
);

INVx2_ASAP7_75t_SL g5406 ( 
.A(n_5398),
.Y(n_5406)
);

OR2x6_ASAP7_75t_L g5407 ( 
.A(n_5406),
.B(n_539),
.Y(n_5407)
);

OAI22xp5_ASAP7_75t_L g5408 ( 
.A1(n_5404),
.A2(n_5403),
.B1(n_5402),
.B2(n_5405),
.Y(n_5408)
);

AOI22x1_ASAP7_75t_L g5409 ( 
.A1(n_5406),
.A2(n_540),
.B1(n_541),
.B2(n_542),
.Y(n_5409)
);

OR2x6_ASAP7_75t_L g5410 ( 
.A(n_5406),
.B(n_540),
.Y(n_5410)
);

AOI221xp5_ASAP7_75t_L g5411 ( 
.A1(n_5403),
.A2(n_542),
.B1(n_543),
.B2(n_545),
.C(n_547),
.Y(n_5411)
);

OAI21xp5_ASAP7_75t_L g5412 ( 
.A1(n_5403),
.A2(n_543),
.B(n_548),
.Y(n_5412)
);

INVx2_ASAP7_75t_L g5413 ( 
.A(n_5406),
.Y(n_5413)
);

AND2x2_ASAP7_75t_L g5414 ( 
.A(n_5406),
.B(n_549),
.Y(n_5414)
);

AOI21xp5_ASAP7_75t_L g5415 ( 
.A1(n_5406),
.A2(n_549),
.B(n_550),
.Y(n_5415)
);

AOI22xp5_ASAP7_75t_L g5416 ( 
.A1(n_5406),
.A2(n_552),
.B1(n_553),
.B2(n_554),
.Y(n_5416)
);

INVxp67_ASAP7_75t_SL g5417 ( 
.A(n_5413),
.Y(n_5417)
);

AOI321xp33_ASAP7_75t_L g5418 ( 
.A1(n_5408),
.A2(n_552),
.A3(n_554),
.B1(n_555),
.B2(n_556),
.C(n_557),
.Y(n_5418)
);

AOI21xp5_ASAP7_75t_SL g5419 ( 
.A1(n_5407),
.A2(n_555),
.B(n_558),
.Y(n_5419)
);

OAI222xp33_ASAP7_75t_L g5420 ( 
.A1(n_5410),
.A2(n_559),
.B1(n_560),
.B2(n_562),
.C1(n_563),
.C2(n_564),
.Y(n_5420)
);

AOI22xp5_ASAP7_75t_L g5421 ( 
.A1(n_5414),
.A2(n_563),
.B1(n_565),
.B2(n_567),
.Y(n_5421)
);

AOI22xp5_ASAP7_75t_L g5422 ( 
.A1(n_5412),
.A2(n_565),
.B1(n_568),
.B2(n_569),
.Y(n_5422)
);

OAI21xp5_ASAP7_75t_SL g5423 ( 
.A1(n_5415),
.A2(n_5416),
.B(n_5411),
.Y(n_5423)
);

AOI222xp33_ASAP7_75t_SL g5424 ( 
.A1(n_5409),
.A2(n_568),
.B1(n_570),
.B2(n_571),
.C1(n_572),
.C2(n_573),
.Y(n_5424)
);

AOI32xp33_ASAP7_75t_L g5425 ( 
.A1(n_5413),
.A2(n_570),
.A3(n_571),
.B1(n_573),
.B2(n_574),
.Y(n_5425)
);

INVxp67_ASAP7_75t_SL g5426 ( 
.A(n_5417),
.Y(n_5426)
);

HB1xp67_ASAP7_75t_L g5427 ( 
.A(n_5423),
.Y(n_5427)
);

OR2x2_ASAP7_75t_L g5428 ( 
.A(n_5419),
.B(n_575),
.Y(n_5428)
);

OAI222xp33_ASAP7_75t_L g5429 ( 
.A1(n_5425),
.A2(n_577),
.B1(n_578),
.B2(n_579),
.C1(n_580),
.C2(n_581),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_5422),
.Y(n_5430)
);

XOR2xp5_ASAP7_75t_L g5431 ( 
.A(n_5421),
.B(n_577),
.Y(n_5431)
);

AOI22xp33_ASAP7_75t_L g5432 ( 
.A1(n_5426),
.A2(n_5424),
.B1(n_5418),
.B2(n_5420),
.Y(n_5432)
);

AOI322xp5_ASAP7_75t_L g5433 ( 
.A1(n_5427),
.A2(n_580),
.A3(n_582),
.B1(n_583),
.B2(n_585),
.C1(n_586),
.C2(n_587),
.Y(n_5433)
);

AOI22x1_ASAP7_75t_L g5434 ( 
.A1(n_5430),
.A2(n_583),
.B1(n_586),
.B2(n_588),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5428),
.Y(n_5435)
);

AOI22xp33_ASAP7_75t_L g5436 ( 
.A1(n_5435),
.A2(n_5431),
.B1(n_5429),
.B2(n_590),
.Y(n_5436)
);

OAI221xp5_ASAP7_75t_R g5437 ( 
.A1(n_5432),
.A2(n_5434),
.B1(n_5433),
.B2(n_591),
.C(n_592),
.Y(n_5437)
);

AOI22xp33_ASAP7_75t_SL g5438 ( 
.A1(n_5437),
.A2(n_588),
.B1(n_589),
.B2(n_591),
.Y(n_5438)
);

AOI211xp5_ASAP7_75t_L g5439 ( 
.A1(n_5438),
.A2(n_5436),
.B(n_592),
.C(n_593),
.Y(n_5439)
);


endmodule