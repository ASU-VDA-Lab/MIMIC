module fake_jpeg_14498_n_431 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_431);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_431;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_46),
.B(n_56),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_47),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_48),
.B(n_50),
.Y(n_136)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_49),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_15),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_17),
.B(n_0),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_57),
.Y(n_103)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_66),
.B(n_67),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_30),
.B(n_2),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_39),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_82),
.Y(n_89)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_77),
.Y(n_131)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_23),
.B(n_3),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_88),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_31),
.B1(n_38),
.B2(n_22),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_92),
.A2(n_73),
.B(n_71),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_43),
.B1(n_22),
.B2(n_42),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_99),
.A2(n_121),
.B1(n_133),
.B2(n_60),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_26),
.B(n_40),
.C(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_102),
.B(n_124),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_74),
.A2(n_42),
.B1(n_28),
.B2(n_38),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_107),
.A2(n_113),
.B1(n_132),
.B2(n_47),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_26),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_114),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_49),
.A2(n_38),
.B1(n_34),
.B2(n_43),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_45),
.B(n_40),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_59),
.A2(n_43),
.B1(n_22),
.B2(n_23),
.Y(n_121)
);

HAxp5_ASAP7_75t_SL g122 ( 
.A(n_57),
.B(n_36),
.CON(n_122),
.SN(n_122)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_122),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_55),
.A2(n_34),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_128),
.C(n_6),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_54),
.B(n_34),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_139),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_47),
.B(n_34),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_135),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_58),
.B(n_3),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_81),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_65),
.A2(n_14),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_3),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_5),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_157),
.Y(n_201)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_145),
.Y(n_239)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_72),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_147),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_78),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_150),
.B(n_160),
.Y(n_219)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

AO22x1_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_70),
.B1(n_72),
.B2(n_51),
.Y(n_152)
);

AO22x2_ASAP7_75t_L g237 ( 
.A1(n_152),
.A2(n_165),
.B1(n_155),
.B2(n_194),
.Y(n_237)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_156),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_100),
.B(n_86),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_162),
.B(n_172),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_166),
.B1(n_175),
.B2(n_180),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_114),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_174),
.Y(n_203)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_84),
.B1(n_79),
.B2(n_69),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_169),
.B(n_189),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_89),
.B(n_77),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_103),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_98),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_176),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_7),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_182),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_7),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_97),
.B(n_7),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_135),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_13),
.C(n_11),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_191),
.C(n_182),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_11),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_94),
.B(n_11),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_91),
.A2(n_12),
.B1(n_13),
.B2(n_112),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_185),
.A2(n_123),
.B1(n_104),
.B2(n_130),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_138),
.A2(n_12),
.B1(n_13),
.B2(n_104),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_188),
.A2(n_153),
.B1(n_171),
.B2(n_180),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_94),
.B(n_12),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_108),
.B(n_112),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_108),
.C(n_93),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_116),
.A2(n_134),
.B1(n_96),
.B2(n_106),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_192),
.A2(n_110),
.B1(n_96),
.B2(n_106),
.Y(n_200)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_90),
.B(n_93),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_196),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_90),
.B(n_93),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_200),
.A2(n_218),
.B1(n_152),
.B2(n_157),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_153),
.A2(n_129),
.B1(n_110),
.B2(n_125),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_202),
.A2(n_225),
.B1(n_152),
.B2(n_184),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_215),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_144),
.B(n_129),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_SL g216 ( 
.A(n_177),
.B(n_138),
.C(n_105),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_SL g264 ( 
.A(n_216),
.B(n_186),
.C(n_211),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_160),
.A2(n_120),
.B(n_143),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_233),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_222),
.A2(n_230),
.B1(n_242),
.B2(n_154),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_148),
.B(n_149),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_241),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_164),
.A2(n_130),
.B1(n_143),
.B2(n_120),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_175),
.A2(n_166),
.B1(n_161),
.B2(n_147),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_161),
.B(n_189),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_159),
.Y(n_258)
);

AO21x2_ASAP7_75t_L g274 ( 
.A1(n_237),
.A2(n_200),
.B(n_206),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_173),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_147),
.A2(n_185),
.B1(n_169),
.B2(n_189),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_243),
.A2(n_245),
.B1(n_251),
.B2(n_265),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_244),
.B(n_272),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_191),
.B1(n_146),
.B2(n_151),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_158),
.C(n_181),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_255),
.C(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_199),
.A2(n_168),
.B1(n_167),
.B2(n_193),
.Y(n_251)
);

AOI22x1_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_173),
.B1(n_145),
.B2(n_170),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_253),
.A2(n_232),
.B(n_231),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_254),
.A2(n_267),
.B1(n_272),
.B2(n_281),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_170),
.C(n_173),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_198),
.Y(n_256)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_187),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_258),
.B(n_268),
.Y(n_295)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_198),
.Y(n_259)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_186),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_261),
.B(n_262),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_186),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_213),
.B(n_201),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_269),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_264),
.A2(n_255),
.B(n_253),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_199),
.A2(n_219),
.B1(n_214),
.B2(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_224),
.Y(n_266)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_219),
.A2(n_242),
.B1(n_218),
.B2(n_197),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_208),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_270),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_197),
.A2(n_233),
.B1(n_234),
.B2(n_225),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_274),
.B1(n_240),
.B2(n_210),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_217),
.A2(n_222),
.B1(n_237),
.B2(n_234),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_227),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_273),
.A2(n_276),
.B1(n_279),
.B2(n_231),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_205),
.B(n_241),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_275),
.Y(n_293)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_237),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_210),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_235),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_216),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_267),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_237),
.A2(n_212),
.B1(n_207),
.B2(n_206),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_212),
.A2(n_235),
.B1(n_240),
.B2(n_220),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_276),
.B1(n_274),
.B2(n_279),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_287),
.A2(n_292),
.B1(n_296),
.B2(n_302),
.Y(n_321)
);

AO22x1_ASAP7_75t_L g288 ( 
.A1(n_246),
.A2(n_239),
.B1(n_232),
.B2(n_238),
.Y(n_288)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_288),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_277),
.A2(n_235),
.B1(n_220),
.B2(n_239),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_265),
.A2(n_209),
.B1(n_204),
.B2(n_238),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_305),
.B(n_282),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_298),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_246),
.A2(n_204),
.B(n_209),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_307),
.B(n_289),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_301),
.Y(n_333)
);

OAI32xp33_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_254),
.A3(n_245),
.B1(n_258),
.B2(n_248),
.Y(n_301)
);

XOR2x2_ASAP7_75t_SL g341 ( 
.A(n_301),
.B(n_295),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_244),
.B(n_251),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_303),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_264),
.A2(n_253),
.B(n_271),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_249),
.C(n_252),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_286),
.C(n_295),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_259),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_310),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_260),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_274),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_303),
.Y(n_330)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_274),
.A2(n_277),
.B1(n_265),
.B2(n_230),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_315),
.A2(n_302),
.B1(n_287),
.B2(n_303),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_274),
.A2(n_254),
.B1(n_272),
.B2(n_281),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_316),
.A2(n_290),
.B1(n_300),
.B2(n_313),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_318),
.A2(n_319),
.B(n_320),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_307),
.B(n_297),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_311),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_322),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_312),
.B(n_293),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_324),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_310),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_332),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_328),
.A2(n_329),
.B1(n_343),
.B2(n_326),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_290),
.B1(n_289),
.B2(n_302),
.Y(n_329)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_330),
.Y(n_350)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_331),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_296),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_334),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_292),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_335),
.A2(n_336),
.B1(n_288),
.B2(n_314),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_309),
.A2(n_293),
.B1(n_299),
.B2(n_308),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_338),
.Y(n_360)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_338),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_288),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_344),
.C(n_284),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_286),
.A2(n_285),
.B1(n_306),
.B2(n_291),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_285),
.B(n_283),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_291),
.B(n_283),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_329),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_351),
.A2(n_356),
.B1(n_361),
.B2(n_368),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_353),
.C(n_355),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_284),
.C(n_294),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_344),
.Y(n_354)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_354),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_294),
.C(n_317),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_322),
.A2(n_317),
.B1(n_335),
.B2(n_325),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_327),
.C(n_336),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_365),
.C(n_323),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_322),
.A2(n_326),
.B1(n_321),
.B2(n_332),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_330),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_363),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_327),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_364),
.A2(n_321),
.B1(n_337),
.B2(n_334),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_320),
.C(n_319),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_333),
.A2(n_318),
.B1(n_323),
.B2(n_337),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_380),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_367),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_378),
.Y(n_386)
);

XNOR2x1_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_358),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_346),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_375),
.A2(n_351),
.B1(n_368),
.B2(n_361),
.Y(n_390)
);

XOR2x2_ASAP7_75t_SL g394 ( 
.A(n_376),
.B(n_348),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_367),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_328),
.B1(n_340),
.B2(n_345),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_379),
.A2(n_348),
.B1(n_346),
.B2(n_349),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_331),
.C(n_339),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_340),
.C(n_355),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_383),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_366),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_382),
.B(n_385),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_347),
.C(n_350),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_359),
.Y(n_384)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_384),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_362),
.C(n_363),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_384),
.A2(n_357),
.B1(n_360),
.B2(n_349),
.Y(n_389)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_389),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_390),
.A2(n_379),
.B1(n_373),
.B2(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_377),
.Y(n_391)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_393),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_376),
.C(n_373),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_383),
.Y(n_408)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_385),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_397),
.B(n_380),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_372),
.A2(n_360),
.B(n_378),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_398),
.A2(n_386),
.B(n_393),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_399),
.A2(n_396),
.B1(n_386),
.B2(n_369),
.Y(n_413)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_400),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_395),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_387),
.B(n_370),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_388),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_370),
.C(n_381),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_392),
.Y(n_414)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_407),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_408),
.B(n_402),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_411),
.B(n_414),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_405),
.B(n_392),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_413),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_415),
.B(n_408),
.C(n_399),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_416),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_418),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_409),
.A2(n_410),
.B(n_398),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_419),
.B(n_406),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_423),
.Y(n_425)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_420),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_424),
.B(n_421),
.C(n_412),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_426),
.A2(n_422),
.B(n_417),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_427),
.A2(n_424),
.B(n_415),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_428),
.A2(n_425),
.B(n_401),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_403),
.B(n_407),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_430),
.A2(n_411),
.B(n_401),
.Y(n_431)
);


endmodule