module fake_jpeg_4260_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_20),
.B(n_24),
.Y(n_56)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_26),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_39),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_26),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_22),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_24),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_48),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_SL g54 ( 
.A(n_33),
.B(n_22),
.C(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_31),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_37),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_20),
.B1(n_24),
.B2(n_28),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_20),
.B1(n_34),
.B2(n_38),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_20),
.B1(n_15),
.B2(n_28),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_62),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_65),
.Y(n_87)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_76),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_72),
.Y(n_96)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_15),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_29),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_69),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_50),
.B1(n_43),
.B2(n_49),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_45),
.B1(n_60),
.B2(n_66),
.Y(n_116)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_86),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_46),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_93),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_72),
.Y(n_98)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_42),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_0),
.B(n_1),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_70),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_78),
.C(n_58),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_105),
.C(n_108),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_55),
.C(n_63),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_73),
.B(n_43),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_99),
.B(n_80),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_44),
.B1(n_36),
.B2(n_54),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_114),
.B1(n_112),
.B2(n_104),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_63),
.C(n_36),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_115),
.B(n_91),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_23),
.B(n_60),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_83),
.B1(n_44),
.B2(n_96),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_99),
.Y(n_130)
);

NOR4xp25_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_89),
.C(n_100),
.D(n_87),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_121),
.B(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_133),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_115),
.A2(n_100),
.B(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_87),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_129),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_137),
.B1(n_113),
.B2(n_111),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_85),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_119),
.B(n_105),
.C(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_136),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_135),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_101),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_128),
.B(n_124),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_147),
.B(n_135),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_112),
.C(n_108),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_151),
.C(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_144),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_134),
.B1(n_132),
.B2(n_137),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_153),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_109),
.C(n_83),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_109),
.A3(n_88),
.B1(n_31),
.B2(n_45),
.C1(n_19),
.C2(n_18),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_23),
.Y(n_164)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_157),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_160),
.C(n_162),
.Y(n_171)
);

XOR2x2_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_130),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_133),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_140),
.B1(n_147),
.B2(n_138),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_127),
.C(n_103),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_101),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_166),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_127),
.C(n_70),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_21),
.B1(n_18),
.B2(n_19),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_21),
.B1(n_17),
.B2(n_12),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_147),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_29),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_143),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_1),
.Y(n_183)
);

INVxp33_ASAP7_75t_SL g169 ( 
.A(n_165),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g184 ( 
.A(n_169),
.B(n_1),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_147),
.C(n_153),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_160),
.C(n_162),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g176 ( 
.A(n_166),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_180),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_29),
.C(n_11),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_29),
.C(n_11),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_8),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_184),
.B(n_3),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_185),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_189),
.Y(n_195)
);

AOI21x1_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_177),
.B(n_168),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_188),
.A2(n_190),
.B1(n_13),
.B2(n_14),
.Y(n_194)
);

OAI321xp33_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_167),
.A3(n_177),
.B1(n_13),
.B2(n_10),
.C(n_12),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_191),
.B(n_193),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_178),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_197),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_187),
.B(n_14),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_8),
.B1(n_9),
.B2(n_35),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_9),
.B1(n_40),
.B2(n_35),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_SL g202 ( 
.A(n_196),
.B(n_9),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_35),
.B(n_40),
.C(n_199),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_203),
.A2(n_204),
.B(n_201),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_202),
.Y(n_206)
);


endmodule