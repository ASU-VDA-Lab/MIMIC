module fake_jpeg_15499_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx6_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_7),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_17),
.B1(n_5),
.B2(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

OA22x2_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

MAJx2_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_13),
.C(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_23),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_17),
.B1(n_10),
.B2(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_8),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_27),
.C(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_15),
.B1(n_19),
.B2(n_27),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_20),
.C(n_21),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_31),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_18),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_25),
.B(n_28),
.Y(n_34)
);

BUFx24_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_10),
.Y(n_36)
);

NOR2x1_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_33),
.Y(n_39)
);

AOI322xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_12),
.A3(n_16),
.B1(n_9),
.B2(n_5),
.C1(n_0),
.C2(n_18),
.Y(n_40)
);

NOR3xp33_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_12),
.C(n_38),
.Y(n_41)
);

NAND4xp25_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_0),
.C(n_39),
.D(n_40),
.Y(n_42)
);


endmodule