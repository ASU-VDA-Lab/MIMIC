module real_aes_8371_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g185 ( .A1(n_0), .A2(n_186), .B(n_189), .C(n_193), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_1), .B(n_177), .Y(n_196) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g460 ( .A(n_2), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_3), .B(n_187), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_4), .A2(n_150), .B(n_153), .C(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_5), .A2(n_145), .B(n_567), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_6), .A2(n_145), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_7), .B(n_177), .Y(n_573) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_8), .A2(n_179), .B(n_251), .Y(n_250) );
AND2x6_ASAP7_75t_L g150 ( .A(n_9), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_10), .A2(n_150), .B(n_153), .C(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g534 ( .A(n_11), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_12), .B(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_12), .B(n_39), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_13), .B(n_192), .Y(n_545) );
INVx1_ASAP7_75t_L g171 ( .A(n_14), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_15), .B(n_187), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_16), .A2(n_188), .B(n_553), .C(n_555), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_17), .B(n_177), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_18), .B(n_165), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_19), .A2(n_153), .B(n_156), .C(n_164), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_20), .A2(n_191), .B(n_259), .C(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_21), .B(n_192), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_22), .B(n_192), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_23), .Y(n_515) );
INVx1_ASAP7_75t_L g495 ( .A(n_24), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_25), .A2(n_153), .B(n_164), .C(n_254), .Y(n_253) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_26), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_27), .Y(n_541) );
INVx1_ASAP7_75t_L g509 ( .A(n_28), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_29), .A2(n_145), .B(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g148 ( .A(n_30), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_31), .A2(n_203), .B(n_204), .C(n_208), .Y(n_202) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_32), .A2(n_33), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_32), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_33), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_34), .A2(n_191), .B(n_570), .C(n_572), .Y(n_569) );
INVxp67_ASAP7_75t_L g510 ( .A(n_35), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_36), .B(n_256), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_37), .A2(n_153), .B(n_164), .C(n_494), .Y(n_493) );
CKINVDCx14_ASAP7_75t_R g568 ( .A(n_38), .Y(n_568) );
INVx1_ASAP7_75t_L g108 ( .A(n_39), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_40), .A2(n_193), .B(n_532), .C(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_41), .B(n_144), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_42), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_43), .B(n_187), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_44), .B(n_145), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_45), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_46), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_47), .A2(n_203), .B(n_208), .C(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g190 ( .A(n_48), .Y(n_190) );
INVx1_ASAP7_75t_L g234 ( .A(n_49), .Y(n_234) );
INVx1_ASAP7_75t_L g581 ( .A(n_50), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_51), .B(n_145), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_52), .Y(n_173) );
CKINVDCx14_ASAP7_75t_R g530 ( .A(n_53), .Y(n_530) );
AOI22xp5_ASAP7_75t_SL g467 ( .A1(n_54), .A2(n_458), .B1(n_468), .B2(n_764), .Y(n_467) );
INVx1_ASAP7_75t_L g151 ( .A(n_55), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_56), .B(n_145), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_57), .B(n_177), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_58), .A2(n_163), .B(n_219), .C(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g170 ( .A(n_59), .Y(n_170) );
INVx1_ASAP7_75t_SL g571 ( .A(n_60), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_61), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_62), .B(n_187), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_63), .A2(n_105), .B1(n_114), .B2(n_769), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_64), .B(n_177), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_65), .B(n_188), .Y(n_269) );
INVx1_ASAP7_75t_L g518 ( .A(n_66), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_67), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_68), .B(n_158), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_69), .A2(n_153), .B(n_208), .C(n_217), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_70), .Y(n_243) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_72), .A2(n_145), .B(n_529), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_73), .A2(n_95), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_73), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_74), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_75), .A2(n_103), .B1(n_477), .B2(n_478), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_75), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_76), .A2(n_145), .B(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_77), .A2(n_144), .B(n_505), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_78), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_79), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_79), .Y(n_474) );
INVx1_ASAP7_75t_L g551 ( .A(n_80), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_81), .B(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_82), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_83), .A2(n_145), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g554 ( .A(n_84), .Y(n_554) );
INVx2_ASAP7_75t_L g168 ( .A(n_85), .Y(n_168) );
INVx1_ASAP7_75t_L g544 ( .A(n_86), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_87), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_88), .B(n_192), .Y(n_270) );
INVx2_ASAP7_75t_L g110 ( .A(n_89), .Y(n_110) );
OR2x2_ASAP7_75t_L g457 ( .A(n_89), .B(n_458), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_90), .A2(n_153), .B(n_208), .C(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_91), .B(n_145), .Y(n_201) );
INVx1_ASAP7_75t_L g205 ( .A(n_92), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_93), .B(n_463), .Y(n_462) );
INVxp67_ASAP7_75t_L g246 ( .A(n_94), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_95), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_96), .A2(n_473), .B1(n_479), .B2(n_480), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_96), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_97), .B(n_179), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_98), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g218 ( .A(n_99), .Y(n_218) );
INVx1_ASAP7_75t_L g265 ( .A(n_100), .Y(n_265) );
INVx2_ASAP7_75t_L g584 ( .A(n_101), .Y(n_584) );
AND2x2_ASAP7_75t_L g236 ( .A(n_102), .B(n_167), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_103), .Y(n_477) );
INVx1_ASAP7_75t_L g769 ( .A(n_105), .Y(n_769) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx2_ASAP7_75t_L g469 ( .A(n_110), .Y(n_469) );
INVx1_ASAP7_75t_L g482 ( .A(n_110), .Y(n_482) );
NOR2x2_ASAP7_75t_L g766 ( .A(n_110), .B(n_458), .Y(n_766) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_466), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g768 ( .A(n_119), .Y(n_768) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_455), .B(n_462), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_126), .B2(n_127), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_124), .B(n_178), .Y(n_546) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B1(n_132), .B2(n_133), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_132), .A2(n_133), .B1(n_471), .B2(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_410), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_345), .Y(n_134) );
NAND4xp25_ASAP7_75t_SL g135 ( .A(n_136), .B(n_290), .C(n_314), .D(n_337), .Y(n_135) );
AOI221xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_227), .B1(n_261), .B2(n_274), .C(n_277), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_197), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_139), .A2(n_175), .B1(n_228), .B2(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_139), .B(n_198), .Y(n_348) );
AND2x2_ASAP7_75t_L g367 ( .A(n_139), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_139), .B(n_351), .Y(n_437) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_175), .Y(n_139) );
AND2x2_ASAP7_75t_L g305 ( .A(n_140), .B(n_198), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_140), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g328 ( .A(n_140), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g333 ( .A(n_140), .B(n_176), .Y(n_333) );
INVx2_ASAP7_75t_L g365 ( .A(n_140), .Y(n_365) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_140), .Y(n_409) );
AND2x2_ASAP7_75t_L g426 ( .A(n_140), .B(n_303), .Y(n_426) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g344 ( .A(n_141), .B(n_303), .Y(n_344) );
AND2x4_ASAP7_75t_L g358 ( .A(n_141), .B(n_175), .Y(n_358) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_141), .Y(n_362) );
AND2x2_ASAP7_75t_L g382 ( .A(n_141), .B(n_297), .Y(n_382) );
AND2x2_ASAP7_75t_L g432 ( .A(n_141), .B(n_199), .Y(n_432) );
AND2x2_ASAP7_75t_L g442 ( .A(n_141), .B(n_176), .Y(n_442) );
OR2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_172), .Y(n_141) );
AOI21xp5_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_152), .B(n_165), .Y(n_142) );
BUFx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_146), .B(n_150), .Y(n_266) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx1_ASAP7_75t_L g260 ( .A(n_148), .Y(n_260) );
INVx1_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
INVx3_ASAP7_75t_L g188 ( .A(n_149), .Y(n_188) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_149), .Y(n_192) );
INVx1_ASAP7_75t_L g256 ( .A(n_149), .Y(n_256) );
BUFx3_ASAP7_75t_L g164 ( .A(n_150), .Y(n_164) );
INVx4_ASAP7_75t_SL g195 ( .A(n_150), .Y(n_195) );
INVx5_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx3_ASAP7_75t_L g194 ( .A(n_154), .Y(n_194) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_154), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_160), .B(n_162), .Y(n_156) );
INVx2_ASAP7_75t_L g161 ( .A(n_158), .Y(n_161) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g220 ( .A(n_159), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_161), .A2(n_205), .B(n_206), .C(n_207), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_161), .A2(n_207), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_161), .A2(n_518), .B(n_519), .C(n_520), .Y(n_517) );
O2A1O1Ixp5_ASAP7_75t_L g543 ( .A1(n_161), .A2(n_520), .B(n_544), .C(n_545), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_162), .A2(n_187), .B(n_495), .C(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_163), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_166), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g174 ( .A(n_167), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_167), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_167), .A2(n_231), .B(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_167), .A2(n_266), .B(n_492), .C(n_493), .Y(n_491) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_167), .A2(n_528), .B(n_535), .Y(n_527) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_168), .B(n_169), .Y(n_167) );
AND2x2_ASAP7_75t_L g180 ( .A(n_168), .B(n_169), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_174), .A2(n_540), .B(n_546), .Y(n_539) );
AND2x2_ASAP7_75t_L g298 ( .A(n_175), .B(n_198), .Y(n_298) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_175), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_175), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g388 ( .A(n_175), .Y(n_388) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g276 ( .A(n_176), .B(n_213), .Y(n_276) );
AND2x2_ASAP7_75t_L g303 ( .A(n_176), .B(n_214), .Y(n_303) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_181), .B(n_196), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_178), .B(n_210), .Y(n_209) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_178), .A2(n_215), .B(n_225), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_178), .B(n_226), .Y(n_225) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_178), .A2(n_264), .B(n_271), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_178), .B(n_498), .Y(n_497) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_178), .A2(n_514), .B(n_521), .Y(n_513) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_179), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_179), .A2(n_252), .B(n_253), .Y(n_251) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g273 ( .A(n_180), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_SL g182 ( .A1(n_183), .A2(n_184), .B(n_185), .C(n_195), .Y(n_182) );
INVx2_ASAP7_75t_L g203 ( .A(n_184), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_184), .A2(n_195), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_184), .A2(n_195), .B(n_506), .C(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_184), .A2(n_195), .B(n_530), .C(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_SL g550 ( .A1(n_184), .A2(n_195), .B(n_551), .C(n_552), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g567 ( .A1(n_184), .A2(n_195), .B(n_568), .C(n_569), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_SL g580 ( .A1(n_184), .A2(n_195), .B(n_581), .C(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_187), .B(n_246), .Y(n_245) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_187), .A2(n_220), .B1(n_509), .B2(n_510), .Y(n_508) );
INVx5_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_188), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_191), .B(n_571), .Y(n_570) );
INVx4_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g532 ( .A(n_192), .Y(n_532) );
INVx2_ASAP7_75t_L g520 ( .A(n_193), .Y(n_520) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_194), .Y(n_207) );
INVx1_ASAP7_75t_L g555 ( .A(n_194), .Y(n_555) );
INVx1_ASAP7_75t_L g208 ( .A(n_195), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_197), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_211), .Y(n_197) );
OR2x2_ASAP7_75t_L g329 ( .A(n_198), .B(n_212), .Y(n_329) );
AND2x2_ASAP7_75t_L g366 ( .A(n_198), .B(n_276), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_198), .B(n_297), .Y(n_377) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_198), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_198), .B(n_333), .Y(n_450) );
INVx5_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
BUFx2_ASAP7_75t_L g275 ( .A(n_199), .Y(n_275) );
AND2x2_ASAP7_75t_L g284 ( .A(n_199), .B(n_212), .Y(n_284) );
AND2x2_ASAP7_75t_L g400 ( .A(n_199), .B(n_295), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_199), .B(n_333), .Y(n_422) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_209), .Y(n_199) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_212), .Y(n_368) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_213), .Y(n_320) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
BUFx2_ASAP7_75t_L g297 ( .A(n_214), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_224), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_221), .C(n_222), .Y(n_217) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_220), .B(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_220), .B(n_584), .Y(n_583) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx3_ASAP7_75t_L g572 ( .A(n_223), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_237), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_228), .B(n_310), .Y(n_429) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_229), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g281 ( .A(n_229), .B(n_282), .Y(n_281) );
INVx5_ASAP7_75t_SL g289 ( .A(n_229), .Y(n_289) );
OR2x2_ASAP7_75t_L g312 ( .A(n_229), .B(n_282), .Y(n_312) );
OR2x2_ASAP7_75t_L g322 ( .A(n_229), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g385 ( .A(n_229), .B(n_239), .Y(n_385) );
AND2x2_ASAP7_75t_SL g423 ( .A(n_229), .B(n_238), .Y(n_423) );
NOR4xp25_ASAP7_75t_L g444 ( .A(n_229), .B(n_365), .C(n_445), .D(n_446), .Y(n_444) );
AND2x2_ASAP7_75t_L g454 ( .A(n_229), .B(n_286), .Y(n_454) );
OR2x6_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g279 ( .A(n_238), .B(n_275), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_238), .B(n_281), .Y(n_448) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_248), .Y(n_238) );
OR2x2_ASAP7_75t_L g288 ( .A(n_239), .B(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g295 ( .A(n_239), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_239), .B(n_263), .Y(n_307) );
INVxp67_ASAP7_75t_L g310 ( .A(n_239), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_239), .B(n_282), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_239), .B(n_249), .Y(n_376) );
AND2x2_ASAP7_75t_L g391 ( .A(n_239), .B(n_286), .Y(n_391) );
OR2x2_ASAP7_75t_L g420 ( .A(n_239), .B(n_249), .Y(n_420) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_247), .Y(n_239) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_240), .A2(n_549), .B(n_556), .Y(n_548) );
OA21x2_ASAP7_75t_L g565 ( .A1(n_240), .A2(n_566), .B(n_573), .Y(n_565) );
OA21x2_ASAP7_75t_L g578 ( .A1(n_240), .A2(n_579), .B(n_585), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_248), .B(n_325), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_248), .B(n_289), .Y(n_428) );
OR2x2_ASAP7_75t_L g449 ( .A(n_248), .B(n_326), .Y(n_449) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g262 ( .A(n_249), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g286 ( .A(n_249), .B(n_282), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_249), .B(n_263), .Y(n_301) );
AND2x2_ASAP7_75t_L g371 ( .A(n_249), .B(n_295), .Y(n_371) );
AND2x2_ASAP7_75t_L g405 ( .A(n_249), .B(n_289), .Y(n_405) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_250), .B(n_289), .Y(n_308) );
AND2x2_ASAP7_75t_L g336 ( .A(n_250), .B(n_263), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_257), .B(n_258), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_258), .A2(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_261), .B(n_344), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_262), .A2(n_351), .B1(n_387), .B2(n_404), .C(n_406), .Y(n_403) );
INVx5_ASAP7_75t_SL g282 ( .A(n_263), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_266), .B(n_267), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_266), .A2(n_515), .B(n_516), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_266), .A2(n_541), .B(n_542), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g503 ( .A(n_273), .Y(n_503) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
OAI33xp33_ASAP7_75t_L g302 ( .A1(n_275), .A2(n_303), .A3(n_304), .B1(n_306), .B2(n_309), .B3(n_313), .Y(n_302) );
OR2x2_ASAP7_75t_L g318 ( .A(n_275), .B(n_319), .Y(n_318) );
AOI322xp5_ASAP7_75t_L g427 ( .A1(n_275), .A2(n_344), .A3(n_351), .B1(n_428), .B2(n_429), .C1(n_430), .C2(n_433), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_275), .B(n_303), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_SL g451 ( .A1(n_275), .A2(n_303), .B(n_452), .C(n_454), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_276), .A2(n_291), .B1(n_296), .B2(n_299), .C(n_302), .Y(n_290) );
INVx1_ASAP7_75t_L g383 ( .A(n_276), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_276), .B(n_432), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_280), .B1(n_283), .B2(n_285), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g360 ( .A(n_281), .B(n_295), .Y(n_360) );
AND2x2_ASAP7_75t_L g418 ( .A(n_281), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g326 ( .A(n_282), .B(n_289), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_282), .B(n_295), .Y(n_354) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_284), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_284), .B(n_362), .Y(n_416) );
OAI321xp33_ASAP7_75t_L g435 ( .A1(n_284), .A2(n_357), .A3(n_436), .B1(n_437), .B2(n_438), .C(n_439), .Y(n_435) );
INVx1_ASAP7_75t_L g402 ( .A(n_285), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_286), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g341 ( .A(n_286), .B(n_289), .Y(n_341) );
AOI321xp33_ASAP7_75t_L g399 ( .A1(n_286), .A2(n_303), .A3(n_400), .B1(n_401), .B2(n_402), .C(n_403), .Y(n_399) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_301), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_289), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_289), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_289), .B(n_375), .Y(n_412) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g335 ( .A(n_293), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g300 ( .A(n_294), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g408 ( .A(n_295), .Y(n_408) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_298), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_305), .B(n_340), .Y(n_389) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
OR2x2_ASAP7_75t_L g353 ( .A(n_308), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g398 ( .A(n_308), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_309), .A2(n_356), .B1(n_359), .B2(n_361), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g453 ( .A(n_312), .B(n_376), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B1(n_321), .B2(n_327), .C(n_330), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_L g351 ( .A(n_320), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_SL g397 ( .A(n_323), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_325), .B(n_375), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_325), .A2(n_393), .B(n_395), .Y(n_392) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g438 ( .A(n_326), .B(n_420), .Y(n_438) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_SL g340 ( .A(n_329), .Y(n_340) );
AOI21xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B(n_334), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g384 ( .A(n_336), .B(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g446 ( .A(n_336), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_341), .B(n_342), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_340), .B(n_358), .Y(n_394) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g415 ( .A(n_344), .Y(n_415) );
NAND5xp2_ASAP7_75t_L g345 ( .A(n_346), .B(n_363), .C(n_372), .D(n_392), .E(n_399), .Y(n_345) );
O2A1O1Ixp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B(n_352), .C(n_355), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g387 ( .A(n_351), .Y(n_387) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_359), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g401 ( .A(n_361), .Y(n_401) );
OAI21xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_367), .B(n_369), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_364), .A2(n_418), .B1(n_421), .B2(n_423), .C(n_424), .Y(n_417) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AOI321xp33_ASAP7_75t_L g372 ( .A1(n_365), .A2(n_373), .A3(n_377), .B1(n_378), .B2(n_384), .C(n_386), .Y(n_372) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g443 ( .A(n_377), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_379), .B(n_383), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g395 ( .A(n_380), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
NOR2xp67_ASAP7_75t_SL g407 ( .A(n_381), .B(n_388), .Y(n_407) );
AOI321xp33_ASAP7_75t_SL g439 ( .A1(n_384), .A2(n_440), .A3(n_441), .B1(n_442), .B2(n_443), .C(n_444), .Y(n_439) );
O2A1O1Ixp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_389), .C(n_390), .Y(n_386) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_397), .B(n_405), .Y(n_434) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .C(n_409), .Y(n_406) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_435), .C(n_447), .Y(n_410) );
OAI211xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_413), .B(n_417), .C(n_427), .Y(n_411) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_415), .B(n_416), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_416), .A2(n_448), .B1(n_449), .B2(n_450), .C(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g436 ( .A(n_418), .Y(n_436) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g440 ( .A(n_438), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
CKINVDCx14_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g465 ( .A(n_457), .Y(n_465) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_462), .A2(n_467), .B(n_767), .Y(n_466) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B1(n_481), .B2(n_483), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_471), .A2(n_472), .B1(n_484), .B2(n_485), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g480 ( .A(n_473), .Y(n_480) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR4x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_654), .C(n_701), .D(n_741), .Y(n_485) );
NAND3xp33_ASAP7_75t_SL g486 ( .A(n_487), .B(n_600), .C(n_629), .Y(n_486) );
AOI211xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_523), .B(n_557), .C(n_593), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_488), .A2(n_613), .B(n_630), .C(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_490), .B(n_592), .Y(n_591) );
INVx3_ASAP7_75t_SL g596 ( .A(n_490), .Y(n_596) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_490), .Y(n_608) );
AND2x4_ASAP7_75t_L g612 ( .A(n_490), .B(n_564), .Y(n_612) );
AND2x2_ASAP7_75t_L g623 ( .A(n_490), .B(n_513), .Y(n_623) );
OR2x2_ASAP7_75t_L g647 ( .A(n_490), .B(n_560), .Y(n_647) );
AND2x2_ASAP7_75t_L g660 ( .A(n_490), .B(n_565), .Y(n_660) );
AND2x2_ASAP7_75t_L g700 ( .A(n_490), .B(n_686), .Y(n_700) );
AND2x2_ASAP7_75t_L g707 ( .A(n_490), .B(n_670), .Y(n_707) );
AND2x2_ASAP7_75t_L g737 ( .A(n_490), .B(n_500), .Y(n_737) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_497), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_499), .B(n_664), .Y(n_676) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_512), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_500), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g614 ( .A(n_500), .B(n_512), .Y(n_614) );
BUFx3_ASAP7_75t_L g622 ( .A(n_500), .Y(n_622) );
OR2x2_ASAP7_75t_L g643 ( .A(n_500), .B(n_526), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_500), .B(n_664), .Y(n_754) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_504), .B(n_511), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_502), .A2(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g561 ( .A(n_504), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_511), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_512), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g607 ( .A(n_512), .Y(n_607) );
AND2x2_ASAP7_75t_L g670 ( .A(n_512), .B(n_565), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_512), .A2(n_673), .B1(n_675), .B2(n_677), .C(n_678), .Y(n_672) );
AND2x2_ASAP7_75t_L g686 ( .A(n_512), .B(n_560), .Y(n_686) );
AND2x2_ASAP7_75t_L g712 ( .A(n_512), .B(n_596), .Y(n_712) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g592 ( .A(n_513), .B(n_565), .Y(n_592) );
BUFx2_ASAP7_75t_L g726 ( .A(n_513), .Y(n_726) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI32xp33_ASAP7_75t_L g692 ( .A1(n_524), .A2(n_653), .A3(n_667), .B1(n_693), .B2(n_694), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_536), .Y(n_524) );
AND2x2_ASAP7_75t_L g633 ( .A(n_525), .B(n_577), .Y(n_633) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g615 ( .A(n_526), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_526), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g687 ( .A(n_526), .B(n_577), .Y(n_687) );
AND2x2_ASAP7_75t_L g698 ( .A(n_526), .B(n_590), .Y(n_698) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g599 ( .A(n_527), .B(n_578), .Y(n_599) );
AND2x2_ASAP7_75t_L g603 ( .A(n_527), .B(n_578), .Y(n_603) );
AND2x2_ASAP7_75t_L g638 ( .A(n_527), .B(n_589), .Y(n_638) );
AND2x2_ASAP7_75t_L g645 ( .A(n_527), .B(n_547), .Y(n_645) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_527), .A2(n_596), .B(n_607), .C(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g704 ( .A(n_527), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_527), .B(n_538), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_536), .B(n_587), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_536), .B(n_603), .Y(n_693) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g598 ( .A(n_537), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
AND2x2_ASAP7_75t_L g590 ( .A(n_538), .B(n_548), .Y(n_590) );
OR2x2_ASAP7_75t_L g605 ( .A(n_538), .B(n_548), .Y(n_605) );
AND2x2_ASAP7_75t_L g628 ( .A(n_538), .B(n_589), .Y(n_628) );
INVx1_ASAP7_75t_L g632 ( .A(n_538), .Y(n_632) );
AND2x2_ASAP7_75t_L g651 ( .A(n_538), .B(n_588), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g661 ( .A1(n_538), .A2(n_616), .B1(n_662), .B2(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_538), .B(n_704), .Y(n_728) );
AND2x2_ASAP7_75t_L g743 ( .A(n_538), .B(n_603), .Y(n_743) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g575 ( .A(n_539), .Y(n_575) );
AND2x2_ASAP7_75t_L g617 ( .A(n_539), .B(n_548), .Y(n_617) );
AND2x2_ASAP7_75t_L g619 ( .A(n_539), .B(n_577), .Y(n_619) );
AND3x2_ASAP7_75t_L g681 ( .A(n_539), .B(n_645), .C(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g716 ( .A(n_547), .B(n_588), .Y(n_716) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g577 ( .A(n_548), .B(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_548), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_548), .B(n_587), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_548), .B(n_628), .C(n_704), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_574), .B1(n_586), .B2(n_591), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_560), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g668 ( .A(n_560), .Y(n_668) );
OAI31xp33_ASAP7_75t_L g684 ( .A1(n_563), .A2(n_685), .A3(n_686), .B(n_687), .Y(n_684) );
AND2x2_ASAP7_75t_L g709 ( .A(n_563), .B(n_596), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_563), .B(n_622), .Y(n_755) );
AND2x2_ASAP7_75t_L g664 ( .A(n_564), .B(n_596), .Y(n_664) );
AND2x2_ASAP7_75t_L g725 ( .A(n_564), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g595 ( .A(n_565), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g653 ( .A(n_565), .Y(n_653) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
CKINVDCx16_ASAP7_75t_R g674 ( .A(n_575), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_576), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AOI221x1_ASAP7_75t_SL g641 ( .A1(n_577), .A2(n_642), .B1(n_644), .B2(n_646), .C(n_648), .Y(n_641) );
INVx2_ASAP7_75t_L g589 ( .A(n_578), .Y(n_589) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_578), .Y(n_683) );
INVx1_ASAP7_75t_L g671 ( .A(n_586), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_587), .B(n_604), .Y(n_696) );
INVx1_ASAP7_75t_SL g759 ( .A(n_587), .Y(n_759) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g677 ( .A(n_590), .B(n_603), .Y(n_677) );
INVx1_ASAP7_75t_L g745 ( .A(n_591), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_591), .B(n_674), .Y(n_758) );
INVx2_ASAP7_75t_SL g597 ( .A(n_592), .Y(n_597) );
AND2x2_ASAP7_75t_L g640 ( .A(n_592), .B(n_596), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_592), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_592), .B(n_667), .Y(n_694) );
AOI21xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_597), .B(n_598), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_595), .B(n_667), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_595), .B(n_622), .Y(n_763) );
OR2x2_ASAP7_75t_L g635 ( .A(n_596), .B(n_614), .Y(n_635) );
AND2x2_ASAP7_75t_L g734 ( .A(n_596), .B(n_725), .Y(n_734) );
OAI22xp5_ASAP7_75t_SL g609 ( .A1(n_597), .A2(n_610), .B1(n_615), .B2(n_618), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_597), .B(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g657 ( .A(n_599), .B(n_605), .Y(n_657) );
INVx1_ASAP7_75t_L g721 ( .A(n_599), .Y(n_721) );
AOI311xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_606), .A3(n_608), .B(n_609), .C(n_620), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_604), .A2(n_736), .B1(n_748), .B2(n_751), .C(n_753), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_604), .B(n_759), .Y(n_761) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g658 ( .A(n_606), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g648 ( .A1(n_607), .A2(n_649), .B(n_650), .C(n_652), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_SL g717 ( .A1(n_611), .A2(n_613), .B(n_718), .C(n_719), .Y(n_717) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_612), .B(n_686), .Y(n_752) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_615), .A2(n_635), .B1(n_636), .B2(n_639), .C(n_641), .Y(n_634) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g637 ( .A(n_617), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g720 ( .A(n_617), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_621), .A2(n_679), .B(n_680), .C(n_684), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_622), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_622), .B(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVxp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g644 ( .A(n_628), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_632), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g746 ( .A(n_635), .Y(n_746) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_638), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g673 ( .A(n_638), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g750 ( .A(n_638), .Y(n_750) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g691 ( .A(n_640), .B(n_667), .Y(n_691) );
INVx1_ASAP7_75t_SL g685 ( .A(n_647), .Y(n_685) );
INVx1_ASAP7_75t_L g662 ( .A(n_653), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_672), .C(n_688), .Y(n_654) );
AOI322xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .A3(n_659), .B1(n_661), .B2(n_665), .C1(n_669), .C2(n_671), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g708 ( .A1(n_656), .A2(n_709), .B(n_710), .C(n_717), .Y(n_708) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_659), .A2(n_680), .B1(n_711), .B2(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g669 ( .A(n_667), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g706 ( .A(n_667), .B(n_707), .Y(n_706) );
AOI32xp33_ASAP7_75t_L g757 ( .A1(n_667), .A2(n_758), .A3(n_759), .B1(n_760), .B2(n_762), .Y(n_757) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g679 ( .A(n_670), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_670), .A2(n_723), .B1(n_727), .B2(n_729), .C(n_732), .Y(n_722) );
AND2x2_ASAP7_75t_L g736 ( .A(n_670), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g739 ( .A(n_674), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g749 ( .A(n_674), .B(n_750), .Y(n_749) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g740 ( .A(n_683), .B(n_704), .Y(n_740) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_692), .C(n_695), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI211xp5_ASAP7_75t_SL g701 ( .A1(n_702), .A2(n_705), .B(n_708), .C(n_722), .Y(n_701) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_716), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g731 ( .A(n_728), .Y(n_731) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_735), .B(n_738), .Y(n_732) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI211xp5_ASAP7_75t_SL g741 ( .A1(n_742), .A2(n_744), .B(n_747), .C(n_757), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AOI21xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx3_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
endmodule