module fake_jpeg_32052_n_129 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_44),
.Y(n_47)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_38),
.Y(n_59)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_52),
.B1(n_1),
.B2(n_5),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_19),
.B(n_4),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_25),
.B(n_23),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_22),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_21),
.B(n_29),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_21),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_28),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_75),
.B(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_77),
.Y(n_81)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_73),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_48),
.Y(n_70)
);

NAND2x1_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_29),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_72),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_6),
.B1(n_7),
.B2(n_11),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_13),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_7),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_55),
.C(n_49),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_11),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_84),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_90),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_SL g84 ( 
.A(n_78),
.B(n_59),
.C(n_53),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_55),
.B(n_60),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_76),
.B(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_60),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_91),
.Y(n_93)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_71),
.B(n_63),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_91),
.C(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_97),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_86),
.B(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_88),
.B1(n_82),
.B2(n_70),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_93),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_81),
.B1(n_72),
.B2(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_108),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_83),
.B1(n_84),
.B2(n_66),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_97),
.B(n_99),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_111),
.B(n_101),
.Y(n_118)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_114),
.C(n_66),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_104),
.A2(n_95),
.B(n_94),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_103),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_113),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_93),
.C(n_100),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_112),
.A2(n_107),
.B1(n_102),
.B2(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_105),
.B(n_101),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_118),
.B(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_122),
.Y(n_123)
);

AOI321xp33_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_53),
.A3(n_80),
.B1(n_56),
.B2(n_68),
.C(n_74),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_117),
.B1(n_58),
.B2(n_49),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_58),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_65),
.B(n_54),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_124),
.Y(n_129)
);


endmodule