module fake_jpeg_4554_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_44),
.Y(n_69)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_42),
.B(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_25),
.Y(n_67)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_53),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_50),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_52),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_56),
.Y(n_98)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_33),
.B1(n_37),
.B2(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_6),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_30),
.B(n_20),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_61),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_62),
.A2(n_70),
.B1(n_87),
.B2(n_88),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_63),
.A2(n_64),
.B(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_33),
.B1(n_35),
.B2(n_34),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_68),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_25),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_77),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_26),
.B1(n_22),
.B2(n_28),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_75),
.A2(n_78),
.B1(n_89),
.B2(n_95),
.Y(n_133)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_18),
.B1(n_16),
.B2(n_30),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_81),
.Y(n_116)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_92),
.Y(n_121)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_12),
.B(n_14),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_9),
.B(n_2),
.C(n_3),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_39),
.A2(n_18),
.B1(n_27),
.B2(n_24),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_41),
.A2(n_27),
.B1(n_24),
.B2(n_29),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_41),
.A2(n_36),
.B1(n_32),
.B2(n_29),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_36),
.B1(n_32),
.B2(n_0),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_97),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_40),
.A2(n_36),
.B1(n_32),
.B2(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_10),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_51),
.A2(n_36),
.B1(n_32),
.B2(n_1),
.Y(n_103)
);

CKINVDCx9p33_ASAP7_75t_R g128 ( 
.A(n_103),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_51),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_106),
.Y(n_127)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_38),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_4),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_111),
.B(n_114),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_67),
.B(n_1),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_138),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_72),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_118),
.B(n_119),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_126),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_61),
.B(n_2),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_125),
.A2(n_119),
.B1(n_113),
.B2(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_13),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g129 ( 
.A(n_71),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

CKINVDCx12_ASAP7_75t_R g134 ( 
.A(n_71),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_12),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_73),
.B(n_12),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_9),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_65),
.B(n_5),
.Y(n_138)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_141),
.Y(n_205)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_148),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_80),
.B1(n_81),
.B2(n_99),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_143),
.A2(n_129),
.B1(n_119),
.B2(n_140),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_91),
.B1(n_105),
.B2(n_102),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_147),
.A2(n_172),
.B1(n_129),
.B2(n_136),
.Y(n_190)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_149),
.B(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_114),
.Y(n_150)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_86),
.Y(n_151)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_79),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_164),
.Y(n_187)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_64),
.B1(n_95),
.B2(n_63),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_88),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_166),
.Y(n_200)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_171),
.B1(n_128),
.B2(n_123),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_65),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_169),
.B(n_175),
.Y(n_193)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_89),
.B1(n_90),
.B2(n_103),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_112),
.A2(n_125),
.B1(n_128),
.B2(n_117),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_116),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_173),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_84),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_9),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_10),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_115),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_142),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_192),
.B1(n_146),
.B2(n_145),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_195),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_185),
.A2(n_190),
.B1(n_211),
.B2(n_149),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_126),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_191),
.A2(n_204),
.B(n_212),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_135),
.B(n_132),
.C(n_140),
.Y(n_192)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_155),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_197),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_143),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_173),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_163),
.B(n_167),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_202),
.B(n_158),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_163),
.A2(n_116),
.B(n_127),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_210),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_134),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_158),
.A2(n_139),
.B1(n_109),
.B2(n_123),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_154),
.C(n_146),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_161),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_109),
.B1(n_124),
.B2(n_82),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_159),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_153),
.B(n_109),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_144),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_175),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_214),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_235),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_217),
.A2(n_239),
.B(n_207),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_220),
.B(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_224),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_152),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_152),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_229),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_209),
.B(n_158),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_192),
.B(n_204),
.Y(n_256)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_232),
.B(n_233),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_178),
.Y(n_233)
);

OAI22x1_ASAP7_75t_SL g234 ( 
.A1(n_177),
.A2(n_211),
.B1(n_201),
.B2(n_182),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_234),
.A2(n_241),
.B1(n_188),
.B2(n_205),
.Y(n_265)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_236),
.B(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_238),
.B(n_240),
.Y(n_267)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_145),
.Y(n_242)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_180),
.C(n_191),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_249),
.B(n_251),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_210),
.Y(n_250)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_236),
.B(n_181),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_177),
.B1(n_192),
.B2(n_184),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_255),
.B1(n_265),
.B2(n_242),
.Y(n_282)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_254),
.B(n_264),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_230),
.A2(n_192),
.B1(n_185),
.B2(n_202),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_239),
.Y(n_274)
);

AND2x4_ASAP7_75t_SL g257 ( 
.A(n_223),
.B(n_204),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_SL g261 ( 
.A1(n_218),
.A2(n_191),
.B(n_82),
.C(n_100),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_261),
.A2(n_226),
.B1(n_240),
.B2(n_233),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_189),
.Y(n_262)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_260),
.C(n_217),
.Y(n_272)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_280),
.B1(n_248),
.B2(n_245),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_274),
.B(n_282),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_257),
.C(n_263),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_275),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_227),
.C(n_238),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_244),
.Y(n_278)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_281),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_247),
.A2(n_225),
.B1(n_237),
.B2(n_224),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_246),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_283),
.B(n_285),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_228),
.B1(n_222),
.B2(n_235),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_284),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_244),
.B(n_216),
.Y(n_285)
);

OA21x2_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_256),
.B(n_253),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_294),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_170),
.Y(n_289)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_274),
.B(n_253),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_296),
.Y(n_301)
);

AOI321xp33_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_243),
.A3(n_252),
.B1(n_229),
.B2(n_248),
.C(n_249),
.Y(n_294)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_267),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_282),
.B(n_284),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_298),
.A2(n_275),
.B(n_278),
.Y(n_302)
);

BUFx4f_ASAP7_75t_SL g299 ( 
.A(n_283),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_270),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_270),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_302),
.A2(n_305),
.B(n_306),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_272),
.C(n_292),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_308),
.C(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_277),
.C(n_293),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_271),
.C(n_268),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_266),
.C(n_228),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_299),
.C(n_290),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_286),
.B1(n_298),
.B2(n_296),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_290),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_316),
.C(n_317),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_319),
.B(n_254),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_300),
.C(n_169),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_301),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_261),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_318),
.B(n_311),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_261),
.C(n_195),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_310),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_323),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_315),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_120),
.B(n_189),
.Y(n_329)
);

AO22x1_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_261),
.B1(n_215),
.B2(n_303),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_11),
.B1(n_166),
.B2(n_120),
.Y(n_331)
);

NOR2x1_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_313),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_331),
.B1(n_325),
.B2(n_11),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_332),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_333),
.C(n_100),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);


endmodule