module fake_jpeg_17030_n_282 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_17),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_31),
.B1(n_19),
.B2(n_17),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_30),
.B1(n_27),
.B2(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_49),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_51),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_21),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_53),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_26),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_59),
.B1(n_64),
.B2(n_46),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_19),
.B1(n_30),
.B2(n_26),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_31),
.B1(n_19),
.B2(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_30),
.B1(n_22),
.B2(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_32),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_30),
.B1(n_27),
.B2(n_23),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_SL g101 ( 
.A1(n_70),
.A2(n_83),
.B(n_90),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_84),
.B1(n_12),
.B2(n_2),
.Y(n_113)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_75),
.Y(n_102)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_78),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_95),
.B1(n_34),
.B2(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_81),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_33),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_47),
.B(n_62),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_43),
.B1(n_42),
.B2(n_25),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_37),
.B(n_42),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_53),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_93),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_34),
.B(n_29),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_96),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_34),
.B1(n_29),
.B2(n_3),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_34),
.B1(n_29),
.B2(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_63),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_99),
.B(n_119),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_113),
.B1(n_71),
.B2(n_72),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_64),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_107),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_24),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_48),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_53),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_125),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_64),
.B1(n_48),
.B2(n_24),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_120),
.A2(n_124),
.B1(n_95),
.B2(n_93),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_33),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_94),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_68),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_64),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_67),
.B(n_24),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_130),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_69),
.B1(n_81),
.B2(n_116),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_85),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_94),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_74),
.C(n_67),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_139),
.C(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_142),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_110),
.C(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_73),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_152),
.B1(n_115),
.B2(n_111),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_101),
.A2(n_105),
.B(n_123),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_115),
.B(n_108),
.Y(n_159)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_147),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_88),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_116),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_80),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_154),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_98),
.A2(n_72),
.B1(n_69),
.B2(n_97),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_93),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_164),
.C(n_168),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_124),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_128),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_100),
.B(n_120),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_167),
.B(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_161),
.B1(n_163),
.B2(n_166),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_146),
.B(n_142),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_152),
.A2(n_116),
.B1(n_81),
.B2(n_114),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_20),
.B1(n_33),
.B2(n_5),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_20),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_114),
.B1(n_33),
.B2(n_20),
.Y(n_171)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_114),
.C(n_33),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_181),
.C(n_130),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_0),
.Y(n_207)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_145),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_146),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_12),
.C(n_6),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_135),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_129),
.A2(n_7),
.B1(n_9),
.B2(n_13),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_154),
.C(n_151),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_188),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_128),
.Y(n_186)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_136),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_169),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_170),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_197),
.B(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_194),
.B(n_203),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_170),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_134),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_171),
.C(n_181),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_168),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_0),
.B(n_9),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_208),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_0),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_196),
.B(n_182),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_203),
.B(n_198),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_222),
.C(n_204),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_155),
.CI(n_174),
.CON(n_216),
.SN(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_186),
.B(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_200),
.B1(n_187),
.B2(n_197),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_187),
.B1(n_206),
.B2(n_198),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_157),
.B1(n_156),
.B2(n_173),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_226),
.B1(n_212),
.B2(n_210),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_159),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_225),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_167),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_191),
.Y(n_227)
);

NOR2xp67_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_163),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_184),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_13),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_231),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_232),
.B1(n_240),
.B2(n_241),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_225),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_200),
.B1(n_193),
.B2(n_190),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_190),
.C(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_236),
.C(n_237),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_195),
.C(n_205),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_195),
.C(n_172),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_221),
.B1(n_224),
.B2(n_220),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_211),
.A2(n_157),
.B1(n_169),
.B2(n_15),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_222),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_14),
.C(n_16),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_14),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_254),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_209),
.B1(n_231),
.B2(n_235),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_213),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_255),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_209),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_229),
.C(n_235),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_248),
.A2(n_215),
.B(n_243),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_260),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_234),
.B(n_215),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_213),
.B(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_251),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_242),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_266),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_250),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_273),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_261),
.A2(n_250),
.B1(n_251),
.B2(n_14),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_272),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_16),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_276),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_265),
.B(n_258),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_277),
.A2(n_268),
.B(n_185),
.C(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_279),
.B(n_274),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_278),
.Y(n_282)
);


endmodule