module fake_netlist_6_3418_n_191 (n_16, n_1, n_34, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_33, n_27, n_3, n_14, n_0, n_32, n_4, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_191);

input n_16;
input n_1;
input n_34;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_0;
input n_32;
input n_4;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_191;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_39;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_189;
wire n_85;
wire n_66;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_108;
wire n_97;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVxp33_ASAP7_75t_SL g59 ( 
.A(n_19),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_0),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

OR2x6_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_3),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_57),
.B1(n_63),
.B2(n_62),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_4),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_SL g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_5),
.Y(n_82)
);

AND3x4_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_6),
.C(n_8),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_59),
.B1(n_51),
.B2(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

AOI221xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_57),
.B1(n_51),
.B2(n_50),
.C(n_46),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_46),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_12),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NOR2x1p5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_17),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

BUFx4f_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2x1p5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_18),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_34),
.C(n_22),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_29),
.C(n_72),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_82),
.B(n_72),
.C(n_66),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_69),
.B(n_85),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_69),
.Y(n_112)
);

NOR4xp25_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_67),
.C(n_79),
.D(n_76),
.Y(n_113)
);

OAI21x1_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_75),
.B(n_71),
.Y(n_114)
);

OAI21x1_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_68),
.B(n_83),
.Y(n_115)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_95),
.Y(n_117)
);

AND2x6_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_109),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_97),
.B1(n_109),
.B2(n_93),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_107),
.C(n_89),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_104),
.B(n_100),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_87),
.B(n_95),
.Y(n_123)
);

AOI221x1_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_108),
.B1(n_106),
.B2(n_103),
.C(n_92),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_105),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_98),
.B1(n_105),
.B2(n_112),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_98),
.B(n_105),
.C(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_110),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_112),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_116),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_111),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_121),
.B1(n_120),
.B2(n_118),
.Y(n_137)
);

OAI22x1_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_83),
.B1(n_66),
.B2(n_112),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_116),
.B1(n_112),
.B2(n_88),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_125),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_99),
.B(n_124),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_110),
.Y(n_142)
);

AOI221x1_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_70),
.B1(n_55),
.B2(n_58),
.C(n_62),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_112),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_132),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

AND2x4_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_144),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_147),
.B(n_127),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

OR2x6_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_137),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_138),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_131),
.B(n_141),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_131),
.B(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_155),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_138),
.B(n_152),
.Y(n_172)
);

NOR2x1p5_ASAP7_75t_SL g173 ( 
.A(n_160),
.B(n_153),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_149),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_155),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_165),
.B(n_164),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_174),
.Y(n_179)
);

OR2x6_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_147),
.Y(n_180)
);

AOI221x1_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_172),
.B1(n_175),
.B2(n_166),
.C(n_169),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_143),
.B1(n_128),
.B2(n_159),
.C(n_158),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_176),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_181),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_180),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_183),
.B1(n_177),
.B2(n_180),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_185),
.B1(n_161),
.B2(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_188),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_143),
.B(n_161),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_161),
.B1(n_150),
.B2(n_145),
.Y(n_191)
);


endmodule