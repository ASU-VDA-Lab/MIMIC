module fake_netlist_1_11639_n_685 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_685);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_685;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx14_ASAP7_75t_R g77 ( .A(n_1), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_37), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_32), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_29), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_20), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_10), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_42), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_46), .Y(n_84) );
NOR2xp67_ASAP7_75t_L g85 ( .A(n_74), .B(n_18), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_39), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_73), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_68), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_12), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_13), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_56), .Y(n_91) );
BUFx2_ASAP7_75t_SL g92 ( .A(n_64), .Y(n_92) );
BUFx3_ASAP7_75t_L g93 ( .A(n_13), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_63), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_23), .Y(n_95) );
BUFx3_ASAP7_75t_L g96 ( .A(n_17), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_20), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_5), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_26), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_1), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_19), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_57), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_41), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_62), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_21), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_30), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_49), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_14), .Y(n_108) );
INVxp33_ASAP7_75t_L g109 ( .A(n_60), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_33), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_50), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_28), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_75), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_34), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_51), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_69), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_61), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_58), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_47), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_70), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_52), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_78), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_93), .B(n_0), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_102), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_88), .B(n_2), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_93), .Y(n_128) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_111), .B(n_113), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_78), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_102), .Y(n_131) );
INVx1_ASAP7_75t_SL g132 ( .A(n_81), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_79), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_111), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_120), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_113), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_120), .Y(n_141) );
NAND3xp33_ASAP7_75t_L g142 ( .A(n_82), .B(n_25), .C(n_72), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_86), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_81), .B(n_3), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_77), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_96), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_96), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_82), .B(n_4), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_86), .Y(n_151) );
NAND2xp33_ASAP7_75t_SL g152 ( .A(n_103), .B(n_5), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_98), .B(n_6), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_94), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_95), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_95), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_106), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_106), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_110), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_110), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_89), .B(n_6), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_112), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_129), .B(n_109), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_146), .B(n_107), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_149), .B(n_108), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_149), .B(n_123), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_136), .B(n_104), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_129), .B(n_99), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_125), .B(n_123), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_125), .B(n_89), .Y(n_180) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_128), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_129), .B(n_121), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_125), .B(n_90), .Y(n_183) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_150), .B(n_122), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
INVx5_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_125), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_138), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_156), .B(n_90), .Y(n_191) );
BUFx2_ASAP7_75t_L g192 ( .A(n_132), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_124), .B(n_91), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_124), .B(n_116), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_147), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_144), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_154), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_150), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_154), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_130), .B(n_100), .Y(n_203) );
INVxp67_ASAP7_75t_SL g204 ( .A(n_130), .Y(n_204) );
BUFx2_ASAP7_75t_L g205 ( .A(n_145), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_152), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_133), .B(n_122), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_154), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_154), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_164), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_164), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_164), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_148), .Y(n_214) );
NOR2xp33_ASAP7_75t_SL g215 ( .A(n_142), .B(n_119), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_133), .B(n_118), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_134), .B(n_118), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_134), .B(n_115), .Y(n_218) );
INVx4_ASAP7_75t_SL g219 ( .A(n_135), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_126), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_135), .B(n_115), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_137), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_126), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_137), .B(n_114), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_131), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_131), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_222), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_201), .Y(n_228) );
AND2x6_ASAP7_75t_L g229 ( .A(n_211), .B(n_140), .Y(n_229) );
CKINVDCx6p67_ASAP7_75t_R g230 ( .A(n_192), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_211), .A2(n_157), .B(n_163), .Y(n_231) );
INVx4_ASAP7_75t_L g232 ( .A(n_219), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_222), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_167), .B(n_127), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_184), .A2(n_165), .B1(n_163), .B2(n_162), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_184), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_192), .B(n_165), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_197), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_172), .Y(n_239) );
INVx4_ASAP7_75t_L g240 ( .A(n_219), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_204), .B(n_162), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_191), .B(n_161), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_182), .B(n_139), .Y(n_243) );
OR2x2_ASAP7_75t_SL g244 ( .A(n_168), .B(n_97), .Y(n_244) );
INVx5_ASAP7_75t_L g245 ( .A(n_189), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_184), .B(n_161), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_212), .A2(n_139), .B(n_159), .C(n_158), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_166), .B(n_155), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_210), .B(n_143), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_201), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_212), .B(n_155), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_174), .B(n_153), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_181), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_196), .Y(n_254) );
AND2x2_ASAP7_75t_SL g255 ( .A(n_197), .B(n_97), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_196), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_196), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_214), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_179), .A2(n_143), .B1(n_159), .B2(n_158), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_214), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_225), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_214), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_172), .Y(n_263) );
BUFx4f_ASAP7_75t_L g264 ( .A(n_179), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_172), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_220), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_220), .Y(n_267) );
AND2x6_ASAP7_75t_L g268 ( .A(n_174), .B(n_114), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_173), .B(n_157), .Y(n_269) );
NOR2x1_ASAP7_75t_L g270 ( .A(n_168), .B(n_153), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_205), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_174), .B(n_151), .Y(n_272) );
INVx5_ASAP7_75t_L g273 ( .A(n_189), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_179), .Y(n_274) );
AND2x2_ASAP7_75t_SL g275 ( .A(n_189), .B(n_105), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_201), .B(n_151), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_225), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_205), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_179), .A2(n_160), .B1(n_105), .B2(n_101), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_180), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_176), .B(n_160), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_169), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_180), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_180), .A2(n_101), .B1(n_141), .B2(n_112), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_180), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_169), .Y(n_286) );
AND2x4_ASAP7_75t_SL g287 ( .A(n_191), .B(n_141), .Y(n_287) );
INVx4_ASAP7_75t_L g288 ( .A(n_219), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_174), .B(n_80), .Y(n_289) );
OR2x6_ASAP7_75t_SL g290 ( .A(n_206), .B(n_7), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_189), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g292 ( .A1(n_282), .A2(n_203), .B1(n_193), .B2(n_216), .C(n_207), .Y(n_292) );
NOR2xp67_ASAP7_75t_SL g293 ( .A(n_236), .B(n_201), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_286), .B(n_183), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_266), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_229), .A2(n_183), .B1(n_177), .B2(n_213), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_236), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_242), .B(n_183), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_236), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_230), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_251), .A2(n_213), .B(n_177), .Y(n_301) );
AOI21xp5_ASAP7_75t_SL g302 ( .A1(n_235), .A2(n_183), .B(n_224), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_229), .A2(n_177), .B1(n_213), .B2(n_225), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_267), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_246), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_232), .Y(n_307) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_247), .A2(n_221), .B(n_218), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_228), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_271), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_274), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_228), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_229), .A2(n_213), .B1(n_177), .B2(n_175), .Y(n_313) );
CKINVDCx6p67_ASAP7_75t_R g314 ( .A(n_275), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_237), .B(n_195), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_227), .B(n_219), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_245), .Y(n_317) );
OAI22xp33_ASAP7_75t_L g318 ( .A1(n_278), .A2(n_226), .B1(n_223), .B2(n_217), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_280), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_238), .A2(n_226), .B1(n_223), .B2(n_175), .C(n_117), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_242), .B(n_226), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_283), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_287), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_233), .B(n_175), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_235), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_232), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_245), .Y(n_328) );
INVx2_ASAP7_75t_SL g329 ( .A(n_245), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_250), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_243), .A2(n_223), .B(n_226), .C(n_215), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_229), .A2(n_85), .B1(n_92), .B2(n_219), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_264), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_255), .Y(n_334) );
NAND2x2_ASAP7_75t_L g335 ( .A(n_290), .B(n_92), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_273), .B(n_187), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_259), .B(n_187), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_273), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_250), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_252), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_259), .B(n_187), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_326), .A2(n_264), .B1(n_284), .B2(n_279), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_305), .A2(n_284), .B1(n_279), .B2(n_251), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_328), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_314), .A2(n_241), .B1(n_270), .B2(n_269), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_315), .A2(n_248), .B1(n_268), .B2(n_281), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_314), .A2(n_234), .B1(n_249), .B2(n_268), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_301), .A2(n_252), .B(n_272), .Y(n_348) );
NOR4xp25_ASAP7_75t_L g349 ( .A(n_318), .B(n_289), .C(n_272), .D(n_244), .Y(n_349) );
AOI22xp33_ASAP7_75t_SL g350 ( .A1(n_334), .A2(n_268), .B1(n_289), .B2(n_273), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_321), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_340), .A2(n_268), .B1(n_253), .B2(n_231), .Y(n_352) );
CKINVDCx11_ASAP7_75t_R g353 ( .A(n_310), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_331), .A2(n_257), .B(n_258), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_300), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_321), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_302), .A2(n_276), .B(n_291), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g358 ( .A1(n_292), .A2(n_254), .B1(n_262), .B2(n_256), .C(n_260), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_310), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_307), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_296), .B(n_277), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_300), .Y(n_362) );
NAND2xp33_ASAP7_75t_L g363 ( .A(n_305), .B(n_261), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_340), .B(n_277), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_298), .A2(n_277), .B1(n_261), .B2(n_265), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g366 ( .A1(n_335), .A2(n_261), .B1(n_263), .B2(n_239), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_328), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_295), .Y(n_368) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_335), .A2(n_288), .B1(n_240), .B2(n_187), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_306), .A2(n_288), .B1(n_240), .B2(n_194), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_306), .A2(n_187), .B1(n_170), .B2(n_194), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_323), .B(n_7), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_368), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_342), .A2(n_295), .B1(n_304), .B2(n_332), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_349), .A2(n_303), .B(n_313), .C(n_302), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_343), .A2(n_304), .B1(n_294), .B2(n_298), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_345), .A2(n_308), .B1(n_322), .B2(n_311), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_351), .Y(n_378) );
OAI211xp5_ASAP7_75t_SL g379 ( .A1(n_353), .A2(n_320), .B(n_311), .C(n_319), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g380 ( .A1(n_359), .A2(n_333), .B1(n_328), .B2(n_338), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_346), .A2(n_333), .B1(n_325), .B2(n_322), .C(n_324), .Y(n_381) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_347), .A2(n_319), .B1(n_324), .B2(n_341), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_372), .B(n_317), .Y(n_383) );
OAI211xp5_ASAP7_75t_L g384 ( .A1(n_366), .A2(n_338), .B(n_329), .C(n_317), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_344), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_356), .B(n_329), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_344), .B(n_338), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_346), .A2(n_308), .B1(n_337), .B2(n_312), .Y(n_389) );
AOI222xp33_ASAP7_75t_L g390 ( .A1(n_353), .A2(n_339), .B1(n_309), .B2(n_330), .C1(n_312), .C2(n_293), .Y(n_390) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_363), .B(n_293), .C(n_198), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_355), .B(n_336), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_362), .A2(n_308), .B1(n_297), .B2(n_299), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_361), .A2(n_339), .B1(n_309), .B2(n_330), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_367), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_361), .A2(n_297), .B1(n_299), .B2(n_316), .Y(n_397) );
BUFx2_ASAP7_75t_SL g398 ( .A(n_360), .Y(n_398) );
OR2x6_ASAP7_75t_L g399 ( .A(n_357), .B(n_336), .Y(n_399) );
OAI21xp33_ASAP7_75t_L g400 ( .A1(n_377), .A2(n_352), .B(n_350), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_388), .A2(n_369), .B1(n_348), .B2(n_352), .C(n_364), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_376), .A2(n_365), .B1(n_364), .B2(n_370), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_373), .Y(n_403) );
AOI211xp5_ASAP7_75t_SL g404 ( .A1(n_374), .A2(n_297), .B(n_299), .C(n_371), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_392), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_373), .Y(n_406) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_384), .B(n_360), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_378), .B(n_365), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_374), .A2(n_360), .B1(n_316), .B2(n_327), .Y(n_409) );
OR2x6_ASAP7_75t_L g410 ( .A(n_399), .B(n_354), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_379), .A2(n_198), .B1(n_185), .B2(n_170), .C(n_199), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_387), .B(n_8), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_394), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_387), .Y(n_415) );
OAI211xp5_ASAP7_75t_L g416 ( .A1(n_393), .A2(n_185), .B(n_200), .C(n_199), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_394), .Y(n_417) );
OA21x2_ASAP7_75t_L g418 ( .A1(n_389), .A2(n_171), .B(n_200), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_396), .B(n_336), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_377), .A2(n_316), .B1(n_327), .B2(n_307), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_389), .B(n_178), .C(n_186), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_381), .A2(n_316), .B1(n_327), .B2(n_307), .Y(n_422) );
OAI211xp5_ASAP7_75t_L g423 ( .A1(n_380), .A2(n_187), .B(n_209), .C(n_208), .Y(n_423) );
OAI22xp5_ASAP7_75t_SL g424 ( .A1(n_397), .A2(n_327), .B1(n_307), .B2(n_336), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_386), .B(n_8), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_387), .B(n_9), .Y(n_426) );
AO21x2_ASAP7_75t_L g427 ( .A1(n_382), .A2(n_171), .B(n_209), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_390), .B(n_178), .C(n_186), .Y(n_428) );
OR2x6_ASAP7_75t_L g429 ( .A(n_399), .B(n_327), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_382), .A2(n_209), .B1(n_202), .B2(n_208), .C(n_190), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_385), .B(n_9), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_399), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_385), .Y(n_433) );
INVx4_ASAP7_75t_R g434 ( .A(n_398), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_403), .B(n_395), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_429), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_403), .B(n_395), .Y(n_437) );
OAI22xp5_ASAP7_75t_SL g438 ( .A1(n_424), .A2(n_375), .B1(n_391), .B2(n_12), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_424), .A2(n_307), .B1(n_202), .B2(n_190), .Y(n_439) );
OAI31xp33_ASAP7_75t_L g440 ( .A1(n_404), .A2(n_10), .A3(n_11), .B(n_14), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_415), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_406), .Y(n_442) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_421), .A2(n_190), .B(n_188), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_429), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_428), .B(n_190), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_412), .Y(n_446) );
BUFx2_ASAP7_75t_L g447 ( .A(n_410), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_406), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_432), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_432), .Y(n_450) );
NAND3xp33_ASAP7_75t_SL g451 ( .A(n_425), .B(n_11), .C(n_15), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_410), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_410), .B(n_15), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_410), .B(n_16), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_427), .B(n_16), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_433), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_431), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_427), .B(n_17), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_408), .B(n_18), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_415), .B(n_19), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_427), .B(n_21), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_414), .B(n_190), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_425), .B(n_190), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_418), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_418), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_414), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_417), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_400), .A2(n_188), .B1(n_186), .B2(n_178), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_417), .B(n_188), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_418), .Y(n_470) );
OAI31xp33_ASAP7_75t_L g471 ( .A1(n_400), .A2(n_22), .A3(n_24), .B(n_27), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_418), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_415), .B(n_188), .Y(n_473) );
NAND3xp33_ASAP7_75t_L g474 ( .A(n_426), .B(n_188), .C(n_186), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_413), .B(n_188), .Y(n_475) );
INVx5_ASAP7_75t_SL g476 ( .A(n_429), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_405), .B(n_31), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_413), .B(n_186), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_429), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_431), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_419), .B(n_35), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_419), .B(n_409), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_422), .A2(n_186), .B1(n_178), .B2(n_40), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_401), .A2(n_178), .B(n_38), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_464), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_446), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_449), .B(n_420), .Y(n_487) );
OAI33xp33_ASAP7_75t_L g488 ( .A1(n_459), .A2(n_402), .A3(n_421), .B1(n_434), .B2(n_416), .B3(n_411), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_445), .A2(n_484), .B(n_474), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_456), .B(n_407), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_456), .B(n_407), .Y(n_491) );
NAND2xp33_ASAP7_75t_L g492 ( .A(n_438), .B(n_434), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_442), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_448), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_448), .Y(n_495) );
AND2x2_ASAP7_75t_SL g496 ( .A(n_447), .B(n_430), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_452), .B(n_36), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_449), .B(n_178), .Y(n_498) );
NOR3xp33_ASAP7_75t_SL g499 ( .A(n_451), .B(n_423), .C(n_44), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_451), .B(n_43), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_448), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_452), .B(n_45), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_453), .A2(n_48), .B1(n_53), .B2(n_54), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_442), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_466), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_457), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_449), .B(n_55), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_450), .B(n_59), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_480), .B(n_65), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_450), .B(n_66), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_466), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_467), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_450), .B(n_67), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_438), .A2(n_76), .B1(n_454), .B2(n_453), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_437), .B(n_452), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_480), .B(n_437), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_437), .B(n_454), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_467), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_457), .B(n_435), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_455), .B(n_461), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_455), .B(n_461), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_455), .B(n_461), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_459), .A2(n_453), .B1(n_454), .B2(n_440), .C(n_458), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_458), .B(n_479), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_464), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_458), .B(n_479), .Y(n_526) );
NAND4xp25_ASAP7_75t_L g527 ( .A(n_440), .B(n_477), .C(n_471), .D(n_447), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_470), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_460), .A2(n_481), .B1(n_436), .B2(n_444), .C(n_475), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_435), .B(n_460), .Y(n_530) );
OAI221xp5_ASAP7_75t_L g531 ( .A1(n_471), .A2(n_439), .B1(n_484), .B2(n_474), .C(n_436), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_470), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_436), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_472), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_463), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_479), .B(n_472), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_475), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_463), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_444), .B(n_478), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_475), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_464), .B(n_465), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_465), .B(n_444), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_515), .B(n_465), .Y(n_543) );
NOR3xp33_ASAP7_75t_L g544 ( .A(n_492), .B(n_478), .C(n_473), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_486), .B(n_482), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_516), .B(n_482), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_527), .B(n_441), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_492), .A2(n_439), .B1(n_476), .B2(n_478), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_485), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_533), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_504), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_519), .B(n_476), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_514), .A2(n_476), .B1(n_441), .B2(n_483), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_533), .B(n_441), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_515), .B(n_476), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_504), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_493), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_519), .B(n_476), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_506), .B(n_476), .Y(n_559) );
AOI211xp5_ASAP7_75t_L g560 ( .A1(n_523), .A2(n_473), .B(n_462), .C(n_469), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_530), .B(n_462), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_520), .B(n_443), .Y(n_562) );
AND4x1_ASAP7_75t_L g563 ( .A(n_499), .B(n_468), .C(n_462), .D(n_469), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_489), .B(n_469), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_520), .B(n_443), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_517), .B(n_443), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_488), .A2(n_443), .B1(n_521), .B2(n_522), .Y(n_567) );
NAND2xp67_ASAP7_75t_L g568 ( .A(n_521), .B(n_522), .Y(n_568) );
NOR2xp67_ASAP7_75t_L g569 ( .A(n_531), .B(n_485), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_537), .B(n_540), .Y(n_570) );
AND4x1_ASAP7_75t_L g571 ( .A(n_500), .B(n_529), .C(n_503), .D(n_490), .Y(n_571) );
XOR2xp5_ASAP7_75t_L g572 ( .A(n_539), .B(n_526), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_524), .B(n_526), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_505), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_542), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_505), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_524), .B(n_542), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_536), .B(n_528), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_511), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_535), .B(n_538), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_511), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_512), .Y(n_582) );
AOI21xp33_ASAP7_75t_SL g583 ( .A1(n_496), .A2(n_491), .B(n_512), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_501), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_536), .B(n_541), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_518), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_494), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_518), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_541), .B(n_485), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_528), .B(n_534), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_532), .B(n_534), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_494), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_532), .B(n_495), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_585), .B(n_487), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_590), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_590), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_591), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_557), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_547), .B(n_496), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_545), .B(n_495), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_585), .B(n_487), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_546), .B(n_501), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_551), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_587), .Y(n_604) );
NAND2x1_ASAP7_75t_L g605 ( .A(n_569), .B(n_497), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_578), .B(n_525), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_556), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_574), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_570), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_575), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_547), .A2(n_497), .B1(n_502), .B2(n_509), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_576), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_584), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_578), .B(n_497), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_579), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_577), .B(n_498), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_592), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_578), .B(n_498), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_580), .B(n_502), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_573), .B(n_502), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_573), .B(n_507), .Y(n_621) );
INVx2_ASAP7_75t_SL g622 ( .A(n_589), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_581), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_589), .B(n_507), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_582), .Y(n_625) );
XNOR2xp5_ASAP7_75t_L g626 ( .A(n_572), .B(n_508), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_561), .B(n_513), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_586), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_568), .B(n_513), .Y(n_629) );
XOR2x2_ASAP7_75t_L g630 ( .A(n_544), .B(n_508), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_550), .Y(n_631) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_564), .B(n_510), .Y(n_632) );
AO22x2_ASAP7_75t_L g633 ( .A1(n_550), .A2(n_510), .B1(n_588), .B2(n_552), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_593), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_584), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_564), .A2(n_560), .B(n_553), .Y(n_636) );
AOI222xp33_ASAP7_75t_L g637 ( .A1(n_567), .A2(n_562), .B1(n_565), .B2(n_543), .C1(n_555), .C2(n_554), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_548), .A2(n_567), .B1(n_562), .B2(n_565), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_543), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_552), .Y(n_640) );
INVx2_ASAP7_75t_SL g641 ( .A(n_559), .Y(n_641) );
CKINVDCx5p33_ASAP7_75t_R g642 ( .A(n_559), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_558), .Y(n_643) );
XNOR2x2_ASAP7_75t_L g644 ( .A(n_566), .B(n_555), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_583), .A2(n_566), .B1(n_549), .B2(n_554), .C(n_571), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_549), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_554), .A2(n_549), .B(n_563), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_590), .Y(n_648) );
NOR2x1_ASAP7_75t_L g649 ( .A(n_569), .B(n_492), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_569), .B(n_544), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_599), .A2(n_649), .B1(n_650), .B2(n_636), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_610), .B(n_606), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_645), .A2(n_609), .B1(n_633), .B2(n_597), .C(n_638), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_617), .Y(n_654) );
NOR4xp75_ASAP7_75t_L g655 ( .A(n_605), .B(n_629), .C(n_614), .D(n_631), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_637), .B(n_638), .Y(n_656) );
NOR2xp33_ASAP7_75t_R g657 ( .A(n_626), .B(n_642), .Y(n_657) );
INVxp67_ASAP7_75t_SL g658 ( .A(n_644), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_633), .A2(n_605), .B(n_626), .Y(n_659) );
AOI21xp33_ASAP7_75t_L g660 ( .A1(n_637), .A2(n_617), .B(n_604), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_632), .A2(n_647), .B(n_630), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_640), .A2(n_643), .B1(n_622), .B2(n_641), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_604), .A2(n_600), .B(n_602), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_654), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_658), .A2(n_611), .B1(n_634), .B2(n_622), .C(n_598), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_659), .B(n_618), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_653), .A2(n_620), .B(n_616), .C(n_618), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_656), .B(n_646), .C(n_608), .Y(n_668) );
AND4x2_ASAP7_75t_L g669 ( .A(n_651), .B(n_620), .C(n_594), .D(n_601), .Y(n_669) );
AO22x2_ASAP7_75t_L g670 ( .A1(n_661), .A2(n_603), .B1(n_615), .B2(n_625), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_663), .B(n_594), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_664), .Y(n_672) );
OAI211xp5_ASAP7_75t_SL g673 ( .A1(n_666), .A2(n_660), .B(n_662), .C(n_652), .Y(n_673) );
NAND5xp2_ASAP7_75t_L g674 ( .A(n_667), .B(n_655), .C(n_657), .D(n_619), .E(n_624), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_665), .A2(n_668), .B1(n_671), .B2(n_669), .C(n_670), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_674), .B(n_595), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_672), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_673), .B(n_670), .Y(n_678) );
NOR2xp67_ASAP7_75t_L g679 ( .A(n_677), .B(n_675), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_676), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_679), .A2(n_678), .B1(n_596), .B2(n_648), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_680), .B(n_628), .Y(n_682) );
AOI222xp33_ASAP7_75t_L g683 ( .A1(n_681), .A2(n_623), .B1(n_607), .B2(n_612), .C1(n_601), .C2(n_639), .Y(n_683) );
OAI22xp33_ASAP7_75t_L g684 ( .A1(n_683), .A2(n_682), .B1(n_621), .B2(n_627), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_684), .A2(n_635), .B(n_613), .Y(n_685) );
endmodule