module fake_jpeg_22260_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_30),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_0),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_33),
.Y(n_37)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_27),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_17),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_19),
.B1(n_22),
.B2(n_13),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_26),
.B1(n_19),
.B2(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_14),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_43),
.B1(n_35),
.B2(n_13),
.Y(n_76)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_59),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_28),
.B(n_31),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_40),
.B(n_24),
.Y(n_62)
);

NOR4xp25_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_28),
.C(n_17),
.D(n_21),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_55),
.B(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_28),
.B(n_20),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

OR2x2_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_13),
.Y(n_58)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_43),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_53),
.C(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_52),
.B1(n_51),
.B2(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_86),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_52),
.B1(n_58),
.B2(n_50),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_76),
.B1(n_63),
.B2(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_87),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_91),
.B1(n_70),
.B2(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_92),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_68),
.B(n_64),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_100),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_102),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_90),
.B(n_68),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_80),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_79),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_79),
.C(n_92),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_96),
.C(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_93),
.B(n_73),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_95),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_117),
.C(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_111),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_114),
.B(n_96),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_106),
.B(n_91),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_112),
.B(n_121),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_127),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_126),
.C(n_15),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_103),
.B1(n_117),
.B2(n_61),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_131),
.C(n_132),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_7),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_12),
.A3(n_6),
.B1(n_11),
.B2(n_3),
.C1(n_5),
.C2(n_9),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_136),
.C(n_0),
.Y(n_137)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_6),
.A3(n_8),
.B1(n_24),
.B2(n_0),
.C1(n_1),
.C2(n_2),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.C(n_135),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_139),
.Y(n_140)
);


endmodule