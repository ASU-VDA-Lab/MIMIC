module real_jpeg_24117_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_210;
wire n_127;
wire n_53;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_2),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_2),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_2),
.B(n_66),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_2),
.B(n_35),
.C(n_37),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_28),
.B1(n_30),
.B2(n_69),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_2),
.B(n_40),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_69),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_2),
.B(n_48),
.C(n_50),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_2),
.A2(n_79),
.B(n_171),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_4),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_5),
.A2(n_42),
.B1(n_48),
.B2(n_51),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_6),
.A2(n_48),
.B1(n_51),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_83),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_8),
.A2(n_56),
.B1(n_68),
.B2(n_75),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_56),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_8),
.A2(n_48),
.B1(n_51),
.B2(n_56),
.Y(n_140)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_48),
.B1(n_51),
.B2(n_87),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_10),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_11),
.A2(n_46),
.B1(n_48),
.B2(n_51),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_12),
.A2(n_48),
.B1(n_51),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_12),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_14),
.A2(n_27),
.B1(n_68),
.B2(n_109),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_14),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_14),
.A2(n_27),
.B1(n_48),
.B2(n_51),
.Y(n_183)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_15),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_99),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_20),
.B(n_99),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.C(n_90),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_21),
.A2(n_22),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_44),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_25),
.B(n_43),
.C(n_57),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_26),
.Y(n_92)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_28),
.A2(n_30),
.B1(n_61),
.B2(n_62),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_28),
.B(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_28),
.B(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g88 ( 
.A1(n_30),
.A2(n_62),
.A3(n_64),
.B1(n_71),
.B2(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_31),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_32),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_32),
.A2(n_105),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_33),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_35),
.B(n_178),
.Y(n_177)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_40),
.B(n_94),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_41),
.Y(n_104)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_52),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_45),
.A2(n_47),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_47),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_47),
.A2(n_52),
.B(n_143),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_47),
.B(n_69),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_51),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_53),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_55),
.B(n_145),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_67),
.B(n_73),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_59)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_107),
.B(n_111),
.Y(n_106)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_67)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_69),
.B(n_85),
.Y(n_195)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_76),
.B(n_90),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_88),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_88),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_84),
.B2(n_86),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_78),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_79),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_80),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_97),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_91),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_113),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_124),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_122),
.A2(n_159),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_207),
.B(n_212),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_160),
.B(n_206),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_149),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_130),
.B(n_149),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_141),
.C(n_146),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_131),
.B(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_134),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B(n_139),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_183),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_139),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_141),
.A2(n_146),
.B1(n_147),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_150),
.B(n_156),
.C(n_157),
.Y(n_211)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_200),
.B(n_205),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_179),
.B(n_199),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_173),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_173),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_170),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_177),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_188),
.B(n_198),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_186),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_193),
.B(n_197),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_204),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_211),
.Y(n_212)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);


endmodule