module fake_netlist_6_3607_n_107 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_107);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_107;

wire n_52;
wire n_91;
wire n_46;
wire n_18;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVxp33_ASAP7_75t_SL g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx8_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_18),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_43)
);

OAI221xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_20),
.B1(n_30),
.B2(n_23),
.C(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_31),
.B1(n_21),
.B2(n_30),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_31),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_34),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_48),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_50),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_50),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_65),
.Y(n_67)
);

AND2x4_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_58),
.Y(n_68)
);

AND2x4_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_58),
.Y(n_69)
);

AOI221xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_43),
.B1(n_44),
.B2(n_62),
.C(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_62),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_64),
.B(n_66),
.C(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

OAI211xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_41),
.B(n_36),
.C(n_38),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_67),
.B1(n_69),
.B2(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_68),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_64),
.B1(n_63),
.B2(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_76),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_38),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_82),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_75),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_81),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_90),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_95),
.Y(n_96)
);

OR4x1_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_51),
.C(n_3),
.D(n_4),
.Y(n_97)
);

NOR2x1p5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_89),
.B1(n_41),
.B2(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_98),
.Y(n_100)
);

AOI221xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_42),
.B1(n_89),
.B2(n_8),
.C(n_9),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_42),
.B1(n_53),
.B2(n_52),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_2),
.Y(n_103)
);

OAI322xp33_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_103),
.A3(n_99),
.B1(n_10),
.B2(n_11),
.C1(n_6),
.C2(n_8),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_10),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_14),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_104),
.B1(n_55),
.B2(n_71),
.C(n_63),
.Y(n_107)
);


endmodule