module fake_jpeg_28711_n_505 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_505);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_505;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_53),
.B(n_72),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_16),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_77),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_38),
.Y(n_67)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_71),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_40),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_74),
.B(n_42),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_30),
.B(n_8),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_90),
.Y(n_132)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_32),
.B(n_9),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_100),
.Y(n_119)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

CKINVDCx9p33_ASAP7_75t_R g106 ( 
.A(n_57),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g175 ( 
.A(n_106),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_141),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_62),
.A2(n_67),
.B1(n_90),
.B2(n_20),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_109),
.A2(n_145),
.B1(n_89),
.B2(n_92),
.Y(n_194)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_26),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_57),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_79),
.A2(n_43),
.B1(n_50),
.B2(n_45),
.Y(n_145)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_54),
.Y(n_152)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_160),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_65),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_161),
.B(n_164),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_74),
.B1(n_66),
.B2(n_56),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_163),
.B(n_132),
.Y(n_213)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_168),
.Y(n_253)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_170),
.B(n_174),
.Y(n_245)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_171),
.Y(n_219)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_119),
.B(n_64),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_102),
.A2(n_137),
.B1(n_68),
.B2(n_85),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_177),
.B(n_187),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_179),
.Y(n_229)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_74),
.B(n_99),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_181),
.A2(n_60),
.B(n_24),
.Y(n_255)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_182),
.B(n_184),
.Y(n_251)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_118),
.A2(n_101),
.B1(n_98),
.B2(n_97),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_202),
.B1(n_149),
.B2(n_159),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_158),
.A2(n_95),
.B1(n_88),
.B2(n_61),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_186),
.A2(n_196),
.B1(n_207),
.B2(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_121),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_201),
.C(n_29),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_133),
.B(n_34),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_189),
.B(n_211),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_34),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_195),
.Y(n_241)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_194),
.A2(n_33),
.B1(n_48),
.B2(n_51),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_109),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_158),
.A2(n_60),
.B1(n_61),
.B2(n_78),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_44),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_198),
.Y(n_234)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_103),
.Y(n_199)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_124),
.B(n_140),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_145),
.A2(n_70),
.B1(n_82),
.B2(n_76),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_132),
.A2(n_32),
.B1(n_44),
.B2(n_49),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_51),
.B(n_48),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_205),
.Y(n_237)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_206),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_87),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_208),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_134),
.B(n_49),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_147),
.B(n_87),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_217),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_214),
.A2(n_122),
.B1(n_112),
.B2(n_144),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_108),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_75),
.B1(n_73),
.B2(n_58),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_231),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_104),
.B1(n_146),
.B2(n_135),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_227),
.B(n_243),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_163),
.B(n_181),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_163),
.B(n_33),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_232),
.B(n_238),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_147),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_177),
.B(n_114),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_166),
.B(n_29),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_168),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_185),
.A2(n_108),
.B1(n_144),
.B2(n_142),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_244),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_209),
.A2(n_134),
.B1(n_50),
.B2(n_25),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_248),
.A2(n_167),
.B(n_190),
.Y(n_287)
);

OR2x2_ASAP7_75t_SL g257 ( 
.A(n_255),
.B(n_186),
.Y(n_257)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_256),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_257),
.A2(n_280),
.B(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_253),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_246),
.Y(n_304)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_259),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_270),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_262),
.B(n_267),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_251),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_263),
.Y(n_317)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_199),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_268),
.A2(n_219),
.B1(n_114),
.B2(n_127),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_187),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_160),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_217),
.B(n_180),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_285),
.Y(n_300)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_216),
.B(n_160),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_282),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_231),
.B(n_236),
.C(n_213),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_279),
.C(n_292),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_165),
.C(n_205),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_238),
.A2(n_196),
.B(n_16),
.C(n_9),
.Y(n_280)
);

INVx2_ASAP7_75t_R g281 ( 
.A(n_233),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_281),
.A2(n_248),
.B(n_222),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g282 ( 
.A(n_228),
.B(n_216),
.C(n_241),
.Y(n_282)
);

CKINVDCx10_ASAP7_75t_R g283 ( 
.A(n_229),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_283),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_228),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_284),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_245),
.Y(n_285)
);

AND2x6_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_175),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_287),
.A2(n_240),
.B(n_244),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_200),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_229),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_165),
.C(n_191),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

AO22x2_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_214),
.B1(n_243),
.B2(n_233),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_313),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_264),
.A2(n_232),
.B1(n_224),
.B2(n_230),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_302),
.A2(n_311),
.B1(n_280),
.B2(n_258),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_242),
.C(n_226),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_320),
.C(n_266),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_312),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_264),
.A2(n_290),
.B1(n_291),
.B2(n_289),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_242),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_290),
.A2(n_249),
.B1(n_207),
.B2(n_123),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_325),
.B1(n_329),
.B2(n_175),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_269),
.B(n_281),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_318),
.B(n_257),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_287),
.A2(n_237),
.B(n_249),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_319),
.A2(n_321),
.B(n_323),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_220),
.C(n_223),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_246),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_288),
.A2(n_250),
.B(n_220),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_263),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_283),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_276),
.A2(n_122),
.B1(n_112),
.B2(n_142),
.Y(n_325)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_330),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_331),
.A2(n_335),
.B1(n_361),
.B2(n_321),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_302),
.A2(n_285),
.B1(n_273),
.B2(n_262),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_317),
.B(n_292),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_336),
.B(n_339),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_307),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_345),
.Y(n_362)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_338),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_250),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_260),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_340),
.B(n_342),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_279),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_351),
.C(n_223),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_260),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_360),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_307),
.Y(n_345)
);

INVx13_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_265),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_347),
.B(n_359),
.Y(n_369)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_348),
.Y(n_385)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_316),
.Y(n_349)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_328),
.B(n_272),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_350),
.B(n_355),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_310),
.B(n_286),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_352),
.B(n_294),
.Y(n_368)
);

CKINVDCx10_ASAP7_75t_R g354 ( 
.A(n_327),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_354),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_299),
.B(n_237),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_316),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_356),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_265),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_357),
.B(n_301),
.Y(n_390)
);

CKINVDCx10_ASAP7_75t_R g358 ( 
.A(n_327),
.Y(n_358)
);

OAI21x1_ASAP7_75t_R g384 ( 
.A1(n_358),
.A2(n_179),
.B(n_304),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_298),
.B(n_303),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_313),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_332),
.A2(n_319),
.B(n_294),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_363),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_306),
.B(n_311),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_366),
.B(n_368),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_333),
.A2(n_321),
.B(n_312),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_370),
.B(n_383),
.Y(n_415)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_373),
.A2(n_382),
.B1(n_358),
.B2(n_356),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_361),
.A2(n_301),
.B1(n_318),
.B2(n_329),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_375),
.A2(n_386),
.B1(n_190),
.B2(n_167),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_320),
.Y(n_376)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_376),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_346),
.B(n_296),
.Y(n_379)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_379),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_300),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_381),
.B(n_389),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_354),
.A2(n_295),
.B1(n_326),
.B2(n_309),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_323),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_384),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_333),
.A2(n_301),
.B1(n_305),
.B2(n_304),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_344),
.B(n_301),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_343),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_305),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_390),
.A2(n_337),
.B1(n_348),
.B2(n_275),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_333),
.C(n_353),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_365),
.B(n_351),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_395),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_383),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_347),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_414),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_402),
.C(n_406),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_334),
.C(n_353),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_375),
.A2(n_334),
.B1(n_343),
.B2(n_349),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_403),
.A2(n_408),
.B1(n_411),
.B2(n_384),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_404),
.A2(n_416),
.B1(n_384),
.B2(n_364),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_330),
.C(n_338),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_293),
.C(n_345),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_412),
.C(n_364),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_373),
.A2(n_259),
.B1(n_256),
.B2(n_221),
.Y(n_409)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_409),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_378),
.A2(n_50),
.B1(n_116),
.B2(n_127),
.Y(n_410)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_410),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_388),
.A2(n_215),
.B1(n_221),
.B2(n_218),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_369),
.B(n_215),
.C(n_218),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_386),
.A2(n_116),
.B1(n_123),
.B2(n_247),
.Y(n_413)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_366),
.B(n_370),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_418),
.B(n_419),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_420),
.B(n_424),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_431),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_401),
.A2(n_403),
.B1(n_392),
.B2(n_397),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_428),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_363),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_415),
.Y(n_425)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_425),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_394),
.A2(n_377),
.B1(n_371),
.B2(n_374),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_416),
.A2(n_368),
.B1(n_362),
.B2(n_380),
.Y(n_429)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_429),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_377),
.C(n_374),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_430),
.B(n_407),
.C(n_414),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_387),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_387),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_433),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_396),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_405),
.B(n_380),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_436),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_446),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_399),
.C(n_402),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_440),
.C(n_444),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_412),
.C(n_393),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_435),
.A2(n_393),
.B(n_367),
.Y(n_441)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_441),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_411),
.C(n_367),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_430),
.A2(n_385),
.B(n_169),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_448),
.B(n_418),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_385),
.C(n_191),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_449),
.B(n_451),
.C(n_431),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_197),
.C(n_169),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_447),
.A2(n_429),
.B1(n_420),
.B2(n_423),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_455),
.A2(n_465),
.B1(n_450),
.B2(n_15),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g457 ( 
.A(n_445),
.B(n_424),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_14),
.Y(n_477)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_458),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_432),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_463),
.C(n_466),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_434),
.Y(n_460)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_460),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_462),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_442),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_179),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g464 ( 
.A1(n_439),
.A2(n_197),
.B1(n_13),
.B2(n_14),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_464),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_444),
.A2(n_25),
.B1(n_10),
.B2(n_16),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_437),
.B(n_15),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_28),
.C(n_24),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_24),
.C(n_28),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_468),
.A2(n_438),
.B1(n_449),
.B2(n_439),
.Y(n_469)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_454),
.A2(n_451),
.B(n_453),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_470),
.A2(n_477),
.B(n_479),
.Y(n_490)
);

INVx6_ASAP7_75t_L g473 ( 
.A(n_456),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_473),
.A2(n_456),
.B1(n_461),
.B2(n_459),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_476),
.B(n_478),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_455),
.A2(n_2),
.B(n_3),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_467),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_481),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_463),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_483),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_466),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_485),
.B(n_486),
.Y(n_492)
);

O2A1O1Ixp33_ASAP7_75t_L g486 ( 
.A1(n_472),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_473),
.A2(n_4),
.B(n_6),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_489),
.A2(n_477),
.B1(n_490),
.B2(n_479),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_487),
.A2(n_474),
.B1(n_475),
.B2(n_470),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_494),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_482),
.C(n_485),
.Y(n_498)
);

O2A1O1Ixp33_ASAP7_75t_SL g497 ( 
.A1(n_491),
.A2(n_486),
.B(n_488),
.C(n_484),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_498),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_496),
.B(n_493),
.C(n_492),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_499),
.B(n_481),
.Y(n_501)
);

OAI211xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_500),
.B(n_4),
.C(n_28),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_24),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_503),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_504),
.B(n_28),
.Y(n_505)
);


endmodule