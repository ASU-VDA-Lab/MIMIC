module fake_netlist_6_1292_n_788 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_788);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_788;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_154),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_26),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_40),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_10),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_28),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_7),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_80),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_122),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_59),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_147),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_30),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_108),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_103),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_69),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_101),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_4),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_56),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_42),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_8),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_49),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_72),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_57),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_152),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_6),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_96),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_25),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_109),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_92),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_79),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_94),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_8),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_74),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_9),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_31),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_29),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_6),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_3),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_L g209 ( 
.A(n_102),
.B(n_104),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_15),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_85),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_58),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_162),
.B(n_16),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_0),
.Y(n_217)
);

CKINVDCx8_ASAP7_75t_R g218 ( 
.A(n_205),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_1),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

CKINVDCx6p67_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_2),
.Y(n_222)
);

OAI22x1_ASAP7_75t_R g223 ( 
.A1(n_164),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_166),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

CKINVDCx11_ASAP7_75t_R g228 ( 
.A(n_181),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

AOI22x1_ASAP7_75t_SL g231 ( 
.A1(n_179),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

BUFx8_ASAP7_75t_SL g233 ( 
.A(n_181),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_159),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_191),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g239 ( 
.A1(n_162),
.A2(n_11),
.B(n_12),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

BUFx8_ASAP7_75t_L g241 ( 
.A(n_165),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_163),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_165),
.B(n_170),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_12),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_169),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_13),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_173),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_174),
.Y(n_254)
);

OA21x2_ASAP7_75t_L g255 ( 
.A1(n_177),
.A2(n_13),
.B(n_14),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_168),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_233),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_256),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_251),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_185),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_233),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_251),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_186),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_228),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_171),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_237),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_228),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_218),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_249),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_237),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_221),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_250),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_241),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_220),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_224),
.B(n_172),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_227),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_220),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_188),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_241),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_196),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_244),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_229),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_R g292 ( 
.A(n_254),
.B(n_175),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_229),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_229),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_230),
.B(n_176),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_215),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_230),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_230),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_254),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_245),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_232),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_232),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_247),
.Y(n_306)
);

AO221x1_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_202),
.B1(n_211),
.B2(n_206),
.C(n_210),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_304),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_240),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_240),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_286),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_292),
.B(n_217),
.Y(n_315)
);

NAND2xp33_ASAP7_75t_SL g316 ( 
.A(n_292),
.B(n_248),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_260),
.B(n_302),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_291),
.B(n_217),
.Y(n_320)
);

NAND2x1p5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_239),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_268),
.Y(n_322)
);

NOR3xp33_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_248),
.C(n_215),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_298),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_294),
.B(n_219),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_L g329 ( 
.A(n_258),
.B(n_243),
.C(n_252),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_219),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_272),
.B(n_187),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_SL g333 ( 
.A(n_296),
.B(n_222),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_274),
.B(n_262),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_L g335 ( 
.A(n_269),
.B(n_253),
.C(n_236),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_222),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_264),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_L g341 ( 
.A(n_276),
.B(n_216),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_265),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_275),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_214),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_259),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_271),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_284),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_285),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_266),
.B(n_242),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_263),
.B(n_235),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_289),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_263),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_287),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_273),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_280),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_278),
.B(n_252),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_257),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_278),
.B(n_216),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_L g363 ( 
.A(n_288),
.B(n_214),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_267),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_261),
.B(n_247),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_270),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_281),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_295),
.B(n_216),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_292),
.B(n_178),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_295),
.B(n_216),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_308),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_306),
.B(n_247),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_339),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_317),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_312),
.Y(n_376)
);

A2O1A1Ixp33_ASAP7_75t_SL g377 ( 
.A1(n_336),
.A2(n_214),
.B(n_255),
.C(n_239),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_331),
.B(n_223),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_R g379 ( 
.A(n_343),
.B(n_182),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_214),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_306),
.B(n_318),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_323),
.A2(n_255),
.B1(n_209),
.B2(n_213),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_318),
.B(n_190),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_192),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_367),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_323),
.A2(n_212),
.B1(n_200),
.B2(n_198),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_344),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_337),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_314),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_321),
.A2(n_197),
.B1(n_194),
.B2(n_193),
.Y(n_391)
);

OR2x2_ASAP7_75t_SL g392 ( 
.A(n_361),
.B(n_231),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_321),
.A2(n_84),
.B(n_17),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g394 ( 
.A(n_309),
.B(n_18),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_346),
.B(n_14),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_19),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_R g398 ( 
.A(n_316),
.B(n_20),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_329),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_330),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_311),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_315),
.A2(n_322),
.B1(n_320),
.B2(n_326),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_310),
.B(n_24),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_340),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_329),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_359),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_352),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_347),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_334),
.B(n_34),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_324),
.B(n_35),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_338),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_354),
.B(n_341),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_328),
.B(n_36),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_328),
.B(n_37),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_319),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_354),
.B(n_38),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_325),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_325),
.B(n_327),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_319),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_362),
.B(n_365),
.Y(n_423)
);

OR2x6_ASAP7_75t_L g424 ( 
.A(n_355),
.B(n_357),
.Y(n_424)
);

NAND2x1p5_ASAP7_75t_L g425 ( 
.A(n_350),
.B(n_39),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_319),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_327),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_365),
.B(n_41),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_366),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_354),
.B(n_46),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_356),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_349),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_354),
.B(n_369),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_358),
.B(n_47),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_364),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_355),
.B(n_48),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_335),
.B(n_50),
.Y(n_439)
);

O2A1O1Ixp5_ASAP7_75t_L g440 ( 
.A1(n_381),
.A2(n_307),
.B(n_363),
.C(n_354),
.Y(n_440)
);

NAND3xp33_ASAP7_75t_SL g441 ( 
.A(n_387),
.B(n_407),
.C(n_423),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_388),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_373),
.Y(n_443)
);

AOI21x1_ASAP7_75t_L g444 ( 
.A1(n_434),
.A2(n_51),
.B(n_52),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_372),
.A2(n_357),
.B(n_360),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_383),
.B(n_360),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_435),
.A2(n_53),
.B(n_54),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_400),
.B(n_411),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_55),
.Y(n_449)
);

AO21x2_ASAP7_75t_L g450 ( 
.A1(n_377),
.A2(n_157),
.B(n_61),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_60),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_379),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_414),
.B(n_62),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_402),
.B(n_63),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_424),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_404),
.Y(n_456)
);

NAND2x1p5_ASAP7_75t_L g457 ( 
.A(n_412),
.B(n_64),
.Y(n_457)
);

O2A1O1Ixp33_ASAP7_75t_L g458 ( 
.A1(n_396),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_458)
);

OA21x2_ASAP7_75t_L g459 ( 
.A1(n_382),
.A2(n_68),
.B(n_70),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_395),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_71),
.Y(n_461)
);

O2A1O1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_391),
.A2(n_73),
.B(n_75),
.C(n_77),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_380),
.A2(n_421),
.B(n_415),
.Y(n_463)
);

OAI21xp33_ASAP7_75t_SL g464 ( 
.A1(n_403),
.A2(n_81),
.B(n_82),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_405),
.Y(n_465)
);

O2A1O1Ixp33_ASAP7_75t_SL g466 ( 
.A1(n_419),
.A2(n_83),
.B(n_87),
.C(n_89),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_384),
.B(n_90),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_412),
.B(n_91),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_410),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_401),
.B(n_93),
.Y(n_470)
);

AO22x2_ASAP7_75t_L g471 ( 
.A1(n_439),
.A2(n_438),
.B1(n_376),
.B2(n_385),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_437),
.B(n_95),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_413),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_416),
.B(n_97),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_431),
.A2(n_98),
.B(n_99),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_100),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

NOR3xp33_ASAP7_75t_SL g478 ( 
.A(n_430),
.B(n_105),
.C(n_106),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_432),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_406),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_392),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_416),
.B(n_113),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_394),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_418),
.Y(n_484)
);

OR2x6_ASAP7_75t_L g485 ( 
.A(n_424),
.B(n_425),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_422),
.A2(n_117),
.B(n_119),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_422),
.Y(n_487)
);

AOI21x1_ASAP7_75t_L g488 ( 
.A1(n_417),
.A2(n_120),
.B(n_121),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_428),
.B(n_123),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_386),
.B(n_124),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_SL g491 ( 
.A1(n_397),
.A2(n_389),
.B(n_390),
.C(n_409),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_439),
.Y(n_492)
);

A2O1A1Ixp33_ASAP7_75t_L g493 ( 
.A1(n_371),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_420),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_374),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_422),
.A2(n_132),
.B(n_133),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_375),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_460),
.Y(n_498)
);

AO21x2_ASAP7_75t_L g499 ( 
.A1(n_448),
.A2(n_393),
.B(n_398),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_456),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_452),
.B(n_394),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_457),
.Y(n_502)
);

AO21x2_ASAP7_75t_L g503 ( 
.A1(n_489),
.A2(n_399),
.B(n_427),
.Y(n_503)
);

AO21x2_ASAP7_75t_L g504 ( 
.A1(n_454),
.A2(n_426),
.B(n_394),
.Y(n_504)
);

AO21x2_ASAP7_75t_L g505 ( 
.A1(n_491),
.A2(n_394),
.B(n_436),
.Y(n_505)
);

AO21x2_ASAP7_75t_L g506 ( 
.A1(n_450),
.A2(n_441),
.B(n_463),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_446),
.B(n_436),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_444),
.A2(n_436),
.B(n_135),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_465),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_477),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_469),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_492),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_488),
.A2(n_436),
.B(n_138),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_459),
.Y(n_514)
);

BUFx4f_ASAP7_75t_SL g515 ( 
.A(n_481),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_484),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_457),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_473),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_455),
.B(n_378),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_470),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_440),
.A2(n_134),
.B(n_139),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_442),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_443),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_497),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_484),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_495),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_479),
.B(n_141),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_450),
.A2(n_143),
.B(n_144),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_483),
.B(n_145),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_459),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_453),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_468),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_474),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_482),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_449),
.Y(n_535)
);

BUFx2_ASAP7_75t_SL g536 ( 
.A(n_461),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_471),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_483),
.B(n_146),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_485),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_487),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_485),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_485),
.B(n_150),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_447),
.A2(n_151),
.B(n_153),
.Y(n_543)
);

BUFx8_ASAP7_75t_L g544 ( 
.A(n_471),
.Y(n_544)
);

CKINVDCx11_ASAP7_75t_R g545 ( 
.A(n_541),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_529),
.A2(n_480),
.B1(n_464),
.B2(n_451),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_529),
.A2(n_490),
.B1(n_476),
.B2(n_494),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_500),
.B(n_445),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_507),
.A2(n_467),
.B(n_462),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_509),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_522),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_526),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_523),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_510),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_521),
.A2(n_475),
.B(n_496),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_498),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_498),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_512),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_539),
.Y(n_559)
);

INVx6_ASAP7_75t_L g560 ( 
.A(n_517),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_523),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_524),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_525),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_521),
.A2(n_486),
.B(n_458),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_541),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_511),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_532),
.A2(n_478),
.B1(n_472),
.B2(n_493),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_539),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_542),
.B(n_155),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_515),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_538),
.A2(n_156),
.B1(n_466),
.B2(n_520),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_532),
.A2(n_531),
.B(n_527),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_514),
.A2(n_508),
.B(n_530),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_542),
.B(n_538),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_518),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_542),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_517),
.Y(n_577)
);

AO21x2_ASAP7_75t_L g578 ( 
.A1(n_506),
.A2(n_530),
.B(n_505),
.Y(n_578)
);

CKINVDCx11_ASAP7_75t_R g579 ( 
.A(n_517),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_L g580 ( 
.A1(n_501),
.A2(n_537),
.B1(n_502),
.B2(n_517),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_502),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_537),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_544),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_529),
.A2(n_544),
.B1(n_531),
.B2(n_535),
.Y(n_584)
);

NAND2x1p5_ASAP7_75t_L g585 ( 
.A(n_516),
.B(n_502),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_502),
.Y(n_586)
);

BUFx8_ASAP7_75t_L g587 ( 
.A(n_502),
.Y(n_587)
);

INVxp33_ASAP7_75t_SL g588 ( 
.A(n_570),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_556),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_576),
.B(n_525),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_556),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_546),
.B(n_544),
.C(n_535),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_572),
.B(n_529),
.Y(n_593)
);

INVx8_ASAP7_75t_L g594 ( 
.A(n_574),
.Y(n_594)
);

INVxp33_ASAP7_75t_SL g595 ( 
.A(n_545),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_550),
.Y(n_596)
);

BUFx4f_ASAP7_75t_SL g597 ( 
.A(n_559),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_557),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_554),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_547),
.A2(n_499),
.B(n_503),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_545),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_565),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_547),
.A2(n_529),
.B1(n_533),
.B2(n_534),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_551),
.Y(n_604)
);

A2O1A1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_549),
.A2(n_543),
.B(n_535),
.C(n_534),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_R g606 ( 
.A(n_576),
.B(n_519),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_569),
.B(n_540),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_574),
.B(n_533),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_548),
.B(n_529),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_582),
.B(n_535),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_569),
.B(n_535),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_568),
.B(n_534),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_R g613 ( 
.A(n_579),
.B(n_534),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_574),
.B(n_534),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_580),
.B(n_533),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_579),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_557),
.B(n_533),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_552),
.Y(n_618)
);

NAND3xp33_ASAP7_75t_L g619 ( 
.A(n_584),
.B(n_567),
.C(n_571),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_558),
.B(n_566),
.Y(n_620)
);

INVxp33_ASAP7_75t_L g621 ( 
.A(n_558),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_559),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_560),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_575),
.Y(n_624)
);

INVxp33_ASAP7_75t_L g625 ( 
.A(n_583),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_584),
.A2(n_516),
.B1(n_533),
.B2(n_536),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_587),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_562),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_580),
.B(n_499),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_587),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_564),
.A2(n_543),
.B(n_513),
.C(n_508),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_577),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_596),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_609),
.B(n_578),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_598),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_619),
.A2(n_571),
.B1(n_503),
.B2(n_504),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_604),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_608),
.B(n_586),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_610),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_628),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_608),
.B(n_586),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_617),
.B(n_578),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_620),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_618),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_629),
.B(n_506),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_629),
.B(n_506),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_624),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_610),
.B(n_563),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_593),
.B(n_553),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_621),
.B(n_561),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_592),
.A2(n_503),
.B1(n_504),
.B2(n_505),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_593),
.B(n_561),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_615),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_608),
.B(n_581),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_615),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_614),
.B(n_528),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_603),
.B(n_581),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_611),
.B(n_607),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_614),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_632),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_591),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_594),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_612),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_589),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_590),
.B(n_577),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_594),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_626),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_605),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_642),
.B(n_600),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_663),
.B(n_626),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_633),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_664),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_643),
.B(n_639),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_640),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_659),
.B(n_602),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_637),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_644),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_647),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_642),
.B(n_528),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_635),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_640),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_659),
.B(n_528),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_634),
.B(n_594),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_663),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_634),
.B(n_573),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_656),
.B(n_505),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_656),
.B(n_625),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_649),
.B(n_631),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_668),
.A2(n_595),
.B1(n_588),
.B2(n_601),
.Y(n_689)
);

INVxp67_ASAP7_75t_SL g690 ( 
.A(n_667),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_660),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_SL g692 ( 
.A(n_668),
.B(n_613),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_653),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_653),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_655),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_645),
.B(n_622),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_669),
.B(n_646),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_669),
.B(n_646),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_691),
.B(n_661),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_672),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_680),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_673),
.B(n_655),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_674),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_687),
.B(n_652),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_671),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_688),
.B(n_645),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_688),
.B(n_657),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_696),
.B(n_648),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_679),
.B(n_657),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_696),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_670),
.A2(n_692),
.B(n_636),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_691),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_676),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_677),
.B(n_648),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_705),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_700),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_713),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_711),
.A2(n_670),
.B1(n_692),
.B2(n_665),
.Y(n_718)
);

OAI21xp33_ASAP7_75t_L g719 ( 
.A1(n_707),
.A2(n_690),
.B(n_683),
.Y(n_719)
);

AOI32xp33_ASAP7_75t_L g720 ( 
.A1(n_707),
.A2(n_684),
.A3(n_689),
.B1(n_679),
.B2(n_682),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_703),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_710),
.B(n_685),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_703),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_701),
.B(n_685),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_718),
.A2(n_684),
.B1(n_700),
.B2(n_704),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_718),
.B(n_702),
.C(n_684),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_719),
.A2(n_662),
.B1(n_666),
.B2(n_706),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_715),
.A2(n_717),
.B(n_724),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_723),
.Y(n_729)
);

OAI21xp33_ASAP7_75t_L g730 ( 
.A1(n_726),
.A2(n_720),
.B(n_722),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_727),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_725),
.A2(n_716),
.B1(n_675),
.B2(n_708),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_729),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_733),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_732),
.B(n_730),
.Y(n_735)
);

AOI221xp5_ASAP7_75t_L g736 ( 
.A1(n_731),
.A2(n_728),
.B1(n_699),
.B2(n_714),
.C(n_712),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_731),
.B(n_699),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_734),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_735),
.B(n_699),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_R g740 ( 
.A(n_738),
.B(n_616),
.Y(n_740)
);

OAI221xp5_ASAP7_75t_L g741 ( 
.A1(n_739),
.A2(n_736),
.B1(n_737),
.B2(n_712),
.C(n_627),
.Y(n_741)
);

AOI321xp33_ASAP7_75t_L g742 ( 
.A1(n_738),
.A2(n_658),
.A3(n_665),
.B1(n_651),
.B2(n_682),
.C(n_686),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_741),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_740),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_742),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_741),
.A2(n_630),
.B1(n_597),
.B2(n_706),
.Y(n_746)
);

NOR2x1_ASAP7_75t_L g747 ( 
.A(n_741),
.B(n_606),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_740),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_744),
.Y(n_749)
);

AND3x2_ASAP7_75t_L g750 ( 
.A(n_743),
.B(n_599),
.C(n_666),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_748),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_745),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_747),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_746),
.B(n_709),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_744),
.B(n_709),
.Y(n_755)
);

CKINVDCx16_ASAP7_75t_R g756 ( 
.A(n_751),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_R g757 ( 
.A(n_749),
.B(n_599),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_752),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_753),
.B(n_721),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_755),
.Y(n_760)
);

NOR2x1_ASAP7_75t_L g761 ( 
.A(n_752),
.B(n_678),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_760),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_756),
.Y(n_763)
);

XNOR2x2_ASAP7_75t_L g764 ( 
.A(n_761),
.B(n_750),
.Y(n_764)
);

NAND4xp25_ASAP7_75t_L g765 ( 
.A(n_758),
.B(n_754),
.C(n_650),
.D(n_662),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_759),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_757),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_760),
.Y(n_768)
);

NAND4xp25_ASAP7_75t_L g769 ( 
.A(n_758),
.B(n_698),
.C(n_697),
.D(n_638),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_763),
.A2(n_762),
.B1(n_768),
.B2(n_767),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_766),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_764),
.Y(n_772)
);

OAI31xp33_ASAP7_75t_L g773 ( 
.A1(n_765),
.A2(n_585),
.A3(n_623),
.B(n_638),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_769),
.A2(n_654),
.B1(n_641),
.B2(n_638),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_763),
.A2(n_654),
.B1(n_641),
.B2(n_560),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_763),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_763),
.A2(n_654),
.B1(n_641),
.B2(n_560),
.Y(n_777)
);

OAI22x1_ASAP7_75t_L g778 ( 
.A1(n_770),
.A2(n_585),
.B1(n_697),
.B2(n_698),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_776),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_772),
.A2(n_513),
.B(n_555),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_771),
.Y(n_781)
);

OAI22xp33_ASAP7_75t_L g782 ( 
.A1(n_775),
.A2(n_693),
.B1(n_695),
.B2(n_694),
.Y(n_782)
);

OA22x2_ASAP7_75t_L g783 ( 
.A1(n_779),
.A2(n_777),
.B1(n_774),
.B2(n_773),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_781),
.Y(n_784)
);

XNOR2xp5_ASAP7_75t_L g785 ( 
.A(n_783),
.B(n_778),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_785),
.A2(n_784),
.B1(n_782),
.B2(n_780),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_786),
.B(n_681),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_787),
.A2(n_681),
.B1(n_674),
.B2(n_499),
.Y(n_788)
);


endmodule