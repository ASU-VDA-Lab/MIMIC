module real_aes_2550_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_792;
wire n_503;
wire n_673;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_976;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_884;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_961;
wire n_870;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_1078;
wire n_744;
wire n_938;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_559;
wire n_1049;
wire n_466;
wire n_636;
wire n_1053;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_1070;
wire n_726;
wire n_517;
wire n_931;
wire n_683;
wire n_904;
wire n_780;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_529;
wire n_725;
wire n_973;
wire n_455;
wire n_504;
wire n_671;
wire n_960;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_936;
wire n_610;
wire n_581;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_676;
wire n_658;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_853;
wire n_1079;
wire n_843;
wire n_810;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_649;
wire n_663;
wire n_1056;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_899;
wire n_637;
wire n_526;
wire n_653;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_1055;
wire n_988;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_1040;
wire n_703;
wire n_652;
wire n_500;
wire n_1101;
wire n_1102;
wire n_601;
wire n_463;
wire n_661;
wire n_804;
wire n_1076;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
wire n_429;
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_0), .A2(n_246), .B1(n_729), .B2(n_730), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_1), .A2(n_322), .B1(n_446), .B2(n_632), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_2), .A2(n_73), .B1(n_513), .B2(n_650), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_3), .A2(n_128), .B1(n_627), .B2(n_696), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_4), .A2(n_140), .B1(n_822), .B2(n_823), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_5), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_6), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_7), .A2(n_265), .B1(n_483), .B2(n_591), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g933 ( .A1(n_8), .A2(n_83), .B1(n_510), .B2(n_934), .Y(n_933) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_9), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_10), .Y(n_887) );
AOI22xp33_ASAP7_75t_SL g815 ( .A1(n_11), .A2(n_359), .B1(n_816), .B2(n_817), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_12), .A2(n_71), .B1(n_627), .B2(n_628), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_13), .A2(n_392), .B1(n_494), .B2(n_497), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_14), .A2(n_219), .B1(n_722), .B2(n_723), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_15), .A2(n_267), .B1(n_670), .B2(n_1000), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_16), .A2(n_270), .B1(n_512), .B2(n_513), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_17), .A2(n_315), .B1(n_617), .B2(n_619), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_18), .A2(n_330), .B1(n_480), .B2(n_678), .Y(n_1025) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_19), .A2(n_91), .B1(n_936), .B2(n_937), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_20), .A2(n_149), .B1(n_513), .B2(n_650), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_21), .A2(n_198), .B1(n_484), .B2(n_591), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_22), .A2(n_344), .B1(n_544), .B2(n_545), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_23), .A2(n_204), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_24), .A2(n_110), .B1(n_678), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_25), .A2(n_308), .B1(n_718), .B2(n_719), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_26), .A2(n_295), .B1(n_676), .B2(n_921), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_27), .A2(n_158), .B1(n_495), .B2(n_750), .Y(n_955) );
INVx1_ASAP7_75t_SL g426 ( .A(n_28), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g1045 ( .A(n_28), .B(n_48), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_29), .A2(n_130), .B1(n_550), .B2(n_584), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_30), .A2(n_283), .B1(n_715), .B2(n_1005), .Y(n_1004) );
AOI22xp5_ASAP7_75t_SL g1029 ( .A1(n_31), .A2(n_272), .B1(n_670), .B2(n_790), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_32), .A2(n_355), .B1(n_477), .B2(n_618), .Y(n_1094) );
AOI222xp33_ASAP7_75t_L g751 ( .A1(n_33), .A2(n_326), .B1(n_364), .B2(n_599), .C1(n_752), .C2(n_753), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_34), .B(n_580), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g982 ( .A(n_35), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_36), .A2(n_42), .B1(n_678), .B2(n_722), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g1055 ( .A(n_37), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_38), .A2(n_233), .B1(n_783), .B2(n_784), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_39), .A2(n_312), .B1(n_696), .B2(n_748), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_40), .A2(n_255), .B1(n_622), .B2(n_624), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_41), .A2(n_230), .B1(n_873), .B2(n_1098), .Y(n_1097) );
XNOR2x1_ASAP7_75t_SL g925 ( .A(n_43), .B(n_926), .Y(n_925) );
AOI22xp5_ASAP7_75t_SL g963 ( .A1(n_43), .A2(n_926), .B1(n_964), .B2(n_965), .Y(n_963) );
INVx1_ASAP7_75t_L g965 ( .A(n_43), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_44), .A2(n_276), .B1(n_637), .B2(n_638), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_45), .A2(n_120), .B1(n_498), .B2(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_46), .A2(n_113), .B1(n_743), .B2(n_826), .Y(n_825) );
OA21x2_ASAP7_75t_L g413 ( .A1(n_47), .A2(n_414), .B(n_502), .Y(n_413) );
INVx1_ASAP7_75t_L g504 ( .A(n_47), .Y(n_504) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_48), .A2(n_370), .B1(n_425), .B2(n_429), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g1063 ( .A(n_49), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_50), .A2(n_307), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_51), .A2(n_121), .B1(n_624), .B2(n_961), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_52), .A2(n_203), .B1(n_622), .B2(n_623), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_53), .A2(n_106), .B1(n_555), .B2(n_556), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_54), .A2(n_291), .B1(n_682), .B2(n_737), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_55), .A2(n_126), .B1(n_727), .B2(n_946), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_56), .A2(n_294), .B1(n_952), .B2(n_953), .Y(n_951) );
INVx1_ASAP7_75t_L g427 ( .A(n_57), .Y(n_427) );
AO222x2_ASAP7_75t_SL g647 ( .A1(n_58), .A2(n_220), .B1(n_300), .B2(n_543), .C1(n_544), .C2(n_545), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_59), .A2(n_360), .B1(n_439), .B2(n_516), .Y(n_811) );
INVx1_ASAP7_75t_L g1018 ( .A(n_60), .Y(n_1018) );
AOI222xp33_ASAP7_75t_L g1010 ( .A1(n_61), .A2(n_205), .B1(n_354), .B2(n_597), .C1(n_915), .C2(n_1011), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_62), .A2(n_286), .B1(n_699), .B2(n_700), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_63), .B(n_795), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_64), .A2(n_132), .B1(n_936), .B2(n_937), .Y(n_1006) );
AOI22xp33_ASAP7_75t_SL g605 ( .A1(n_65), .A2(n_336), .B1(n_555), .B2(n_556), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_66), .A2(n_133), .B1(n_489), .B2(n_873), .Y(n_872) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_67), .A2(n_399), .B1(n_409), .B2(n_1046), .C(n_1047), .Y(n_398) );
AO222x2_ASAP7_75t_SL g542 ( .A1(n_68), .A2(n_137), .B1(n_181), .B2(n_543), .C1(n_544), .C2(n_545), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_69), .A2(n_153), .B1(n_444), .B2(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_70), .A2(n_310), .B1(n_510), .B2(n_715), .Y(n_916) );
AO22x2_ASAP7_75t_L g435 ( .A1(n_72), .A2(n_212), .B1(n_425), .B2(n_436), .Y(n_435) );
XNOR2x1_ASAP7_75t_L g661 ( .A(n_74), .B(n_662), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_75), .A2(n_79), .B1(n_524), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_76), .A2(n_337), .B1(n_723), .B2(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_77), .A2(n_368), .B1(n_699), .B2(n_700), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_78), .A2(n_177), .B1(n_531), .B2(n_532), .Y(n_530) );
AOI221x1_ASAP7_75t_L g677 ( .A1(n_80), .A2(n_90), .B1(n_534), .B2(n_678), .C(n_679), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_81), .A2(n_293), .B1(n_512), .B2(n_513), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_82), .A2(n_170), .B1(n_727), .B2(n_1092), .Y(n_1091) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_84), .A2(n_347), .B1(n_510), .B2(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_85), .A2(n_141), .B1(n_618), .B2(n_619), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_86), .A2(n_178), .B1(n_618), .B2(n_737), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_87), .A2(n_342), .B1(n_524), .B2(n_559), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_88), .A2(n_211), .B1(n_696), .B2(n_748), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_89), .A2(n_277), .B1(n_470), .B2(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_92), .B(n_752), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_93), .A2(n_1049), .B1(n_1079), .B2(n_1080), .Y(n_1048) );
CKINVDCx20_ASAP7_75t_R g1080 ( .A(n_93), .Y(n_1080) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_94), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_95), .A2(n_264), .B1(n_670), .B2(n_727), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_96), .A2(n_289), .B1(n_524), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_97), .A2(n_297), .B1(n_619), .B2(n_1002), .Y(n_1001) );
AO22x1_ASAP7_75t_L g437 ( .A1(n_98), .A2(n_266), .B1(n_438), .B2(n_444), .Y(n_437) );
INVx1_ASAP7_75t_L g683 ( .A(n_99), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_100), .A2(n_396), .B1(n_531), .B2(n_532), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g898 ( .A1(n_101), .A2(n_127), .B1(n_484), .B2(n_743), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_102), .A2(n_273), .B1(n_559), .B2(n_591), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_103), .A2(n_215), .B1(n_817), .B2(n_873), .Y(n_891) );
AOI22xp33_ASAP7_75t_SL g930 ( .A1(n_104), .A2(n_314), .B1(n_446), .B2(n_931), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_105), .B(n_635), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g990 ( .A1(n_107), .A2(n_151), .B1(n_471), .B2(n_591), .Y(n_990) );
INVx1_ASAP7_75t_L g691 ( .A(n_108), .Y(n_691) );
INVx1_ASAP7_75t_L g668 ( .A(n_109), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_111), .A2(n_251), .B1(n_722), .B2(n_723), .Y(n_1009) );
AO22x2_ASAP7_75t_L g860 ( .A1(n_112), .A2(n_861), .B1(n_879), .B2(n_880), .Y(n_860) );
INVx1_ASAP7_75t_L g880 ( .A(n_112), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_114), .A2(n_258), .B1(n_558), .B2(n_562), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_115), .A2(n_346), .B1(n_548), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_116), .A2(n_373), .B1(n_439), .B2(n_516), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_117), .A2(n_385), .B1(n_438), .B2(n_1011), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_118), .A2(n_313), .B1(n_458), .B2(n_829), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_119), .A2(n_348), .B1(n_524), .B2(n_559), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_122), .A2(n_157), .B1(n_498), .B2(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_123), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_124), .A2(n_268), .B1(n_670), .B2(n_727), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g1030 ( .A1(n_125), .A2(n_284), .B1(n_627), .B2(n_719), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_129), .A2(n_199), .B1(n_678), .B2(n_941), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_131), .A2(n_339), .B1(n_476), .B2(n_725), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_134), .A2(n_351), .B1(n_729), .B2(n_730), .Y(n_1008) );
AO22x2_ASAP7_75t_L g432 ( .A1(n_135), .A2(n_298), .B1(n_425), .B2(n_433), .Y(n_432) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_136), .A2(n_242), .B1(n_512), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_138), .A2(n_350), .B1(n_723), .B2(n_790), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_139), .A2(n_166), .B1(n_458), .B2(n_534), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_142), .A2(n_365), .B1(n_558), .B2(n_559), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_143), .A2(n_192), .B1(n_544), .B2(n_545), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_144), .A2(n_282), .B1(n_619), .B2(n_786), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_145), .A2(n_175), .B1(n_817), .B2(n_873), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_146), .A2(n_184), .B1(n_550), .B2(n_551), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_147), .A2(n_363), .B1(n_480), .B2(n_483), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_148), .A2(n_164), .B1(n_723), .B2(n_727), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_150), .A2(n_250), .B1(n_465), .B2(n_468), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_152), .B(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_154), .A2(n_226), .B1(n_550), .B2(n_584), .Y(n_765) );
INVx1_ASAP7_75t_L g802 ( .A(n_155), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_156), .A2(n_168), .B1(n_438), .B2(n_798), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_159), .A2(n_245), .B1(n_826), .B2(n_941), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_160), .A2(n_328), .B1(n_544), .B2(n_599), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_161), .A2(n_311), .B1(n_532), .B2(n_589), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g1065 ( .A(n_162), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_163), .A2(n_380), .B1(n_498), .B2(n_814), .Y(n_874) );
XOR2x2_ASAP7_75t_L g883 ( .A(n_165), .B(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_167), .A2(n_329), .B1(n_531), .B2(n_532), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g980 ( .A(n_169), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_171), .Y(n_659) );
AO22x1_ASAP7_75t_L g840 ( .A1(n_172), .A2(n_237), .B1(n_446), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_173), .A2(n_188), .B1(n_718), .B2(n_719), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_174), .B(n_597), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g1061 ( .A(n_176), .Y(n_1061) );
AOI22xp33_ASAP7_75t_SL g601 ( .A1(n_179), .A2(n_372), .B1(n_550), .B2(n_551), .Y(n_601) );
OA22x2_ASAP7_75t_L g506 ( .A1(n_180), .A2(n_507), .B1(n_536), .B2(n_537), .Y(n_506) );
INVx1_ASAP7_75t_L g536 ( .A(n_180), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_182), .A2(n_305), .B1(n_826), .B2(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g667 ( .A(n_183), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_185), .A2(n_218), .B1(n_699), .B2(n_700), .Y(n_1078) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_186), .A2(n_259), .B1(n_525), .B2(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_187), .A2(n_229), .B1(n_666), .B2(n_823), .Y(n_878) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_189), .A2(n_299), .B1(n_739), .B2(n_740), .Y(n_738) );
XNOR2x1_ASAP7_75t_L g707 ( .A(n_190), .B(n_708), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g1069 ( .A(n_191), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_193), .B(n_444), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_194), .B(n_597), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_195), .A2(n_234), .B1(n_555), .B2(n_556), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g986 ( .A(n_196), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_197), .A2(n_262), .B1(n_458), .B2(n_739), .Y(n_958) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_200), .B(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_201), .A2(n_249), .B1(n_722), .B2(n_729), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_202), .A2(n_280), .B1(n_510), .B2(n_934), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_206), .A2(n_341), .B1(n_522), .B2(n_525), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_207), .A2(n_303), .B1(n_515), .B2(n_516), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_208), .A2(n_387), .B1(n_555), .B2(n_556), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_209), .A2(n_285), .B1(n_470), .B2(n_524), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_210), .A2(n_260), .B1(n_666), .B2(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1044 ( .A(n_212), .Y(n_1044) );
INVx1_ASAP7_75t_L g673 ( .A(n_213), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_214), .A2(n_274), .B1(n_730), .B2(n_740), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_216), .A2(n_376), .B1(n_532), .B2(n_589), .Y(n_993) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_217), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_221), .A2(n_389), .B1(n_788), .B2(n_853), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_222), .A2(n_320), .B1(n_556), .B2(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_223), .A2(n_390), .B1(n_786), .B2(n_788), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g820 ( .A1(n_224), .A2(n_382), .B1(n_476), .B2(n_787), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_225), .A2(n_261), .B1(n_531), .B2(n_532), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_227), .A2(n_393), .B1(n_624), .B2(n_829), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g1072 ( .A(n_228), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_231), .A2(n_391), .B1(n_544), .B2(n_545), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g1059 ( .A(n_232), .Y(n_1059) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_235), .A2(n_256), .B1(n_446), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_236), .A2(n_397), .B1(n_618), .B2(n_737), .Y(n_959) );
INVx2_ASAP7_75t_L g408 ( .A(n_238), .Y(n_408) );
XOR2x2_ASAP7_75t_L g909 ( .A(n_239), .B(n_910), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_240), .A2(n_253), .B1(n_480), .B2(n_483), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g1053 ( .A(n_241), .Y(n_1053) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_243), .Y(n_1068) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_244), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_247), .A2(n_269), .B1(n_524), .B2(n_559), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_248), .A2(n_357), .B1(n_495), .B2(n_750), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_252), .A2(n_334), .B1(n_452), .B2(n_458), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_254), .A2(n_321), .B1(n_531), .B2(n_532), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_257), .A2(n_343), .B1(n_512), .B2(n_548), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g929 ( .A(n_263), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_271), .A2(n_278), .B1(n_476), .B2(n_725), .Y(n_942) );
XOR2x2_ASAP7_75t_L g996 ( .A(n_275), .B(n_997), .Y(n_996) );
AO22x2_ASAP7_75t_L g1087 ( .A1(n_279), .A2(n_1088), .B1(n_1101), .B2(n_1102), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_279), .Y(n_1101) );
INVx1_ASAP7_75t_L g672 ( .A(n_281), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_287), .A2(n_335), .B1(n_798), .B2(n_915), .Y(n_914) );
OA22x2_ASAP7_75t_L g732 ( .A1(n_288), .A2(n_733), .B1(n_734), .B2(n_755), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_288), .Y(n_733) );
AO21x2_ASAP7_75t_L g758 ( .A1(n_288), .A2(n_734), .B(n_759), .Y(n_758) );
AOI22x1_ASAP7_75t_L g539 ( .A1(n_290), .A2(n_540), .B1(n_564), .B2(n_565), .Y(n_539) );
INVx1_ASAP7_75t_L g565 ( .A(n_290), .Y(n_565) );
XNOR2x1_ASAP7_75t_L g948 ( .A(n_292), .B(n_949), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_296), .B(n_1022), .Y(n_1021) );
NOR2xp33_ASAP7_75t_L g1042 ( .A(n_298), .B(n_1043), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_301), .A2(n_366), .B1(n_516), .B2(n_931), .Y(n_1099) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_302), .A2(n_327), .B1(n_559), .B2(n_591), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_304), .B(n_519), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_306), .A2(n_383), .B1(n_550), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_309), .A2(n_353), .B1(n_676), .B2(n_743), .Y(n_868) );
AND2x2_ASAP7_75t_L g839 ( .A(n_316), .B(n_795), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_317), .A2(n_332), .B1(n_476), .B2(n_528), .Y(n_527) );
OA22x2_ASAP7_75t_L g972 ( .A1(n_318), .A2(n_973), .B1(n_974), .B2(n_995), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_318), .Y(n_973) );
INVx3_ASAP7_75t_L g425 ( .A(n_319), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_323), .Y(n_1075) );
INVx1_ASAP7_75t_L g684 ( .A(n_324), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_325), .A2(n_338), .B1(n_487), .B2(n_489), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_331), .A2(n_384), .B1(n_748), .B2(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g834 ( .A(n_333), .Y(n_834) );
AND2x2_ASAP7_75t_L g417 ( .A(n_340), .B(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_345), .A2(n_379), .B1(n_676), .B2(n_877), .Y(n_1090) );
INVx1_ASAP7_75t_L g693 ( .A(n_349), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_352), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_356), .A2(n_362), .B1(n_1002), .B2(n_1027), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_358), .A2(n_361), .B1(n_473), .B2(n_476), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_367), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_369), .B(n_580), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_371), .A2(n_378), .B1(n_699), .B2(n_1024), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_374), .B(n_635), .Y(n_913) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_375), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g1040 ( .A(n_375), .Y(n_1040) );
INVx1_ASAP7_75t_L g405 ( .A(n_377), .Y(n_405) );
AND2x2_ASAP7_75t_R g1082 ( .A(n_377), .B(n_1040), .Y(n_1082) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_381), .B(n_407), .Y(n_406) );
XNOR2xp5_ASAP7_75t_L g612 ( .A(n_386), .B(n_613), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_388), .Y(n_849) );
INVx1_ASAP7_75t_L g688 ( .A(n_394), .Y(n_688) );
XOR2x2_ASAP7_75t_L g805 ( .A(n_395), .B(n_806), .Y(n_805) );
CKINVDCx6p67_ASAP7_75t_R g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_SL g402 ( .A(n_403), .B(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_404), .B(n_406), .Y(n_1105) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_405), .B(n_1040), .Y(n_1039) );
AOI21xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_904), .B(n_1037), .Y(n_409) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_410), .B(n_904), .Y(n_1046) );
XOR2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_703), .Y(n_410) );
XNOR2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_570), .Y(n_411) );
AO22x2_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_505), .B1(n_568), .B2(n_569), .Y(n_412) );
INVx1_ASAP7_75t_L g568 ( .A(n_413), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_414), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_485), .Y(n_415) );
NOR3xp33_ASAP7_75t_SL g416 ( .A(n_417), .B(n_437), .C(n_450), .Y(n_416) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_SL g519 ( .A(n_420), .Y(n_519) );
INVx4_ASAP7_75t_SL g580 ( .A(n_420), .Y(n_580) );
INVx4_ASAP7_75t_SL g597 ( .A(n_420), .Y(n_597) );
BUFx2_ASAP7_75t_L g796 ( .A(n_420), .Y(n_796) );
INVx3_ASAP7_75t_L g1022 ( .A(n_420), .Y(n_1022) );
INVx6_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_430), .Y(n_421) );
AND2x4_ASAP7_75t_L g491 ( .A(n_422), .B(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g499 ( .A(n_422), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g513 ( .A(n_422), .B(n_492), .Y(n_513) );
AND2x4_ASAP7_75t_L g543 ( .A(n_422), .B(n_430), .Y(n_543) );
AND2x2_ASAP7_75t_L g548 ( .A(n_422), .B(n_492), .Y(n_548) );
AND2x2_ASAP7_75t_L g551 ( .A(n_422), .B(n_500), .Y(n_551) );
AND2x2_ASAP7_75t_L g584 ( .A(n_422), .B(n_500), .Y(n_584) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_428), .Y(n_422) );
AND2x2_ASAP7_75t_L g442 ( .A(n_423), .B(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_423), .Y(n_449) );
INVx2_ASAP7_75t_L g457 ( .A(n_423), .Y(n_457) );
OAI22x1_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_425), .Y(n_429) );
INVx2_ASAP7_75t_L g433 ( .A(n_425), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_425), .Y(n_436) );
INVx2_ASAP7_75t_L g443 ( .A(n_428), .Y(n_443) );
AND2x2_ASAP7_75t_L g456 ( .A(n_428), .B(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g478 ( .A(n_428), .Y(n_478) );
AND2x2_ASAP7_75t_L g455 ( .A(n_430), .B(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g467 ( .A(n_430), .B(n_461), .Y(n_467) );
AND2x4_ASAP7_75t_L g482 ( .A(n_430), .B(n_442), .Y(n_482) );
AND2x6_ASAP7_75t_L g524 ( .A(n_430), .B(n_456), .Y(n_524) );
AND2x2_ASAP7_75t_L g531 ( .A(n_430), .B(n_442), .Y(n_531) );
AND2x2_ASAP7_75t_L g558 ( .A(n_430), .B(n_461), .Y(n_558) );
AND2x2_ASAP7_75t_L g589 ( .A(n_430), .B(n_442), .Y(n_589) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g441 ( .A(n_432), .B(n_434), .Y(n_441) );
AND2x2_ASAP7_75t_L g448 ( .A(n_432), .B(n_435), .Y(n_448) );
INVx1_ASAP7_75t_L g463 ( .A(n_432), .Y(n_463) );
INVxp67_ASAP7_75t_L g492 ( .A(n_434), .Y(n_492) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g462 ( .A(n_435), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g1054 ( .A(n_438), .Y(n_1054) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g515 ( .A(n_440), .Y(n_515) );
INVx2_ASAP7_75t_L g633 ( .A(n_440), .Y(n_633) );
BUFx5_ASAP7_75t_L g931 ( .A(n_440), .Y(n_931) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AND2x4_ASAP7_75t_L g471 ( .A(n_441), .B(n_461), .Y(n_471) );
AND2x4_ASAP7_75t_L g488 ( .A(n_441), .B(n_456), .Y(n_488) );
AND2x2_ASAP7_75t_L g512 ( .A(n_441), .B(n_456), .Y(n_512) );
AND2x4_ASAP7_75t_L g544 ( .A(n_441), .B(n_442), .Y(n_544) );
AND2x2_ASAP7_75t_L g562 ( .A(n_441), .B(n_461), .Y(n_562) );
AND2x2_ASAP7_75t_L g650 ( .A(n_441), .B(n_456), .Y(n_650) );
AND2x2_ASAP7_75t_L g496 ( .A(n_442), .B(n_462), .Y(n_496) );
AND2x4_ASAP7_75t_L g550 ( .A(n_442), .B(n_462), .Y(n_550) );
AND2x4_ASAP7_75t_L g461 ( .A(n_443), .B(n_457), .Y(n_461) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI222xp33_ASAP7_75t_L g687 ( .A1(n_445), .A2(n_688), .B1(n_689), .B2(n_691), .C1(n_692), .C2(n_693), .Y(n_687) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g1011 ( .A(n_446), .Y(n_1011) );
BUFx12f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g517 ( .A(n_447), .Y(n_517) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
AND2x4_ASAP7_75t_L g477 ( .A(n_448), .B(n_478), .Y(n_477) );
AND2x4_ASAP7_75t_L g484 ( .A(n_448), .B(n_461), .Y(n_484) );
AND2x4_ASAP7_75t_L g532 ( .A(n_448), .B(n_461), .Y(n_532) );
AND2x2_ASAP7_75t_SL g545 ( .A(n_448), .B(n_449), .Y(n_545) );
AND2x4_ASAP7_75t_L g556 ( .A(n_448), .B(n_478), .Y(n_556) );
AND2x2_ASAP7_75t_SL g599 ( .A(n_448), .B(n_449), .Y(n_599) );
NAND4xp25_ASAP7_75t_L g450 ( .A(n_451), .B(n_464), .C(n_472), .D(n_479), .Y(n_450) );
INVx1_ASAP7_75t_L g1064 ( .A(n_452), .Y(n_1064) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_SL g727 ( .A(n_454), .Y(n_727) );
INVx3_ASAP7_75t_L g739 ( .A(n_454), .Y(n_739) );
INVx2_ASAP7_75t_L g822 ( .A(n_454), .Y(n_822) );
INVx2_ASAP7_75t_SL g1000 ( .A(n_454), .Y(n_1000) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g622 ( .A(n_455), .Y(n_622) );
BUFx2_ASAP7_75t_L g666 ( .A(n_455), .Y(n_666) );
AND2x2_ASAP7_75t_L g475 ( .A(n_456), .B(n_462), .Y(n_475) );
AND2x2_ASAP7_75t_SL g555 ( .A(n_456), .B(n_462), .Y(n_555) );
AND2x2_ASAP7_75t_L g771 ( .A(n_456), .B(n_462), .Y(n_771) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_SL g535 ( .A(n_459), .Y(n_535) );
INVx2_ASAP7_75t_L g670 ( .A(n_459), .Y(n_670) );
INVx2_ASAP7_75t_L g740 ( .A(n_459), .Y(n_740) );
INVx2_ASAP7_75t_L g784 ( .A(n_459), .Y(n_784) );
INVx2_ASAP7_75t_L g823 ( .A(n_459), .Y(n_823) );
INVx2_ASAP7_75t_SL g946 ( .A(n_459), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_459), .A2(n_1063), .B1(n_1064), .B2(n_1065), .Y(n_1062) );
INVx1_ASAP7_75t_SL g1092 ( .A(n_459), .Y(n_1092) );
INVx8_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AND2x6_ASAP7_75t_L g559 ( .A(n_461), .B(n_462), .Y(n_559) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_463), .Y(n_501) );
INVx2_ASAP7_75t_L g731 ( .A(n_465), .Y(n_731) );
BUFx6f_ASAP7_75t_L g921 ( .A(n_465), .Y(n_921) );
INVx4_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_SL g534 ( .A(n_466), .Y(n_534) );
INVx3_ASAP7_75t_L g591 ( .A(n_466), .Y(n_591) );
INVx2_ASAP7_75t_L g790 ( .A(n_466), .Y(n_790) );
INVx2_ASAP7_75t_SL g829 ( .A(n_466), .Y(n_829) );
INVx2_ASAP7_75t_SL g877 ( .A(n_466), .Y(n_877) );
INVx8_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g1071 ( .A1(n_469), .A2(n_1072), .B1(n_1073), .B2(n_1075), .Y(n_1071) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_470), .Y(n_723) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g526 ( .A(n_471), .Y(n_526) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_471), .Y(n_624) );
BUFx3_ASAP7_75t_L g676 ( .A(n_471), .Y(n_676) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g529 ( .A(n_475), .Y(n_529) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_475), .Y(n_618) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g619 ( .A(n_477), .Y(n_619) );
INVx5_ASAP7_75t_SL g685 ( .A(n_477), .Y(n_685) );
BUFx3_ASAP7_75t_L g1027 ( .A(n_477), .Y(n_1027) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_481), .A2(n_672), .B1(n_673), .B2(n_674), .Y(n_671) );
INVx2_ASAP7_75t_L g722 ( .A(n_481), .Y(n_722) );
INVx1_ASAP7_75t_SL g792 ( .A(n_481), .Y(n_792) );
INVx2_ASAP7_75t_L g941 ( .A(n_481), .Y(n_941) );
INVx3_ASAP7_75t_L g961 ( .A(n_481), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_481), .A2(n_1068), .B1(n_1069), .B2(n_1070), .Y(n_1067) );
INVx6_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx3_ASAP7_75t_L g743 ( .A(n_482), .Y(n_743) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_SL g678 ( .A(n_484), .Y(n_678) );
BUFx2_ASAP7_75t_SL g729 ( .A(n_484), .Y(n_729) );
INVx2_ASAP7_75t_L g827 ( .A(n_484), .Y(n_827) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_493), .Y(n_485) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_488), .Y(n_637) );
BUFx2_ASAP7_75t_L g816 ( .A(n_488), .Y(n_816) );
BUFx3_ASAP7_75t_L g873 ( .A(n_488), .Y(n_873) );
INVx2_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g638 ( .A(n_490), .Y(n_638) );
INVx2_ASAP7_75t_L g700 ( .A(n_490), .Y(n_700) );
INVx2_ASAP7_75t_L g719 ( .A(n_490), .Y(n_719) );
INVx2_ASAP7_75t_L g817 ( .A(n_490), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_490), .A2(n_847), .B1(n_848), .B2(n_849), .Y(n_846) );
INVx2_ASAP7_75t_L g937 ( .A(n_490), .Y(n_937) );
INVx1_ASAP7_75t_L g1098 ( .A(n_490), .Y(n_1098) );
INVx6_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_496), .Y(n_510) );
INVx3_ASAP7_75t_L g749 ( .A(n_496), .Y(n_749) );
BUFx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
BUFx6f_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g629 ( .A(n_499), .Y(n_629) );
INVx1_ASAP7_75t_L g697 ( .A(n_499), .Y(n_697) );
BUFx3_ASAP7_75t_L g750 ( .A(n_499), .Y(n_750) );
BUFx4f_ASAP7_75t_L g934 ( .A(n_499), .Y(n_934) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g569 ( .A(n_505), .Y(n_569) );
AOI22x1_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_538), .B1(n_566), .B2(n_567), .Y(n_505) );
INVx2_ASAP7_75t_L g567 ( .A(n_506), .Y(n_567) );
INVx1_ASAP7_75t_L g537 ( .A(n_507), .Y(n_537) );
NOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_520), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .C(n_514), .D(n_518), .Y(n_508) );
BUFx6f_ASAP7_75t_SL g627 ( .A(n_510), .Y(n_627) );
INVx1_ASAP7_75t_L g981 ( .A(n_510), .Y(n_981) );
INVx1_ASAP7_75t_L g713 ( .A(n_515), .Y(n_713) );
BUFx6f_ASAP7_75t_SL g915 ( .A(n_515), .Y(n_915) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g799 ( .A(n_517), .Y(n_799) );
INVx2_ASAP7_75t_L g953 ( .A(n_517), .Y(n_953) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_519), .Y(n_690) );
INVx2_ASAP7_75t_L g864 ( .A(n_519), .Y(n_864) );
NAND4xp25_ASAP7_75t_L g520 ( .A(n_521), .B(n_527), .C(n_530), .D(n_533), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_525), .Y(n_1033) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g610 ( .A(n_526), .Y(n_610) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g682 ( .A(n_529), .Y(n_682) );
INVx1_ASAP7_75t_L g787 ( .A(n_529), .Y(n_787) );
INVx2_ASAP7_75t_SL g566 ( .A(n_538), .Y(n_566) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AO22x2_ASAP7_75t_L g642 ( .A1(n_539), .A2(n_643), .B1(n_644), .B2(n_660), .Y(n_642) );
INVx1_ASAP7_75t_L g660 ( .A(n_539), .Y(n_660) );
INVx1_ASAP7_75t_L g564 ( .A(n_540), .Y(n_564) );
NAND2x1_ASAP7_75t_SL g540 ( .A(n_541), .B(n_552), .Y(n_540) );
NOR2xp67_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
BUFx2_ASAP7_75t_L g752 ( .A(n_543), .Y(n_752) );
INVx1_ASAP7_75t_SL g754 ( .A(n_544), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
INVxp67_ASAP7_75t_L g987 ( .A(n_548), .Y(n_987) );
NOR2x1_ASAP7_75t_L g552 ( .A(n_553), .B(n_560), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B1(n_640), .B2(n_702), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OA22x2_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_612), .B2(n_639), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
XNOR2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_592), .Y(n_574) );
XNOR2x1_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR2x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_585), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .C(n_582), .D(n_583), .Y(n_578) );
INVx1_ASAP7_75t_SL g809 ( .A(n_580), .Y(n_809) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .C(n_588), .D(n_590), .Y(n_585) );
XOR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_611), .Y(n_592) );
NAND2x1_ASAP7_75t_L g593 ( .A(n_594), .B(n_603), .Y(n_593) );
NOR2x1_ASAP7_75t_L g594 ( .A(n_595), .B(n_600), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
BUFx2_ASAP7_75t_L g635 ( .A(n_597), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NOR2x1_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx2_ASAP7_75t_SL g639 ( .A(n_612), .Y(n_639) );
NOR2xp67_ASAP7_75t_L g613 ( .A(n_614), .B(n_625), .Y(n_613) );
NAND4xp25_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .C(n_620), .D(n_621), .Y(n_614) );
INVx1_ASAP7_75t_L g1060 ( .A(n_617), .Y(n_1060) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND4xp25_ASAP7_75t_L g625 ( .A(n_626), .B(n_630), .C(n_634), .D(n_636), .Y(n_625) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g716 ( .A(n_629), .Y(n_716) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g692 ( .A(n_632), .Y(n_692) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g841 ( .A(n_633), .Y(n_841) );
INVx2_ASAP7_75t_L g952 ( .A(n_633), .Y(n_952) );
BUFx2_ASAP7_75t_L g699 ( .A(n_637), .Y(n_699) );
BUFx2_ASAP7_75t_L g718 ( .A(n_637), .Y(n_718) );
INVx1_ASAP7_75t_L g848 ( .A(n_637), .Y(n_848) );
BUFx4f_ASAP7_75t_SL g936 ( .A(n_637), .Y(n_936) );
INVx2_ASAP7_75t_L g702 ( .A(n_640), .Y(n_702) );
OA22x2_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_661), .B2(n_701), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AO22x2_ASAP7_75t_L g882 ( .A1(n_643), .A2(n_644), .B1(n_883), .B2(n_899), .Y(n_882) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
XOR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_659), .Y(n_644) );
NAND2x1_ASAP7_75t_L g645 ( .A(n_646), .B(n_652), .Y(n_645) );
NOR2x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVxp67_ASAP7_75t_L g985 ( .A(n_650), .Y(n_985) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_653), .B(n_656), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx2_ASAP7_75t_L g701 ( .A(n_661), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_677), .C(n_686), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_671), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B1(n_668), .B2(n_669), .Y(n_664) );
INVx2_ASAP7_75t_L g783 ( .A(n_665), .Y(n_783) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g1070 ( .A(n_678), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_682), .Y(n_725) );
INVx1_ASAP7_75t_L g854 ( .A(n_682), .Y(n_854) );
INVx2_ASAP7_75t_L g737 ( .A(n_685), .Y(n_737) );
INVx2_ASAP7_75t_L g788 ( .A(n_685), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_685), .A2(n_1059), .B1(n_1060), .B2(n_1061), .Y(n_1058) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_694), .Y(n_686) );
OAI221xp5_ASAP7_75t_L g1052 ( .A1(n_689), .A2(n_1053), .B1(n_1054), .B2(n_1055), .C(n_1056), .Y(n_1052) );
INVx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .Y(n_694) );
INVx2_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_697), .A2(n_980), .B1(n_981), .B2(n_982), .Y(n_979) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_777), .B(n_901), .Y(n_703) );
INVx4_ASAP7_75t_L g903 ( .A(n_704), .Y(n_903) );
OA22x2_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_761), .B2(n_776), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_732), .B1(n_756), .B2(n_757), .Y(n_706) );
INVx1_ASAP7_75t_SL g756 ( .A(n_707), .Y(n_756) );
OR2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_720), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .C(n_714), .D(n_717), .Y(n_709) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx3_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_716), .A2(n_843), .B1(n_844), .B2(n_845), .Y(n_842) );
NAND4xp25_ASAP7_75t_L g720 ( .A(n_721), .B(n_724), .C(n_726), .D(n_728), .Y(n_720) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_733), .Y(n_760) );
INVx1_ASAP7_75t_L g755 ( .A(n_734), .Y(n_755) );
NOR2x1_ASAP7_75t_SL g759 ( .A(n_734), .B(n_760), .Y(n_759) );
NAND4xp75_ASAP7_75t_L g734 ( .A(n_735), .B(n_741), .C(n_745), .D(n_751), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
AND2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx2_ASAP7_75t_SL g844 ( .A(n_748), .Y(n_844) );
INVx4_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g814 ( .A(n_749), .Y(n_814) );
BUFx6f_ASAP7_75t_SL g1024 ( .A(n_750), .Y(n_1024) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx3_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g776 ( .A(n_761), .Y(n_776) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
XNOR2x1_ASAP7_75t_L g804 ( .A(n_762), .B(n_805), .Y(n_804) );
XNOR2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_775), .Y(n_762) );
NOR2x1_ASAP7_75t_L g763 ( .A(n_764), .B(n_769), .Y(n_763) );
NAND4xp25_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .C(n_767), .D(n_768), .Y(n_764) );
NAND4xp25_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .C(n_773), .D(n_774), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_777), .B(n_902), .Y(n_901) );
XNOR2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_831), .Y(n_777) );
OA22x2_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_803), .B1(n_804), .B2(n_830), .Y(n_778) );
INVx1_ASAP7_75t_L g830 ( .A(n_779), .Y(n_830) );
XOR2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_802), .Y(n_779) );
NOR2x1_ASAP7_75t_L g780 ( .A(n_781), .B(n_793), .Y(n_780) );
NAND4xp25_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .C(n_789), .D(n_791), .Y(n_781) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND4xp25_ASAP7_75t_L g793 ( .A(n_794), .B(n_797), .C(n_800), .D(n_801), .Y(n_793) );
INVx2_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
OAI21xp5_ASAP7_75t_SL g886 ( .A1(n_796), .A2(n_887), .B(n_888), .Y(n_886) );
BUFx6f_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND2x1_ASAP7_75t_L g806 ( .A(n_807), .B(n_818), .Y(n_806) );
NOR2x1_ASAP7_75t_L g807 ( .A(n_808), .B(n_812), .Y(n_807) );
OAI21xp5_ASAP7_75t_SL g808 ( .A1(n_809), .A2(n_810), .B(n_811), .Y(n_808) );
OAI21xp33_ASAP7_75t_L g928 ( .A1(n_809), .A2(n_929), .B(n_930), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_815), .Y(n_812) );
NOR2x1_ASAP7_75t_L g818 ( .A(n_819), .B(n_824), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_828), .Y(n_824) );
INVx2_ASAP7_75t_SL g826 ( .A(n_827), .Y(n_826) );
BUFx2_ASAP7_75t_L g1074 ( .A(n_829), .Y(n_1074) );
AO22x2_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_881), .B1(n_882), .B2(n_900), .Y(n_831) );
INVx1_ASAP7_75t_L g900 ( .A(n_832), .Y(n_900) );
XNOR2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_860), .Y(n_832) );
OAI21x1_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_835), .B(n_859), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_834), .B(n_837), .Y(n_859) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_850), .Y(n_837) );
NOR4xp75_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .C(n_842), .D(n_846), .Y(n_838) );
INVx1_ASAP7_75t_L g1005 ( .A(n_844), .Y(n_1005) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_856), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_852), .B(n_855), .Y(n_851) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g1002 ( .A(n_854), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
INVx2_ASAP7_75t_SL g879 ( .A(n_861), .Y(n_879) );
AND2x2_ASAP7_75t_L g861 ( .A(n_862), .B(n_870), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_867), .Y(n_862) );
OAI21xp33_ASAP7_75t_SL g863 ( .A1(n_864), .A2(n_865), .B(n_866), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_875), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_874), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_876), .B(n_878), .Y(n_875) );
INVx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx2_ASAP7_75t_L g899 ( .A(n_883), .Y(n_899) );
NAND2x1_ASAP7_75t_SL g884 ( .A(n_885), .B(n_892), .Y(n_884) );
NOR2x1_ASAP7_75t_L g885 ( .A(n_886), .B(n_889), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
NOR2x1_ASAP7_75t_L g892 ( .A(n_893), .B(n_896), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_967), .B1(n_968), .B2(n_1036), .Y(n_904) );
INVx1_ASAP7_75t_L g1036 ( .A(n_905), .Y(n_1036) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_923), .B1(n_924), .B2(n_966), .Y(n_908) );
INVx5_ASAP7_75t_L g966 ( .A(n_909), .Y(n_966) );
NOR2x1_ASAP7_75t_L g910 ( .A(n_911), .B(n_917), .Y(n_910) );
NAND4xp25_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .C(n_914), .D(n_916), .Y(n_911) );
NAND4xp25_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .C(n_920), .D(n_922), .Y(n_917) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_925), .A2(n_947), .B1(n_948), .B2(n_963), .Y(n_924) );
INVx1_ASAP7_75t_SL g964 ( .A(n_926), .Y(n_964) );
AND2x2_ASAP7_75t_L g926 ( .A(n_927), .B(n_938), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_932), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_933), .B(n_935), .Y(n_932) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_943), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_942), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
INVx1_ASAP7_75t_SL g947 ( .A(n_948), .Y(n_947) );
OR2x2_ASAP7_75t_L g949 ( .A(n_950), .B(n_957), .Y(n_949) );
NAND4xp25_ASAP7_75t_L g950 ( .A(n_951), .B(n_954), .C(n_955), .D(n_956), .Y(n_950) );
NAND4xp25_ASAP7_75t_L g957 ( .A(n_958), .B(n_959), .C(n_960), .D(n_962), .Y(n_957) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
OAI22xp5_ASAP7_75t_SL g968 ( .A1(n_969), .A2(n_1016), .B1(n_1034), .B2(n_1035), .Y(n_968) );
INVx2_ASAP7_75t_SL g1034 ( .A(n_969), .Y(n_1034) );
AO22x2_ASAP7_75t_SL g969 ( .A1(n_970), .A2(n_996), .B1(n_1012), .B2(n_1015), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx2_ASAP7_75t_L g1014 ( .A(n_972), .Y(n_1014) );
INVx1_ASAP7_75t_L g995 ( .A(n_974), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_975), .B(n_988), .Y(n_974) );
NOR3xp33_ASAP7_75t_L g975 ( .A(n_976), .B(n_979), .C(n_983), .Y(n_975) );
NAND2xp5_ASAP7_75t_SL g976 ( .A(n_977), .B(n_978), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_984), .A2(n_985), .B1(n_986), .B2(n_987), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_992), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_991), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
INVx2_ASAP7_75t_L g1015 ( .A(n_996), .Y(n_1015) );
NAND4xp75_ASAP7_75t_L g997 ( .A(n_998), .B(n_1003), .C(n_1007), .D(n_1010), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_999), .B(n_1001), .Y(n_998) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1006), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1016), .Y(n_1035) );
INVx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
XNOR2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
NOR2x1_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1028), .Y(n_1019) );
NAND4xp25_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1023), .C(n_1025), .D(n_1026), .Y(n_1020) );
NAND4xp25_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1030), .C(n_1031), .D(n_1032), .Y(n_1028) );
INVx3_ASAP7_75t_SL g1037 ( .A(n_1038), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1041), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1039), .B(n_1042), .Y(n_1085) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .Y(n_1043) );
OAI222xp33_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1081), .B1(n_1083), .B2(n_1086), .C1(n_1101), .C2(n_1103), .Y(n_1047) );
CKINVDCx16_ASAP7_75t_R g1079 ( .A(n_1049), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
NAND4xp75_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1057), .C(n_1066), .D(n_1076), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
NOR2x1_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1062), .Y(n_1057) );
NOR2x1_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1071), .Y(n_1066) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1078), .Y(n_1076) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_SL g1083 ( .A(n_1084), .Y(n_1083) );
CKINVDCx6p67_ASAP7_75t_R g1084 ( .A(n_1085), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_SL g1102 ( .A(n_1088), .Y(n_1102) );
NOR2x1_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1095), .Y(n_1088) );
NAND4xp25_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1091), .C(n_1093), .D(n_1094), .Y(n_1089) );
NAND4xp25_ASAP7_75t_SL g1095 ( .A(n_1096), .B(n_1097), .C(n_1099), .D(n_1100), .Y(n_1095) );
CKINVDCx20_ASAP7_75t_R g1103 ( .A(n_1104), .Y(n_1103) );
CKINVDCx20_ASAP7_75t_R g1104 ( .A(n_1105), .Y(n_1104) );
endmodule