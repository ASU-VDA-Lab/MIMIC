module fake_netlist_1_11110_n_38 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
OAI22xp5_ASAP7_75t_SL g12 ( .A1(n_9), .A2(n_11), .B1(n_0), .B2(n_7), .Y(n_12) );
AOI22x1_ASAP7_75t_SL g13 ( .A1(n_7), .A2(n_10), .B1(n_4), .B2(n_0), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
AND2x6_ASAP7_75t_L g16 ( .A(n_6), .B(n_1), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_10), .B(n_1), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_14), .B(n_2), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_12), .B(n_2), .Y(n_20) );
OA21x2_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_17), .B(n_16), .Y(n_21) );
OAI21xp5_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_16), .B(n_17), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
OAI221xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_20), .B1(n_21), .B2(n_13), .C(n_16), .Y(n_25) );
NAND2xp5_ASAP7_75t_SL g26 ( .A(n_23), .B(n_21), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
AOI222xp33_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_16), .B1(n_23), .B2(n_21), .C1(n_6), .C2(n_3), .Y(n_29) );
OAI322xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_3), .A3(n_4), .B1(n_5), .B2(n_8), .C1(n_16), .C2(n_20), .Y(n_30) );
OAI21xp5_ASAP7_75t_L g31 ( .A1(n_27), .A2(n_16), .B(n_8), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_29), .Y(n_33) );
NOR2xp33_ASAP7_75t_L g34 ( .A(n_31), .B(n_25), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_33), .B(n_32), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_32), .Y(n_36) );
CKINVDCx20_ASAP7_75t_R g37 ( .A(n_36), .Y(n_37) );
AOI22xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_36), .B1(n_35), .B2(n_34), .Y(n_38) );
endmodule