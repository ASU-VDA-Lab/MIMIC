module fake_jpeg_26822_n_270 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_19),
.Y(n_63)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_51),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_27),
.B1(n_18),
.B2(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_42),
.B1(n_46),
.B2(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_68),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_27),
.B1(n_34),
.B2(n_33),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_62),
.B1(n_42),
.B2(n_23),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_74),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_27),
.B1(n_33),
.B2(n_17),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_73),
.B1(n_36),
.B2(n_38),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_31),
.B1(n_22),
.B2(n_21),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_21),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_22),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_72),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_25),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_35),
.B(n_26),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_36),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_43),
.B1(n_35),
.B2(n_26),
.Y(n_97)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_36),
.A2(n_24),
.B1(n_19),
.B2(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_19),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_30),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_75),
.B(n_43),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_86),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_41),
.B(n_39),
.C(n_37),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_88),
.B1(n_92),
.B2(n_95),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_87),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_41),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_56),
.B(n_37),
.CI(n_44),
.CON(n_87),
.SN(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_42),
.B1(n_43),
.B2(n_28),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_96),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_97),
.B1(n_49),
.B2(n_55),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_92)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_25),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_102),
.Y(n_127)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_39),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_108),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_109),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_26),
.B(n_7),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_110),
.B(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_110),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_48),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_124),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_86),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_55),
.B1(n_49),
.B2(n_76),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_135),
.B1(n_137),
.B2(n_92),
.Y(n_138)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_130),
.B(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_65),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_136),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_72),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_80),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_99),
.A2(n_66),
.B1(n_65),
.B2(n_53),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_53),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_86),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_83),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_157),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_115),
.B1(n_119),
.B2(n_118),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_86),
.B1(n_87),
.B2(n_77),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_145),
.B1(n_149),
.B2(n_128),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_106),
.C(n_86),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_130),
.A2(n_87),
.B1(n_94),
.B2(n_85),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_104),
.B1(n_85),
.B2(n_79),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_161),
.B1(n_128),
.B2(n_125),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_152),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_97),
.B1(n_104),
.B2(n_80),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_96),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_154),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_80),
.C(n_89),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_125),
.C(n_1),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_90),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_121),
.B(n_98),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_78),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_162),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_156),
.B(n_3),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_102),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_163),
.Y(n_183)
);

OAI31xp33_ASAP7_75t_SL g160 ( 
.A1(n_117),
.A2(n_95),
.A3(n_81),
.B(n_93),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_115),
.A3(n_118),
.B1(n_131),
.B2(n_119),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_95),
.B1(n_78),
.B2(n_0),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_136),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_3),
.Y(n_185)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_115),
.A3(n_114),
.B1(n_117),
.B2(n_137),
.C1(n_129),
.C2(n_135),
.Y(n_167)
);

OAI322xp33_ASAP7_75t_L g199 ( 
.A1(n_167),
.A2(n_155),
.A3(n_140),
.B1(n_145),
.B2(n_162),
.C1(n_150),
.C2(n_165),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_178),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_175),
.B1(n_176),
.B2(n_182),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_179),
.B(n_171),
.Y(n_197)
);

XOR2x2_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_125),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_184),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_8),
.C(n_11),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_186),
.Y(n_196)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_4),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_190),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_5),
.B(n_6),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_149),
.B1(n_138),
.B2(n_141),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_200),
.B1(n_203),
.B2(n_209),
.Y(n_211)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_202),
.Y(n_216)
);

AOI321xp33_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_186),
.A3(n_170),
.B1(n_178),
.B2(n_173),
.C(n_180),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_166),
.A2(n_142),
.B1(n_151),
.B2(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_142),
.B1(n_163),
.B2(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_158),
.B1(n_6),
.B2(n_7),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_205),
.A2(n_185),
.B1(n_177),
.B2(n_188),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_158),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_210),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_5),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_210),
.C(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_169),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_225),
.C(n_167),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_171),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_219),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_179),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_220),
.B(n_224),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_181),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_174),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_203),
.B1(n_193),
.B2(n_187),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_189),
.B(n_177),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_223),
.A2(n_226),
.B(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_175),
.B(n_182),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_206),
.C(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_229),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_226),
.B(n_214),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_208),
.C(n_168),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_201),
.B1(n_205),
.B2(n_204),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_233),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_174),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_236),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_235),
.A2(n_211),
.B1(n_238),
.B2(n_228),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_168),
.C(n_201),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_212),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_229),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_241),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_231),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_8),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_244),
.B(n_248),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_12),
.C(n_14),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_223),
.B1(n_215),
.B2(n_216),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_218),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_227),
.Y(n_251)
);

NOR2x1_ASAP7_75t_R g250 ( 
.A(n_242),
.B(n_237),
.Y(n_250)
);

AOI21x1_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_245),
.B(n_247),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_256),
.Y(n_259)
);

OAI221xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_187),
.B1(n_236),
.B2(n_13),
.C(n_14),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_14),
.B(n_15),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_254),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_246),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_260),
.B(n_257),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_250),
.B(n_245),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_264),
.B(n_265),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_263),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_255),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_267),
.A2(n_241),
.B1(n_249),
.B2(n_15),
.Y(n_268)
);

AOI211xp5_ASAP7_75t_SL g269 ( 
.A1(n_268),
.A2(n_15),
.B(n_16),
.C(n_266),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_16),
.Y(n_270)
);


endmodule