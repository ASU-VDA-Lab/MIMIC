module real_jpeg_13706_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_330, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_330;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_2),
.A2(n_40),
.B1(n_54),
.B2(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_40),
.B1(n_59),
.B2(n_60),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_2),
.A2(n_30),
.B1(n_36),
.B2(n_40),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_4),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_35),
.B1(n_54),
.B2(n_57),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_4),
.A2(n_35),
.B1(n_59),
.B2(n_60),
.Y(n_325)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_6),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_6),
.A2(n_54),
.B1(n_57),
.B2(n_182),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_182),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_6),
.A2(n_30),
.B1(n_36),
.B2(n_182),
.Y(n_261)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_7),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_7),
.B(n_185),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_7),
.B(n_57),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_7),
.A2(n_59),
.B(n_221),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g239 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_174),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_7),
.A2(n_42),
.B(n_45),
.C(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_7),
.B(n_79),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_7),
.B(n_33),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_7),
.B(n_50),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g275 ( 
.A1(n_7),
.A2(n_57),
.B(n_212),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_9),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_9),
.A2(n_54),
.B1(n_57),
.B2(n_63),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_63),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_9),
.A2(n_30),
.B1(n_36),
.B2(n_63),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_54),
.B1(n_57),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_10),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_10),
.A2(n_30),
.B1(n_36),
.B2(n_71),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_12),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_12),
.A2(n_54),
.B1(n_57),
.B2(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_155),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_12),
.A2(n_30),
.B1(n_36),
.B2(n_155),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_13),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_13),
.A2(n_54),
.B1(n_57),
.B2(n_119),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_119),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_13),
.A2(n_30),
.B1(n_36),
.B2(n_119),
.Y(n_249)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_15),
.A2(n_49),
.B1(n_54),
.B2(n_57),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_15),
.A2(n_30),
.B1(n_36),
.B2(n_49),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_15),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_16),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_16),
.A2(n_54),
.B1(n_57),
.B2(n_65),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_16),
.A2(n_41),
.B1(n_42),
.B2(n_65),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_16),
.A2(n_30),
.B1(n_36),
.B2(n_65),
.Y(n_202)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_321),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_308),
.B(n_320),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_133),
.B(n_305),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_120),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_96),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_23),
.B(n_96),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_66),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_24),
.B(n_82),
.C(n_94),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_51),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_25),
.A2(n_26),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_37),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_27),
.A2(n_28),
.B1(n_51),
.B2(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_27),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_33),
.B(n_34),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_29),
.A2(n_33),
.B1(n_34),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_29),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_29),
.A2(n_33),
.B1(n_146),
.B2(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_29),
.A2(n_33),
.B1(n_170),
.B2(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_29),
.A2(n_33),
.B1(n_202),
.B2(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_29),
.A2(n_33),
.B1(n_215),
.B2(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_29),
.A2(n_33),
.B1(n_174),
.B2(n_261),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_29),
.A2(n_33),
.B1(n_254),
.B2(n_261),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_30),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_30),
.B(n_263),
.Y(n_262)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_32),
.A2(n_110),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_32),
.A2(n_144),
.B1(n_253),
.B2(n_255),
.Y(n_252)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_36),
.A2(n_46),
.B(n_174),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_39),
.A2(n_43),
.B1(n_50),
.B2(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_42),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g210 ( 
.A1(n_41),
.A2(n_57),
.A3(n_75),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_42),
.B(n_76),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_48),
.B1(n_50),
.B2(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_50),
.B(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_43),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_43),
.A2(n_50),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_43),
.A2(n_50),
.B1(n_149),
.B2(n_206),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_43),
.A2(n_50),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_43),
.A2(n_50),
.B1(n_240),
.B2(n_247),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_47),
.A2(n_114),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_47),
.A2(n_150),
.B1(n_205),
.B2(n_277),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_64),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_53),
.B1(n_64),
.B2(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_52),
.A2(n_53),
.B1(n_85),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_52),
.A2(n_53),
.B1(n_118),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_52),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_52),
.A2(n_53),
.B1(n_181),
.B2(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_53),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_57),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_54),
.A2(n_56),
.A3(n_59),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_55),
.B(n_57),
.Y(n_172)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_60),
.B(n_174),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_82),
.B1(n_94),
.B2(n_95),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_68),
.B(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_80),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B1(n_78),
.B2(n_79),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_73),
.B1(n_77),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_78),
.B1(n_79),
.B2(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_72),
.A2(n_79),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_72),
.A2(n_79),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_72),
.A2(n_79),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_73),
.A2(n_77),
.B1(n_92),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_73),
.A2(n_77),
.B1(n_116),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_73),
.A2(n_77),
.B1(n_177),
.B2(n_198),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_73),
.A2(n_77),
.B1(n_196),
.B2(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_84),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_88),
.C(n_90),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_84),
.B(n_123),
.C(n_126),
.Y(n_309)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_93),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_93),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_88),
.B(n_129),
.C(n_131),
.Y(n_319)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.C(n_104),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_157)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.C(n_117),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_106),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_117),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_120),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_121),
.B(n_122),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_130),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_132),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_158),
.B(n_304),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_156),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_135),
.B(n_156),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_140),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_151),
.C(n_153),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_142),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_143),
.B(n_147),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_153),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_188),
.B(n_303),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_186),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_160),
.B(n_186),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.C(n_166),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_165),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_166),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_175),
.C(n_179),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_167),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_173),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_175),
.B(n_179),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_183),
.A2(n_185),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_183),
.A2(n_185),
.B1(n_316),
.B2(n_325),
.Y(n_324)
);

OAI221xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_296),
.B1(n_301),
.B2(n_302),
.C(n_330),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_288),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_232),
.B(n_287),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_216),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_192),
.B(n_216),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_203),
.C(n_207),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_193),
.B(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_200),
.C(n_201),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_203),
.A2(n_207),
.B1(n_208),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_203),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_214),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_227),
.B2(n_231),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_217),
.B(n_228),
.C(n_230),
.Y(n_289)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_219),
.B(n_223),
.C(n_226),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_227),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_281),
.B(n_286),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_270),
.B(n_280),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_250),
.B(n_269),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_243),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_236),
.B(n_243),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_246),
.C(n_248),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_249),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_258),
.B(n_268),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_256),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_264),
.B(n_267),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_265),
.B(n_266),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_271),
.B(n_272),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_276),
.C(n_278),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_290),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.C(n_294),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_298),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_310),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_319),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_314),
.B1(n_317),
.B2(n_318),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_312),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_317),
.C(n_319),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_328),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_327),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_327),
.Y(n_326)
);


endmodule