module fake_ariane_2541_n_2005 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2005);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2005;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_158),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_66),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_91),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_41),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_18),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_32),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_95),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_107),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_65),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_43),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_8),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_61),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_153),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_111),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_139),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_53),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_143),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_13),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_49),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_127),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_99),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_159),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_28),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_46),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_55),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_126),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_68),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_179),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_145),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_124),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_110),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_29),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_108),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_10),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_151),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_148),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_7),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_58),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_10),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_117),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_30),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_152),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_9),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_42),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_50),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_64),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_115),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_27),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_96),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_147),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_150),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_131),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_36),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_78),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_135),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_171),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_144),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_82),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_74),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_90),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_183),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_184),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_57),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_25),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_113),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_167),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_92),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_41),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_128),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_142),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_97),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_3),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_60),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_89),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_70),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_65),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_138),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_132),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_16),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_35),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_76),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_83),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_191),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_67),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_157),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_76),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_130),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_123),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_56),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_149),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_168),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_21),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_4),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_21),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_190),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_121),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_134),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_37),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_50),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_176),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_59),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_109),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_11),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_178),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_141),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_64),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_94),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_63),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_120),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_114),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_162),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_32),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_26),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_51),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_8),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_36),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_56),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_98),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_55),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_23),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_23),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_33),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_52),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_186),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_71),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_60),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_71),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_39),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_2),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_165),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_49),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_53),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_172),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_100),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_181),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_61),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_80),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_88),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_154),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_73),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_25),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_122),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_74),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_105),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_31),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_3),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_119),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_79),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_5),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_140),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_112),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_22),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_16),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_59),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_24),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_18),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_169),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_102),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_81),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_6),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_29),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_31),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_37),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_68),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_33),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_73),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_14),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_69),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_170),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_19),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_5),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_42),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_38),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_84),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_160),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_57),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_20),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_58),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_30),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_1),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_35),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_0),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_200),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_R g389 ( 
.A(n_261),
.B(n_290),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_198),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_346),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_346),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_346),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_340),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_264),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_358),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_201),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_202),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_201),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_358),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_204),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_360),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_333),
.B(n_0),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_204),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_213),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_213),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_219),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_256),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_203),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_222),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_219),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_360),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_223),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_194),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_236),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_264),
.B(n_1),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_333),
.B(n_369),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_196),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_236),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_237),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_237),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_303),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_202),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_308),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_241),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_197),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_205),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_241),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_243),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_211),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_214),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_224),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_198),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_226),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_243),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_334),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_235),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_247),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_247),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_238),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_245),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_256),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_254),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_246),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_254),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_258),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_248),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_337),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_257),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_258),
.B(n_2),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_270),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_270),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_271),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_257),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_251),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_271),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_273),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_263),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_273),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_293),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_267),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_293),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_R g463 ( 
.A(n_193),
.B(n_129),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_275),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_307),
.B(n_6),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_275),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_275),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_307),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_369),
.B(n_7),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_309),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_309),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_314),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_314),
.B(n_9),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_R g474 ( 
.A(n_195),
.B(n_125),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_295),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_216),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_323),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_216),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_323),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_268),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_339),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_280),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_390),
.B(n_198),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_393),
.B(n_339),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_408),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_416),
.B(n_256),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_390),
.B(n_433),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_392),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_391),
.B(n_343),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_397),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_397),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_399),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_399),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_401),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_401),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_433),
.B(n_206),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_404),
.B(n_405),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_404),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_405),
.B(n_206),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_406),
.B(n_206),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_406),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_407),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_407),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_396),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_400),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_411),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_415),
.B(n_419),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_415),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_419),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_420),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_420),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_421),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_421),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_425),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_428),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_428),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_429),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_435),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_389),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_435),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

CKINVDCx8_ASAP7_75t_R g533 ( 
.A(n_388),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_438),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_439),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_439),
.B(n_328),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_443),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_443),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_SL g539 ( 
.A(n_464),
.B(n_369),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_449),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_445),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_445),
.B(n_343),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_446),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_451),
.B(n_344),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_451),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_395),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_452),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_452),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_387),
.B(n_376),
.Y(n_550)
);

BUFx8_ASAP7_75t_L g551 ( 
.A(n_395),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_453),
.B(n_328),
.Y(n_552)
);

BUFx8_ASAP7_75t_L g553 ( 
.A(n_453),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_456),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_456),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_457),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_457),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_459),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_459),
.B(n_328),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_460),
.B(n_295),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_460),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_462),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_496),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_496),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_496),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_533),
.A2(n_409),
.B1(n_422),
.B2(n_410),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_496),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_496),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_496),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_496),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_553),
.B(n_418),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_553),
.B(n_218),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_496),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_496),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_497),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_530),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_553),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_488),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_550),
.B(n_465),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_490),
.B(n_413),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_488),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_488),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_497),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_488),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_553),
.B(n_426),
.Y(n_585)
);

INVx6_ASAP7_75t_L g586 ( 
.A(n_553),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_553),
.B(n_427),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_485),
.B(n_430),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_488),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_560),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_502),
.B(n_432),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_497),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_497),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_502),
.B(n_462),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_502),
.B(n_218),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_502),
.B(n_468),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_SL g597 ( 
.A(n_517),
.B(n_434),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_502),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_497),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_497),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_502),
.B(n_437),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_513),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_485),
.B(n_468),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_497),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_490),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_547),
.B(n_440),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_488),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_513),
.B(n_470),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_513),
.B(n_470),
.Y(n_609)
);

BUFx4f_ASAP7_75t_L g610 ( 
.A(n_560),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_497),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_491),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_560),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_497),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_503),
.B(n_218),
.Y(n_615)
);

CKINVDCx11_ASAP7_75t_R g616 ( 
.A(n_533),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_551),
.B(n_441),
.Y(n_617)
);

INVx6_ASAP7_75t_L g618 ( 
.A(n_505),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_500),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_547),
.B(n_444),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_550),
.A2(n_450),
.B1(n_473),
.B2(n_469),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_491),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_551),
.B(n_455),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_513),
.B(n_471),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_513),
.B(n_471),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_551),
.B(n_458),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_491),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_500),
.Y(n_628)
);

BUFx6f_ASAP7_75t_SL g629 ( 
.A(n_560),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_551),
.B(n_461),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_551),
.B(n_480),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_551),
.B(n_482),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_490),
.B(n_466),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_550),
.A2(n_560),
.B1(n_505),
.B2(n_552),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_500),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_504),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_483),
.B(n_467),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_491),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_513),
.B(n_472),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_536),
.B(n_472),
.Y(n_640)
);

XNOR2x2_ASAP7_75t_R g641 ( 
.A(n_533),
.B(n_424),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_491),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_500),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_500),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_500),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_500),
.Y(n_646)
);

INVxp67_ASAP7_75t_SL g647 ( 
.A(n_515),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_500),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_521),
.B(n_477),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_550),
.B(n_398),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_500),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_550),
.A2(n_560),
.B1(n_505),
.B2(n_552),
.Y(n_652)
);

CKINVDCx6p67_ASAP7_75t_R g653 ( 
.A(n_504),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_507),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_507),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_483),
.B(n_475),
.Y(n_656)
);

AO21x2_ASAP7_75t_L g657 ( 
.A1(n_487),
.A2(n_349),
.B(n_344),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_507),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_504),
.B(n_431),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_L g660 ( 
.A(n_507),
.B(n_256),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_507),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_483),
.B(n_447),
.Y(n_662)
);

BUFx8_ASAP7_75t_SL g663 ( 
.A(n_540),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_491),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_501),
.B(n_454),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_507),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_507),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_507),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_550),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_504),
.B(n_403),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_501),
.B(n_477),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_507),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_516),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_501),
.B(n_524),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_524),
.B(n_479),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_516),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_521),
.B(n_535),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_516),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_516),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_517),
.B(n_479),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_516),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_516),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_550),
.A2(n_240),
.B1(n_244),
.B2(n_239),
.Y(n_683)
);

BUFx8_ASAP7_75t_SL g684 ( 
.A(n_540),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_510),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_516),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_550),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_516),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_527),
.B(n_481),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_527),
.B(n_481),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_516),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_526),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_487),
.A2(n_476),
.B1(n_423),
.B2(n_478),
.Y(n_693)
);

BUFx10_ASAP7_75t_L g694 ( 
.A(n_510),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_536),
.B(n_417),
.Y(n_695)
);

INVxp33_ASAP7_75t_L g696 ( 
.A(n_511),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_526),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_561),
.B(n_253),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_526),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_526),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_517),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_540),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_521),
.B(n_417),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_526),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_536),
.B(n_233),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_521),
.B(n_231),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_521),
.B(n_282),
.Y(n_707)
);

OAI21xp33_ASAP7_75t_SL g708 ( 
.A1(n_515),
.A2(n_276),
.B(n_242),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_526),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_511),
.A2(n_367),
.B1(n_318),
.B2(n_317),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_560),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_514),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_514),
.B(n_233),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_560),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_561),
.B(n_394),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_580),
.B(n_436),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_578),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_588),
.B(n_539),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_578),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_586),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_610),
.B(n_526),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_598),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_650),
.A2(n_463),
.B1(n_474),
.B2(n_560),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_581),
.Y(n_724)
);

AND2x4_ASAP7_75t_SL g725 ( 
.A(n_653),
.B(n_448),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_696),
.B(n_539),
.Y(n_726)
);

BUFx5_ASAP7_75t_L g727 ( 
.A(n_577),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_SL g728 ( 
.A(n_636),
.B(n_653),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_598),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_581),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_606),
.B(n_521),
.Y(n_731)
);

INVxp67_ASAP7_75t_SL g732 ( 
.A(n_577),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_582),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_582),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_669),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_647),
.B(n_535),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_671),
.B(n_535),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_603),
.B(n_535),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_674),
.B(n_535),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_620),
.B(n_535),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_586),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_610),
.B(n_526),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_705),
.B(n_505),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_602),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_712),
.B(n_538),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_584),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_584),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_591),
.B(n_538),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_669),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_640),
.B(n_538),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_601),
.B(n_538),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_580),
.B(n_505),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_680),
.B(n_538),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_640),
.B(n_538),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_715),
.B(n_503),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_633),
.B(n_505),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_705),
.B(n_503),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_610),
.B(n_613),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_589),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_602),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_650),
.B(n_508),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_650),
.B(n_506),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_650),
.B(n_508),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_595),
.B(n_526),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_SL g765 ( 
.A(n_636),
.B(n_335),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_662),
.B(n_508),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_637),
.B(n_506),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_675),
.B(n_518),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_613),
.B(n_529),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_586),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_613),
.B(n_529),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_589),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_656),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_689),
.B(n_518),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_711),
.B(n_529),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_690),
.B(n_518),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_665),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_714),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_698),
.B(n_519),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_607),
.Y(n_780)
);

OAI22x1_ASAP7_75t_SL g781 ( 
.A1(n_641),
.A2(n_285),
.B1(n_297),
.B2(n_281),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_695),
.B(n_687),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_687),
.A2(n_560),
.B1(n_552),
.B2(n_559),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_677),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_695),
.B(n_519),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_711),
.B(n_529),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_605),
.B(n_519),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_607),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_579),
.A2(n_560),
.B1(n_552),
.B2(n_559),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_711),
.B(n_529),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_714),
.B(n_529),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_618),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_605),
.B(n_522),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_594),
.B(n_522),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_612),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_596),
.B(n_522),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_701),
.B(n_506),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_693),
.B(n_523),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_693),
.B(n_523),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_597),
.B(n_336),
.C(n_284),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_572),
.A2(n_560),
.B1(n_506),
.B2(n_559),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_618),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_702),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_621),
.B(n_523),
.Y(n_804)
);

NOR2xp67_ASAP7_75t_L g805 ( 
.A(n_617),
.B(n_542),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_618),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_579),
.A2(n_552),
.B1(n_559),
.B2(n_506),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_706),
.B(n_528),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_618),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_707),
.B(n_528),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_612),
.Y(n_811)
);

NOR2x1_ASAP7_75t_L g812 ( 
.A(n_623),
.B(n_542),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_L g813 ( 
.A(n_710),
.B(n_531),
.C(n_528),
.Y(n_813)
);

INVxp33_ASAP7_75t_L g814 ( 
.A(n_566),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_595),
.B(n_531),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_634),
.B(n_506),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_595),
.B(n_531),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_579),
.A2(n_548),
.B1(n_554),
.B2(n_532),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_713),
.B(n_532),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_595),
.B(n_532),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_595),
.B(n_703),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_622),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_595),
.B(n_548),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_708),
.A2(n_554),
.B(n_555),
.C(n_548),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_572),
.A2(n_559),
.B1(n_552),
.B2(n_555),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_595),
.B(n_554),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_608),
.B(n_555),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_L g828 ( 
.A(n_564),
.B(n_529),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_622),
.Y(n_829)
);

INVx8_ASAP7_75t_L g830 ( 
.A(n_572),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_627),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_685),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_714),
.B(n_529),
.Y(n_833)
);

OAI221xp5_ASAP7_75t_L g834 ( 
.A1(n_683),
.A2(n_361),
.B1(n_277),
.B2(n_279),
.C(n_286),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_652),
.B(n_529),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_627),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_609),
.B(n_556),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_624),
.B(n_556),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_638),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_683),
.B(n_559),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_625),
.A2(n_492),
.B(n_545),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_572),
.A2(n_579),
.B1(n_615),
.B2(n_657),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_659),
.B(n_556),
.Y(n_843)
);

O2A1O1Ixp5_ASAP7_75t_L g844 ( 
.A1(n_567),
.A2(n_558),
.B(n_484),
.C(n_492),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_639),
.B(n_558),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_638),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_564),
.B(n_537),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_663),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_572),
.A2(n_558),
.B1(n_537),
.B2(n_549),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_685),
.B(n_545),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_590),
.B(n_495),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_642),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_670),
.B(n_484),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_685),
.B(n_495),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_685),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_649),
.B(n_495),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_694),
.B(n_495),
.Y(n_857)
);

AOI221xp5_ASAP7_75t_L g858 ( 
.A1(n_708),
.A2(n_351),
.B1(n_276),
.B2(n_242),
.C(n_277),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_642),
.Y(n_859)
);

INVx6_ASAP7_75t_L g860 ( 
.A(n_576),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_664),
.Y(n_861)
);

INVx8_ASAP7_75t_L g862 ( 
.A(n_572),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_664),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_572),
.B(n_498),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_694),
.B(n_576),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_579),
.B(n_498),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_694),
.B(n_498),
.Y(n_867)
);

OAI22xp33_ASAP7_75t_L g868 ( 
.A1(n_586),
.A2(n_702),
.B1(n_630),
.B2(n_631),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_564),
.B(n_537),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_657),
.B(n_498),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_694),
.B(n_499),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_615),
.A2(n_537),
.B1(n_549),
.B2(n_335),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_626),
.B(n_499),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_666),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_666),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_564),
.Y(n_876)
);

NOR2xp67_ASAP7_75t_L g877 ( 
.A(n_632),
.B(n_499),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_567),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_564),
.B(n_575),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_575),
.B(n_537),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_615),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_684),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_615),
.A2(n_537),
.B1(n_549),
.B2(n_335),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_672),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_657),
.B(n_499),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_571),
.B(n_585),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_566),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_587),
.B(n_509),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_879),
.A2(n_565),
.B(n_563),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_718),
.B(n_616),
.C(n_549),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_879),
.A2(n_565),
.B(n_563),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_722),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_717),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_755),
.B(n_576),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_808),
.A2(n_570),
.B(n_568),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_766),
.B(n_576),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_716),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_725),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_731),
.B(n_575),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_725),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_810),
.A2(n_736),
.B(n_737),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_729),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_738),
.A2(n_570),
.B(n_568),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_850),
.B(n_615),
.Y(n_904)
);

AOI21x1_ASAP7_75t_L g905 ( 
.A1(n_721),
.A2(n_574),
.B(n_573),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_762),
.B(n_590),
.Y(n_906)
);

BUFx8_ASAP7_75t_L g907 ( 
.A(n_832),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_773),
.B(n_567),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_740),
.B(n_615),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_781),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_803),
.Y(n_911)
);

O2A1O1Ixp5_ASAP7_75t_L g912 ( 
.A1(n_779),
.A2(n_619),
.B(n_643),
.C(n_569),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_816),
.A2(n_834),
.B1(n_840),
.B2(n_814),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_757),
.B(n_615),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_L g915 ( 
.A(n_777),
.B(n_286),
.C(n_279),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_752),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_756),
.B(n_569),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_769),
.A2(n_574),
.B(n_573),
.Y(n_918)
);

AOI21xp33_ASAP7_75t_L g919 ( 
.A1(n_814),
.A2(n_673),
.B(n_672),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_743),
.B(n_509),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_741),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_844),
.A2(n_592),
.B(n_583),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_769),
.A2(n_775),
.B(n_771),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_771),
.A2(n_592),
.B(n_583),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_775),
.A2(n_599),
.B(n_593),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_750),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_741),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_787),
.A2(n_793),
.B(n_804),
.C(n_858),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_841),
.A2(n_599),
.B(n_593),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_717),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_726),
.B(n_569),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_840),
.B(n_509),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_743),
.B(n_509),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_761),
.A2(n_512),
.B(n_525),
.C(n_520),
.Y(n_934)
);

OAI321xp33_ASAP7_75t_L g935 ( 
.A1(n_868),
.A2(n_373),
.A3(n_351),
.B1(n_313),
.B2(n_306),
.C(n_359),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_848),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_745),
.B(n_512),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_854),
.B(n_512),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_778),
.B(n_575),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_786),
.A2(n_604),
.B(n_600),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_719),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_857),
.B(n_512),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_786),
.A2(n_604),
.B(n_600),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_790),
.A2(n_614),
.B(n_611),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_767),
.B(n_619),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_867),
.B(n_520),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_790),
.A2(n_833),
.B(n_791),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_871),
.B(n_782),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_792),
.B(n_619),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_791),
.A2(n_614),
.B(n_611),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_833),
.A2(n_635),
.B(n_628),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_763),
.B(n_520),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_856),
.A2(n_635),
.B(n_628),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_754),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_816),
.B(n_520),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_797),
.B(n_525),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_819),
.B(n_525),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_802),
.B(n_643),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_887),
.B(n_525),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_806),
.B(n_809),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_719),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_768),
.A2(n_643),
.B1(n_676),
.B2(n_646),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_762),
.B(n_534),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_860),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_721),
.A2(n_645),
.B(n_644),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_762),
.B(n_843),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_741),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_724),
.Y(n_968)
);

NOR2xp67_ASAP7_75t_L g969 ( 
.A(n_882),
.B(n_641),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_741),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_832),
.B(n_534),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_778),
.B(n_575),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_774),
.A2(n_645),
.B(n_644),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_765),
.B(n_646),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_855),
.B(n_534),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_784),
.B(n_646),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_855),
.B(n_534),
.Y(n_977)
);

BUFx12f_ASAP7_75t_L g978 ( 
.A(n_860),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_776),
.A2(n_699),
.B1(n_700),
.B2(n_676),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_785),
.A2(n_651),
.B(n_648),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_873),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_742),
.A2(n_651),
.B(n_648),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_865),
.B(n_735),
.Y(n_983)
);

BUFx8_ASAP7_75t_L g984 ( 
.A(n_873),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_L g985 ( 
.A(n_800),
.B(n_294),
.C(n_289),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_778),
.B(n_655),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_720),
.B(n_590),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_873),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_735),
.B(n_749),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_742),
.A2(n_658),
.B(n_654),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_748),
.A2(n_541),
.B(n_544),
.C(n_543),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_753),
.B(n_541),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_724),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_749),
.B(n_541),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_739),
.B(n_541),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_805),
.A2(n_629),
.B1(n_658),
.B2(n_654),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_827),
.A2(n_667),
.B(n_661),
.Y(n_997)
);

AOI21xp33_ASAP7_75t_L g998 ( 
.A1(n_751),
.A2(n_678),
.B(n_673),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_822),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_837),
.A2(n_845),
.B(n_838),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_818),
.B(n_655),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_860),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_728),
.Y(n_1003)
);

INVxp67_ASAP7_75t_L g1004 ( 
.A(n_798),
.Y(n_1004)
);

OAI21xp33_ASAP7_75t_SL g1005 ( 
.A1(n_815),
.A2(n_667),
.B(n_661),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_794),
.A2(n_686),
.B(n_668),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_796),
.A2(n_686),
.B(n_668),
.Y(n_1007)
);

AO21x1_ASAP7_75t_L g1008 ( 
.A1(n_870),
.A2(n_362),
.B(n_349),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_723),
.A2(n_853),
.B1(n_807),
.B2(n_812),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_799),
.B(n_543),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_732),
.B(n_543),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_744),
.B(n_676),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_813),
.B(n_543),
.Y(n_1013)
);

BUFx4f_ASAP7_75t_L g1014 ( 
.A(n_760),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_824),
.A2(n_544),
.B(n_546),
.C(n_557),
.Y(n_1015)
);

OAI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_789),
.A2(n_376),
.B1(n_291),
.B2(n_384),
.Y(n_1016)
);

BUFx8_ASAP7_75t_L g1017 ( 
.A(n_829),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_876),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_831),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_847),
.A2(n_880),
.B(n_869),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_847),
.A2(n_880),
.B(n_869),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_886),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_876),
.Y(n_1023)
);

AO21x1_ASAP7_75t_L g1024 ( 
.A1(n_885),
.A2(n_374),
.B(n_362),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_828),
.A2(n_704),
.B(n_691),
.Y(n_1025)
);

AO21x1_ASAP7_75t_L g1026 ( 
.A1(n_864),
.A2(n_374),
.B(n_691),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_828),
.A2(n_704),
.B(n_679),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_878),
.B(n_699),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_878),
.A2(n_679),
.B(n_678),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_878),
.A2(n_688),
.B(n_682),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_824),
.A2(n_866),
.B(n_820),
.C(n_823),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_874),
.A2(n_688),
.B(n_682),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_875),
.A2(n_697),
.B(n_692),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_836),
.A2(n_544),
.B(n_546),
.C(n_557),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_839),
.A2(n_546),
.B(n_557),
.C(n_562),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_730),
.B(n_733),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_733),
.B(n_546),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_884),
.A2(n_697),
.B(n_692),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_876),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_835),
.A2(n_821),
.B(n_888),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_734),
.A2(n_709),
.B(n_700),
.Y(n_1041)
);

O2A1O1Ixp5_ASAP7_75t_L g1042 ( 
.A1(n_817),
.A2(n_700),
.B(n_699),
.C(n_709),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_734),
.B(n_557),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_746),
.A2(n_681),
.B(n_655),
.Y(n_1044)
);

OAI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_826),
.A2(n_299),
.B(n_298),
.Y(n_1045)
);

NOR3xp33_ASAP7_75t_L g1046 ( 
.A(n_764),
.B(n_294),
.C(n_289),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_746),
.B(n_562),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_747),
.A2(n_681),
.B(n_655),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_846),
.Y(n_1049)
);

OAI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_852),
.A2(n_311),
.B(n_304),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_747),
.B(n_562),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_759),
.B(n_537),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_772),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_772),
.A2(n_681),
.B(n_655),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_780),
.B(n_537),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_861),
.B(n_681),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_876),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_780),
.B(n_537),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_788),
.B(n_549),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_788),
.B(n_233),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_795),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_835),
.A2(n_629),
.B1(n_376),
.B2(n_233),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_795),
.A2(n_681),
.B(n_590),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_811),
.A2(n_590),
.B(n_660),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_811),
.B(n_549),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_859),
.A2(n_590),
.B(n_262),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_859),
.B(n_306),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_863),
.A2(n_758),
.B(n_764),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_863),
.A2(n_320),
.B(n_319),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_851),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_758),
.A2(n_549),
.B(n_207),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_783),
.A2(n_494),
.B(n_301),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_825),
.B(n_549),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_881),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_877),
.B(n_549),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_881),
.B(n_229),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_801),
.B(n_313),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_842),
.B(n_324),
.Y(n_1078)
);

OAI21xp33_ASAP7_75t_L g1079 ( 
.A1(n_872),
.A2(n_322),
.B(n_321),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_851),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1000),
.A2(n_862),
.B(n_830),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_916),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_894),
.B(n_720),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_911),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_913),
.B(n_883),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_897),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_959),
.B(n_325),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_1039),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_898),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_913),
.B(n_326),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_893),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_896),
.B(n_727),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_928),
.B(n_330),
.C(n_327),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1022),
.B(n_341),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_929),
.A2(n_849),
.B(n_493),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_905),
.A2(n_493),
.B(n_494),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_966),
.B(n_720),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_SL g1098 ( 
.A(n_969),
.B(n_770),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1039),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_928),
.A2(n_862),
.B(n_830),
.C(n_329),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_999),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_SL g1102 ( 
.A1(n_945),
.A2(n_908),
.B(n_917),
.C(n_931),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_932),
.B(n_727),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_909),
.A2(n_862),
.B(n_830),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_948),
.B(n_770),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1060),
.B(n_926),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_931),
.A2(n_862),
.B(n_830),
.C(n_329),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_954),
.B(n_727),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_930),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_901),
.A2(n_770),
.B(n_727),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_SL g1111 ( 
.A1(n_945),
.A2(n_361),
.B(n_331),
.C(n_332),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_900),
.B(n_324),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_981),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_915),
.A2(n_332),
.B(n_373),
.C(n_371),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_906),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1078),
.A2(n_335),
.B1(n_384),
.B2(n_331),
.Y(n_1116)
);

INVx5_ASAP7_75t_L g1117 ( 
.A(n_906),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1009),
.B(n_727),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1003),
.B(n_727),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1039),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_908),
.A2(n_359),
.B(n_365),
.C(n_371),
.Y(n_1121)
);

AO22x1_ASAP7_75t_L g1122 ( 
.A1(n_1017),
.A2(n_378),
.B1(n_350),
.B2(n_357),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_SL g1123 ( 
.A(n_936),
.B(n_629),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_978),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_985),
.A2(n_365),
.B(n_291),
.C(n_301),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_983),
.B(n_345),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_938),
.A2(n_229),
.B(n_301),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_983),
.B(n_229),
.Y(n_1128)
);

OAI21xp33_ASAP7_75t_SL g1129 ( 
.A1(n_1001),
.A2(n_363),
.B(n_232),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_965),
.A2(n_493),
.B(n_494),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_988),
.B(n_348),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_1039),
.Y(n_1132)
);

CKINVDCx10_ASAP7_75t_R g1133 ( 
.A(n_910),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_906),
.Y(n_1134)
);

NOR2x1_ASAP7_75t_L g1135 ( 
.A(n_890),
.B(n_921),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_923),
.A2(n_363),
.B(n_493),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1016),
.A2(n_904),
.B1(n_974),
.B2(n_917),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_970),
.Y(n_1138)
);

NAND2xp33_ASAP7_75t_R g1139 ( 
.A(n_987),
.B(n_199),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_930),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1067),
.B(n_354),
.Y(n_1141)
);

AOI222xp33_ASAP7_75t_L g1142 ( 
.A1(n_935),
.A2(n_377),
.B1(n_386),
.B2(n_385),
.C1(n_383),
.C2(n_382),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_941),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_970),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_970),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_920),
.A2(n_363),
.B(n_232),
.C(n_295),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_R g1147 ( 
.A(n_978),
.B(n_366),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_956),
.B(n_368),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_955),
.B(n_892),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_942),
.A2(n_305),
.B(n_208),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1016),
.B(n_370),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_946),
.A2(n_283),
.B(n_210),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_941),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_899),
.A2(n_287),
.B(n_212),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_984),
.B(n_372),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1019),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1077),
.A2(n_256),
.B1(n_272),
.B2(n_381),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_933),
.A2(n_375),
.B(n_12),
.C(n_13),
.Y(n_1158)
);

AOI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_960),
.A2(n_1045),
.B(n_963),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_961),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_914),
.A2(n_256),
.B1(n_272),
.B2(n_380),
.Y(n_1161)
);

NAND2x1_ASAP7_75t_L g1162 ( 
.A(n_1018),
.B(n_486),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_984),
.B(n_11),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_899),
.A2(n_274),
.B(n_215),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_989),
.A2(n_272),
.B1(n_209),
.B2(n_379),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1029),
.A2(n_278),
.B(n_220),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_902),
.B(n_12),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_L g1168 ( 
.A(n_1050),
.B(n_364),
.C(n_252),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_989),
.A2(n_272),
.B1(n_217),
.B2(n_356),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_R g1170 ( 
.A(n_907),
.B(n_221),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1031),
.A2(n_272),
.B1(n_225),
.B2(n_355),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_961),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1014),
.B(n_272),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1049),
.Y(n_1174)
);

OAI22x1_ASAP7_75t_L g1175 ( 
.A1(n_960),
.A2(n_234),
.B1(n_230),
.B2(n_228),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1014),
.B(n_14),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1030),
.A2(n_300),
.B(n_250),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_968),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1002),
.B(n_15),
.Y(n_1179)
);

OR2x6_ASAP7_75t_SL g1180 ( 
.A(n_1017),
.B(n_227),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_974),
.A2(n_1046),
.B1(n_1069),
.B2(n_907),
.Y(n_1181)
);

OR2x6_ASAP7_75t_SL g1182 ( 
.A(n_971),
.B(n_255),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_964),
.B(n_489),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1047),
.B(n_15),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1031),
.A2(n_310),
.B1(n_260),
.B2(n_353),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1018),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_957),
.B(n_17),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_976),
.A2(n_489),
.B(n_486),
.C(n_352),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1010),
.B(n_17),
.Y(n_1189)
);

NOR3xp33_ASAP7_75t_L g1190 ( 
.A(n_1001),
.B(n_1005),
.C(n_937),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_980),
.A2(n_302),
.B(n_265),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_973),
.A2(n_312),
.B(n_266),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_947),
.A2(n_316),
.B(n_288),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_993),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1061),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_975),
.B(n_19),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1051),
.B(n_20),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_952),
.A2(n_315),
.B1(n_269),
.B2(n_347),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_976),
.A2(n_296),
.B1(n_292),
.B2(n_342),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_993),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_949),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_970),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1079),
.A2(n_489),
.B1(n_486),
.B2(n_259),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1057),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_SL g1205 ( 
.A(n_1034),
.B(n_338),
.C(n_24),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_921),
.Y(n_1206)
);

CKINVDCx11_ASAP7_75t_R g1207 ( 
.A(n_1070),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_995),
.A2(n_259),
.B(n_249),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1053),
.B(n_22),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_927),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_992),
.B(n_1036),
.Y(n_1211)
);

NOR3xp33_ASAP7_75t_SL g1212 ( 
.A(n_934),
.B(n_26),
.C(n_27),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1023),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_991),
.A2(n_28),
.B(n_34),
.C(n_38),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_977),
.A2(n_489),
.B1(n_486),
.B2(n_259),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_L g1216 ( 
.A(n_934),
.B(n_489),
.C(n_486),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1011),
.B(n_34),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1073),
.B(n_1072),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_991),
.A2(n_39),
.B(n_40),
.C(n_43),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1023),
.B(n_40),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1070),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1013),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_987),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1080),
.B(n_44),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1035),
.Y(n_1225)
);

O2A1O1Ixp5_ASAP7_75t_SL g1226 ( 
.A1(n_998),
.A2(n_919),
.B(n_1076),
.C(n_922),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1056),
.A2(n_489),
.B(n_486),
.C(n_259),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1080),
.B(n_489),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_939),
.A2(n_259),
.B(n_249),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1028),
.B(n_45),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1028),
.A2(n_47),
.B(n_48),
.C(n_51),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_949),
.B(n_47),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_958),
.A2(n_489),
.B1(n_486),
.B2(n_259),
.Y(n_1233)
);

AOI221xp5_ASAP7_75t_L g1234 ( 
.A1(n_1062),
.A2(n_489),
.B1(n_486),
.B2(n_249),
.C(n_62),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1037),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_987),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1043),
.Y(n_1237)
);

O2A1O1Ixp5_ASAP7_75t_SL g1238 ( 
.A1(n_1076),
.A2(n_986),
.B(n_939),
.C(n_972),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_958),
.B(n_48),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1188),
.A2(n_1024),
.A3(n_1008),
.B(n_1026),
.Y(n_1240)
);

BUFx4f_ASAP7_75t_L g1241 ( 
.A(n_1223),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1110),
.A2(n_1015),
.B(n_912),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1093),
.A2(n_1062),
.B(n_1056),
.C(n_1068),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1147),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1083),
.A2(n_986),
.B(n_1025),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1083),
.A2(n_1027),
.B(n_997),
.Y(n_1246)
);

BUFx8_ASAP7_75t_L g1247 ( 
.A(n_1086),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1105),
.A2(n_1007),
.B(n_1006),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1238),
.A2(n_1042),
.B(n_895),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1101),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1081),
.A2(n_1038),
.B(n_1033),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1105),
.A2(n_1048),
.B(n_1044),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_1239),
.B(n_1071),
.C(n_1012),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1149),
.B(n_1012),
.Y(n_1254)
);

AOI31xp67_ASAP7_75t_L g1255 ( 
.A1(n_1128),
.A2(n_996),
.A3(n_1075),
.B(n_994),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1156),
.Y(n_1256)
);

O2A1O1Ixp5_ASAP7_75t_SL g1257 ( 
.A1(n_1128),
.A2(n_1032),
.B(n_962),
.C(n_979),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1100),
.A2(n_1020),
.A3(n_1021),
.B(n_953),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1174),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1149),
.A2(n_1074),
.B(n_1066),
.C(n_940),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1097),
.B(n_967),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1171),
.A2(n_903),
.B(n_982),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1096),
.A2(n_1040),
.B(n_889),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1118),
.A2(n_1054),
.B(n_990),
.Y(n_1264)
);

INVxp67_ASAP7_75t_SL g1265 ( 
.A(n_1134),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1223),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1130),
.A2(n_891),
.B(n_1041),
.Y(n_1267)
);

AOI221xp5_ASAP7_75t_L g1268 ( 
.A1(n_1114),
.A2(n_1065),
.B1(n_1052),
.B2(n_1055),
.C(n_1059),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1118),
.A2(n_944),
.B(n_925),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1082),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1084),
.B(n_927),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1207),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1117),
.B(n_967),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1090),
.A2(n_1058),
.B1(n_950),
.B2(n_951),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1227),
.A2(n_1063),
.A3(n_943),
.B(n_924),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1223),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1095),
.A2(n_1136),
.B(n_1226),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1097),
.B(n_1137),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1190),
.A2(n_918),
.B(n_1064),
.Y(n_1279)
);

AOI21xp33_ASAP7_75t_L g1280 ( 
.A1(n_1239),
.A2(n_249),
.B(n_54),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1208),
.A2(n_249),
.A3(n_101),
.B(n_103),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1089),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1133),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1212),
.B(n_52),
.C(n_54),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1223),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1134),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1211),
.A2(n_104),
.A3(n_175),
.B(n_174),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1190),
.A2(n_87),
.B(n_163),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1102),
.A2(n_86),
.B(n_161),
.Y(n_1289)
);

NOR4xp25_ASAP7_75t_L g1290 ( 
.A(n_1222),
.B(n_62),
.C(n_63),
.D(n_66),
.Y(n_1290)
);

OAI22x1_ASAP7_75t_L g1291 ( 
.A1(n_1167),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1229),
.A2(n_116),
.B(n_156),
.Y(n_1292)
);

AOI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1127),
.A2(n_106),
.B(n_146),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1085),
.B(n_72),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1216),
.A2(n_93),
.B(n_137),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1201),
.B(n_72),
.Y(n_1296)
);

NOR3xp33_ASAP7_75t_L g1297 ( 
.A(n_1121),
.B(n_75),
.C(n_77),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1196),
.A2(n_75),
.B(n_77),
.C(n_85),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1201),
.B(n_133),
.Y(n_1299)
);

O2A1O1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1126),
.A2(n_136),
.B(n_189),
.C(n_1102),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1161),
.A2(n_1215),
.A3(n_1108),
.B(n_1200),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1196),
.A2(n_1125),
.B(n_1167),
.C(n_1168),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1087),
.B(n_1141),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1172),
.B(n_1119),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1195),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1091),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1109),
.Y(n_1307)
);

AO21x1_ASAP7_75t_L g1308 ( 
.A1(n_1185),
.A2(n_1193),
.B(n_1187),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1148),
.B(n_1094),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1235),
.A2(n_1237),
.A3(n_1140),
.B(n_1160),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1168),
.A2(n_1234),
.B(n_1106),
.C(n_1158),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1139),
.A2(n_1176),
.B1(n_1131),
.B2(n_1142),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_SL g1313 ( 
.A(n_1117),
.B(n_1123),
.Y(n_1313)
);

NAND3xp33_ASAP7_75t_L g1314 ( 
.A(n_1212),
.B(n_1219),
.C(n_1214),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1104),
.A2(n_1092),
.B(n_1218),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1107),
.A2(n_1103),
.B(n_1217),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1131),
.B(n_1113),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_SL g1318 ( 
.A1(n_1230),
.A2(n_1232),
.B(n_1225),
.C(n_1231),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_L g1319 ( 
.A(n_1181),
.B(n_1169),
.C(n_1165),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1189),
.A2(n_1132),
.B(n_1159),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1119),
.A2(n_1150),
.B(n_1151),
.C(n_1129),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1132),
.A2(n_1162),
.B(n_1191),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1143),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1139),
.A2(n_1163),
.B1(n_1155),
.B2(n_1182),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1153),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1113),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1178),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1135),
.A2(n_1146),
.B(n_1209),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1115),
.B(n_1124),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1172),
.B(n_1221),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1213),
.A2(n_1233),
.B(n_1203),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1194),
.A2(n_1175),
.A3(n_1224),
.B(n_1220),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1228),
.A2(n_1145),
.B(n_1144),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1221),
.B(n_1236),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1192),
.A2(n_1152),
.A3(n_1154),
.B(n_1164),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1116),
.A2(n_1205),
.B(n_1197),
.C(n_1184),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1236),
.B(n_1115),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1179),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1213),
.A2(n_1166),
.B(n_1177),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1111),
.A2(n_1157),
.B(n_1203),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1236),
.B(n_1117),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1111),
.A2(n_1088),
.B(n_1120),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_SL g1343 ( 
.A1(n_1231),
.A2(n_1210),
.B(n_1206),
.C(n_1144),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1116),
.A2(n_1117),
.B1(n_1157),
.B2(n_1236),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1088),
.A2(n_1099),
.B(n_1120),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1186),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1112),
.A2(n_1199),
.B1(n_1173),
.B2(n_1147),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1183),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_SL g1349 ( 
.A1(n_1124),
.A2(n_1198),
.B(n_1145),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1088),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1099),
.B(n_1120),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1099),
.B(n_1138),
.Y(n_1352)
);

AO21x2_ASAP7_75t_L g1353 ( 
.A1(n_1183),
.A2(n_1170),
.B(n_1138),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1098),
.A2(n_1170),
.B1(n_1204),
.B2(n_1202),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1138),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1138),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1122),
.A2(n_1180),
.B(n_1110),
.Y(n_1357)
);

NAND3x1_ASAP7_75t_L g1358 ( 
.A(n_1163),
.B(n_1090),
.C(n_718),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1110),
.A2(n_1000),
.B(n_1083),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1082),
.B(n_777),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1207),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1110),
.A2(n_1000),
.B(n_1083),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1238),
.A2(n_928),
.B(n_1171),
.Y(n_1363)
);

BUFx8_ASAP7_75t_SL g1364 ( 
.A(n_1089),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1239),
.A2(n_928),
.B1(n_755),
.B2(n_718),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1110),
.A2(n_1081),
.B(n_1096),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1110),
.A2(n_1000),
.B(n_1083),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_1147),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1216),
.A2(n_1100),
.B(n_1136),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1216),
.A2(n_1100),
.B(n_1136),
.Y(n_1370)
);

AOI221x1_ASAP7_75t_L g1371 ( 
.A1(n_1171),
.A2(n_1190),
.B1(n_718),
.B2(n_1093),
.C(n_1239),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1133),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1238),
.A2(n_928),
.B(n_1171),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1110),
.A2(n_1000),
.B(n_1083),
.Y(n_1374)
);

CKINVDCx11_ASAP7_75t_R g1375 ( 
.A(n_1180),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1238),
.A2(n_928),
.B(n_1171),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1207),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1149),
.B(n_1004),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1101),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1147),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1101),
.Y(n_1381)
);

NAND3x1_ASAP7_75t_L g1382 ( 
.A(n_1163),
.B(n_1090),
.C(n_718),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1149),
.B(n_1004),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1110),
.A2(n_1081),
.B(n_1096),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1110),
.A2(n_1000),
.B(n_1083),
.Y(n_1385)
);

OAI22x1_ASAP7_75t_L g1386 ( 
.A1(n_1090),
.A2(n_683),
.B1(n_718),
.B2(n_636),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_SL g1387 ( 
.A1(n_1102),
.A2(n_894),
.B(n_928),
.C(n_896),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1119),
.B(n_894),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1149),
.B(n_1004),
.Y(n_1389)
);

CKINVDCx14_ASAP7_75t_R g1390 ( 
.A(n_1147),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1110),
.A2(n_1000),
.B(n_1083),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1149),
.B(n_1004),
.Y(n_1392)
);

OAI221xp5_ASAP7_75t_L g1393 ( 
.A1(n_1114),
.A2(n_777),
.B1(n_773),
.B2(n_718),
.C(n_915),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1110),
.A2(n_1081),
.B(n_1096),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1082),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1101),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1082),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1101),
.Y(n_1398)
);

AOI221x1_ASAP7_75t_L g1399 ( 
.A1(n_1171),
.A2(n_1190),
.B1(n_718),
.B2(n_1093),
.C(n_1239),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1110),
.A2(n_1081),
.B(n_1096),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1101),
.Y(n_1401)
);

O2A1O1Ixp5_ASAP7_75t_L g1402 ( 
.A1(n_1171),
.A2(n_894),
.B(n_718),
.C(n_1239),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1110),
.A2(n_1081),
.B(n_1096),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1304),
.Y(n_1404)
);

BUFx4_ASAP7_75t_SL g1405 ( 
.A(n_1283),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1282),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1365),
.A2(n_1312),
.B1(n_1386),
.B2(n_1297),
.Y(n_1407)
);

CKINVDCx11_ASAP7_75t_R g1408 ( 
.A(n_1244),
.Y(n_1408)
);

INVx6_ASAP7_75t_L g1409 ( 
.A(n_1247),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1304),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1241),
.Y(n_1411)
);

BUFx12f_ASAP7_75t_L g1412 ( 
.A(n_1375),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1395),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1365),
.A2(n_1393),
.B1(n_1302),
.B2(n_1314),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1319),
.A2(n_1344),
.B1(n_1284),
.B2(n_1278),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1358),
.A2(n_1382),
.B1(n_1309),
.B2(n_1347),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1344),
.A2(n_1278),
.B1(n_1340),
.B2(n_1392),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1291),
.A2(n_1280),
.B1(n_1303),
.B2(n_1324),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1378),
.B(n_1383),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1273),
.Y(n_1420)
);

BUFx8_ASAP7_75t_SL g1421 ( 
.A(n_1372),
.Y(n_1421)
);

BUFx12f_ASAP7_75t_L g1422 ( 
.A(n_1272),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1361),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1256),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1259),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1241),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1273),
.Y(n_1427)
);

INVx4_ASAP7_75t_SL g1428 ( 
.A(n_1350),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1340),
.A2(n_1378),
.B1(n_1389),
.B2(n_1383),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1389),
.A2(n_1392),
.B1(n_1317),
.B2(n_1380),
.Y(n_1430)
);

BUFx4_ASAP7_75t_SL g1431 ( 
.A(n_1368),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1350),
.Y(n_1432)
);

BUFx12f_ASAP7_75t_L g1433 ( 
.A(n_1377),
.Y(n_1433)
);

CKINVDCx11_ASAP7_75t_R g1434 ( 
.A(n_1270),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1397),
.A2(n_1254),
.B1(n_1336),
.B2(n_1308),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1397),
.Y(n_1436)
);

INVx6_ASAP7_75t_L g1437 ( 
.A(n_1356),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1326),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1379),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1402),
.B(n_1254),
.Y(n_1440)
);

BUFx2_ASAP7_75t_SL g1441 ( 
.A(n_1266),
.Y(n_1441)
);

CKINVDCx11_ASAP7_75t_R g1442 ( 
.A(n_1390),
.Y(n_1442)
);

CKINVDCx6p67_ASAP7_75t_R g1443 ( 
.A(n_1360),
.Y(n_1443)
);

CKINVDCx11_ASAP7_75t_R g1444 ( 
.A(n_1364),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1286),
.B(n_1296),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1350),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1381),
.Y(n_1447)
);

BUFx8_ASAP7_75t_SL g1448 ( 
.A(n_1266),
.Y(n_1448)
);

OAI21xp33_ASAP7_75t_L g1449 ( 
.A1(n_1280),
.A2(n_1290),
.B(n_1298),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1296),
.A2(n_1311),
.B1(n_1253),
.B2(n_1388),
.Y(n_1450)
);

CKINVDCx6p67_ASAP7_75t_R g1451 ( 
.A(n_1356),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1313),
.A2(n_1363),
.B1(n_1373),
.B2(n_1376),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1371),
.A2(n_1399),
.B1(n_1294),
.B2(n_1338),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1271),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1313),
.A2(n_1363),
.B1(n_1373),
.B2(n_1376),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1396),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1341),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1299),
.A2(n_1294),
.B1(n_1261),
.B2(n_1346),
.Y(n_1458)
);

NAND2x1p5_ASAP7_75t_L g1459 ( 
.A(n_1276),
.B(n_1285),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1398),
.B(n_1401),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1305),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1330),
.A2(n_1323),
.B1(n_1306),
.B2(n_1325),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1354),
.A2(n_1265),
.B1(n_1329),
.B2(n_1353),
.Y(n_1463)
);

INVx6_ASAP7_75t_L g1464 ( 
.A(n_1341),
.Y(n_1464)
);

INVxp67_ASAP7_75t_SL g1465 ( 
.A(n_1330),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1276),
.B(n_1285),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1353),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1337),
.A2(n_1299),
.B1(n_1261),
.B2(n_1348),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1357),
.A2(n_1295),
.B1(n_1288),
.B2(n_1331),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1307),
.A2(n_1327),
.B1(n_1268),
.B2(n_1370),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1295),
.A2(n_1370),
.B1(n_1369),
.B2(n_1349),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1369),
.A2(n_1334),
.B1(n_1320),
.B2(n_1274),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1337),
.A2(n_1334),
.B1(n_1321),
.B2(n_1387),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1310),
.Y(n_1474)
);

BUFx10_ASAP7_75t_L g1475 ( 
.A(n_1343),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_SL g1476 ( 
.A1(n_1262),
.A2(n_1316),
.B1(n_1289),
.B2(n_1328),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1262),
.A2(n_1249),
.B1(n_1248),
.B2(n_1342),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1355),
.B(n_1332),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1243),
.A2(n_1260),
.B1(n_1300),
.B2(n_1245),
.Y(n_1479)
);

CKINVDCx11_ASAP7_75t_R g1480 ( 
.A(n_1332),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1310),
.Y(n_1481)
);

BUFx4f_ASAP7_75t_L g1482 ( 
.A(n_1351),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_1351),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1352),
.Y(n_1484)
);

CKINVDCx6p67_ASAP7_75t_R g1485 ( 
.A(n_1352),
.Y(n_1485)
);

INVx6_ASAP7_75t_L g1486 ( 
.A(n_1345),
.Y(n_1486)
);

OAI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1246),
.A2(n_1279),
.B1(n_1315),
.B2(n_1362),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1333),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1287),
.Y(n_1489)
);

CKINVDCx12_ASAP7_75t_R g1490 ( 
.A(n_1287),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1335),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1359),
.A2(n_1367),
.B(n_1374),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1318),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1249),
.A2(n_1269),
.B1(n_1277),
.B2(n_1322),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1264),
.Y(n_1495)
);

OAI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1385),
.A2(n_1391),
.B1(n_1252),
.B2(n_1339),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1293),
.A2(n_1257),
.B1(n_1255),
.B2(n_1240),
.Y(n_1497)
);

BUFx4_ASAP7_75t_R g1498 ( 
.A(n_1258),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1292),
.A2(n_1242),
.B1(n_1263),
.B2(n_1267),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1281),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1251),
.A2(n_1366),
.B1(n_1400),
.B2(n_1394),
.Y(n_1501)
);

CKINVDCx11_ASAP7_75t_R g1502 ( 
.A(n_1281),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1281),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1258),
.Y(n_1504)
);

CKINVDCx9p33_ASAP7_75t_R g1505 ( 
.A(n_1258),
.Y(n_1505)
);

BUFx2_ASAP7_75t_SL g1506 ( 
.A(n_1275),
.Y(n_1506)
);

INVx6_ASAP7_75t_L g1507 ( 
.A(n_1275),
.Y(n_1507)
);

CKINVDCx12_ASAP7_75t_R g1508 ( 
.A(n_1240),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1240),
.B(n_1301),
.Y(n_1509)
);

BUFx4_ASAP7_75t_R g1510 ( 
.A(n_1301),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_SL g1511 ( 
.A1(n_1301),
.A2(n_1384),
.B1(n_1403),
.B2(n_1275),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1378),
.B(n_1383),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1365),
.A2(n_566),
.B1(n_718),
.B2(n_1090),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1317),
.B(n_1309),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1282),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1365),
.A2(n_1090),
.B1(n_718),
.B2(n_814),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1364),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1250),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1365),
.A2(n_566),
.B1(n_718),
.B2(n_1090),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1378),
.B(n_1383),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1378),
.B(n_1383),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1365),
.A2(n_718),
.B1(n_1312),
.B2(n_633),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1250),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1250),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1250),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1365),
.A2(n_566),
.B1(n_718),
.B2(n_1090),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1364),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1365),
.A2(n_1090),
.B1(n_718),
.B2(n_814),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1365),
.A2(n_1402),
.B(n_718),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1250),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1317),
.B(n_1309),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1364),
.Y(n_1532)
);

BUFx12f_ASAP7_75t_L g1533 ( 
.A(n_1375),
.Y(n_1533)
);

BUFx4f_ASAP7_75t_SL g1534 ( 
.A(n_1244),
.Y(n_1534)
);

OAI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1365),
.A2(n_1312),
.B1(n_1278),
.B2(n_1284),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1364),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1364),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1364),
.Y(n_1538)
);

BUFx12f_ASAP7_75t_L g1539 ( 
.A(n_1375),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1365),
.A2(n_894),
.B1(n_1393),
.B2(n_1302),
.Y(n_1540)
);

CKINVDCx6p67_ASAP7_75t_R g1541 ( 
.A(n_1375),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1365),
.A2(n_1090),
.B1(n_718),
.B2(n_814),
.Y(n_1542)
);

CKINVDCx6p67_ASAP7_75t_R g1543 ( 
.A(n_1375),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1365),
.A2(n_1090),
.B1(n_718),
.B2(n_814),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1365),
.A2(n_1312),
.B1(n_1278),
.B2(n_1284),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1365),
.A2(n_1312),
.B1(n_1278),
.B2(n_1284),
.Y(n_1546)
);

OAI22x1_ASAP7_75t_L g1547 ( 
.A1(n_1312),
.A2(n_1338),
.B1(n_1090),
.B2(n_718),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1364),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1474),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1443),
.B(n_1436),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1419),
.B(n_1512),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1520),
.B(n_1521),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1446),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1492),
.A2(n_1479),
.B(n_1497),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1481),
.Y(n_1555)
);

AOI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1440),
.A2(n_1489),
.B(n_1493),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1513),
.A2(n_1526),
.B1(n_1519),
.B2(n_1522),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1478),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1404),
.Y(n_1559)
);

AO21x2_ASAP7_75t_L g1560 ( 
.A1(n_1503),
.A2(n_1453),
.B(n_1496),
.Y(n_1560)
);

OR2x6_ASAP7_75t_L g1561 ( 
.A(n_1467),
.B(n_1506),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1404),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1410),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1514),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1410),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1531),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1488),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1406),
.B(n_1515),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1486),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1454),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1516),
.A2(n_1544),
.B1(n_1542),
.B2(n_1528),
.Y(n_1571)
);

BUFx2_ASAP7_75t_SL g1572 ( 
.A(n_1475),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1465),
.B(n_1445),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1534),
.B(n_1434),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1509),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1486),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1439),
.B(n_1447),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1494),
.A2(n_1477),
.B(n_1499),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1534),
.B(n_1408),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1494),
.A2(n_1477),
.B(n_1499),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1456),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1461),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1518),
.Y(n_1584)
);

AOI21xp33_ASAP7_75t_L g1585 ( 
.A1(n_1547),
.A2(n_1546),
.B(n_1545),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1516),
.A2(n_1544),
.B1(n_1528),
.B2(n_1542),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1540),
.A2(n_1529),
.B(n_1414),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1495),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1501),
.A2(n_1504),
.B(n_1472),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1413),
.B(n_1438),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1428),
.B(n_1427),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1523),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1524),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1525),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1530),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1491),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1508),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1510),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1510),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1452),
.B(n_1455),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1429),
.B(n_1417),
.Y(n_1601)
);

BUFx4f_ASAP7_75t_SL g1602 ( 
.A(n_1532),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1502),
.A2(n_1407),
.B1(n_1535),
.B2(n_1546),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1460),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1507),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1500),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1407),
.A2(n_1545),
.B1(n_1535),
.B2(n_1449),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1490),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1507),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1507),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1498),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1472),
.B(n_1484),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1498),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1473),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1430),
.B(n_1435),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1440),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1505),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1468),
.B(n_1458),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1505),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1466),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1462),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1432),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1457),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1462),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1487),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1480),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1450),
.A2(n_1415),
.B(n_1453),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1464),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1464),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1416),
.B(n_1418),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1475),
.Y(n_1631)
);

AO21x2_ASAP7_75t_L g1632 ( 
.A1(n_1496),
.A2(n_1487),
.B(n_1463),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1511),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1432),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1470),
.A2(n_1459),
.B(n_1427),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1448),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1459),
.A2(n_1476),
.B(n_1469),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1464),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1485),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1471),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1432),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1432),
.Y(n_1642)
);

AND2x4_ASAP7_75t_SL g1643 ( 
.A(n_1483),
.B(n_1451),
.Y(n_1643)
);

AOI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1441),
.A2(n_1437),
.B(n_1418),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1482),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1411),
.B(n_1426),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1482),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1431),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1437),
.A2(n_1420),
.B(n_1411),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1426),
.A2(n_1409),
.B(n_1541),
.C(n_1543),
.Y(n_1650)
);

CKINVDCx12_ASAP7_75t_R g1651 ( 
.A(n_1405),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1409),
.Y(n_1652)
);

INVxp33_ASAP7_75t_SL g1653 ( 
.A(n_1517),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1422),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1423),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1412),
.A2(n_1533),
.B1(n_1539),
.B2(n_1442),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1433),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1527),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1537),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1536),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1444),
.B(n_1538),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1559),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1587),
.A2(n_1548),
.B(n_1421),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1564),
.B(n_1566),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1562),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1551),
.B(n_1552),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1627),
.A2(n_1557),
.B1(n_1585),
.B2(n_1601),
.C(n_1615),
.Y(n_1667)
);

A2O1A1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1557),
.A2(n_1600),
.B(n_1603),
.C(n_1618),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1605),
.B(n_1611),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1588),
.B(n_1620),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1588),
.B(n_1618),
.Y(n_1671)
);

BUFx4f_ASAP7_75t_SL g1672 ( 
.A(n_1659),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1588),
.B(n_1576),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1607),
.A2(n_1586),
.B1(n_1571),
.B2(n_1600),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1630),
.A2(n_1614),
.B1(n_1615),
.B2(n_1572),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1632),
.A2(n_1625),
.B(n_1554),
.Y(n_1676)
);

AO32x2_ASAP7_75t_L g1677 ( 
.A1(n_1573),
.A2(n_1575),
.A3(n_1565),
.B1(n_1563),
.B2(n_1562),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_SL g1678 ( 
.A(n_1572),
.B(n_1632),
.Y(n_1678)
);

OAI211xp5_ASAP7_75t_L g1679 ( 
.A1(n_1625),
.A2(n_1630),
.B(n_1616),
.C(n_1633),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1614),
.A2(n_1554),
.B(n_1616),
.Y(n_1680)
);

O2A1O1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1633),
.A2(n_1640),
.B(n_1590),
.C(n_1631),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1632),
.B(n_1576),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1568),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1570),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1579),
.A2(n_1581),
.B(n_1637),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1579),
.A2(n_1581),
.B(n_1589),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1591),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1578),
.B(n_1643),
.Y(n_1688)
);

O2A1O1Ixp33_ASAP7_75t_SL g1689 ( 
.A1(n_1650),
.A2(n_1631),
.B(n_1658),
.C(n_1660),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1553),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1560),
.A2(n_1569),
.B(n_1577),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1644),
.A2(n_1556),
.B(n_1635),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1584),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1622),
.B(n_1634),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1621),
.A2(n_1624),
.B1(n_1604),
.B2(n_1593),
.C(n_1595),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1592),
.B(n_1593),
.Y(n_1698)
);

OAI21xp33_ASAP7_75t_SL g1699 ( 
.A1(n_1652),
.A2(n_1550),
.B(n_1647),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_SL g1700 ( 
.A1(n_1658),
.A2(n_1660),
.B(n_1653),
.C(n_1580),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1644),
.A2(n_1635),
.B(n_1577),
.Y(n_1701)
);

NAND4xp25_ASAP7_75t_L g1702 ( 
.A(n_1656),
.B(n_1574),
.C(n_1595),
.D(n_1594),
.Y(n_1702)
);

OA21x2_ASAP7_75t_L g1703 ( 
.A1(n_1606),
.A2(n_1617),
.B(n_1619),
.Y(n_1703)
);

BUFx12f_ASAP7_75t_L g1704 ( 
.A(n_1648),
.Y(n_1704)
);

AND4x1_ASAP7_75t_L g1705 ( 
.A(n_1661),
.B(n_1651),
.C(n_1657),
.D(n_1654),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1648),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1623),
.B(n_1639),
.Y(n_1707)
);

A2O1A1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1598),
.A2(n_1599),
.B(n_1613),
.C(n_1621),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1549),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1598),
.A2(n_1599),
.B(n_1624),
.C(n_1612),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1549),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1641),
.Y(n_1712)
);

BUFx12f_ASAP7_75t_L g1713 ( 
.A(n_1553),
.Y(n_1713)
);

AO32x2_ASAP7_75t_L g1714 ( 
.A1(n_1575),
.A2(n_1558),
.A3(n_1628),
.B1(n_1638),
.B2(n_1629),
.Y(n_1714)
);

CKINVDCx6p67_ASAP7_75t_R g1715 ( 
.A(n_1651),
.Y(n_1715)
);

OR2x6_ASAP7_75t_L g1716 ( 
.A(n_1561),
.B(n_1608),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1605),
.B(n_1608),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1553),
.B(n_1626),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1558),
.B(n_1638),
.Y(n_1719)
);

NOR2xp67_ASAP7_75t_L g1720 ( 
.A(n_1699),
.B(n_1629),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1709),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1711),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1671),
.B(n_1567),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1712),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1673),
.B(n_1641),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1665),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1715),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1667),
.A2(n_1597),
.B1(n_1610),
.B2(n_1609),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1682),
.B(n_1561),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1677),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1671),
.B(n_1666),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1682),
.B(n_1642),
.Y(n_1732)
);

NOR2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1715),
.B(n_1636),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1695),
.Y(n_1734)
);

CKINVDCx6p67_ASAP7_75t_R g1735 ( 
.A(n_1704),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1692),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1670),
.B(n_1596),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1662),
.B(n_1692),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1694),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1696),
.B(n_1596),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1677),
.B(n_1609),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1677),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1677),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1698),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1668),
.A2(n_1645),
.B1(n_1646),
.B2(n_1636),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1668),
.A2(n_1646),
.B1(n_1655),
.B2(n_1657),
.Y(n_1746)
);

INVx4_ASAP7_75t_L g1747 ( 
.A(n_1713),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1703),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1719),
.B(n_1555),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1714),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1714),
.Y(n_1751)
);

INVxp67_ASAP7_75t_SL g1752 ( 
.A(n_1703),
.Y(n_1752)
);

OR2x6_ASAP7_75t_L g1753 ( 
.A(n_1716),
.B(n_1649),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1730),
.B(n_1685),
.Y(n_1754)
);

NOR2xp67_ASAP7_75t_L g1755 ( 
.A(n_1729),
.B(n_1676),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1721),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1721),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1750),
.Y(n_1758)
);

BUFx2_ASAP7_75t_L g1759 ( 
.A(n_1752),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1730),
.B(n_1703),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1748),
.B(n_1736),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1748),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1736),
.B(n_1680),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1745),
.A2(n_1674),
.B1(n_1675),
.B2(n_1679),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1746),
.A2(n_1710),
.B1(n_1708),
.B2(n_1683),
.Y(n_1765)
);

AOI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1742),
.A2(n_1681),
.B1(n_1697),
.B2(n_1710),
.C(n_1702),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1742),
.B(n_1678),
.Y(n_1767)
);

OR2x6_ASAP7_75t_L g1768 ( 
.A(n_1753),
.B(n_1701),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1750),
.B(n_1686),
.Y(n_1769)
);

OAI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1728),
.A2(n_1708),
.B1(n_1705),
.B2(n_1689),
.C(n_1707),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1751),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1743),
.B(n_1691),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1722),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1739),
.B(n_1714),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1741),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1722),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1720),
.B(n_1687),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1733),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1744),
.B(n_1664),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1729),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1732),
.B(n_1688),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1725),
.B(n_1669),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1725),
.B(n_1669),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1778),
.B(n_1735),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1763),
.B(n_1726),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1759),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1759),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1756),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1772),
.B(n_1731),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1782),
.B(n_1783),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1756),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1757),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1763),
.B(n_1726),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1758),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1775),
.B(n_1724),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1772),
.B(n_1738),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1757),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1773),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1778),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1775),
.B(n_1723),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1773),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1780),
.B(n_1720),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1774),
.B(n_1737),
.Y(n_1803)
);

NOR3xp33_ASAP7_75t_L g1804 ( 
.A(n_1764),
.B(n_1689),
.C(n_1663),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1776),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1776),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1780),
.B(n_1755),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1763),
.B(n_1734),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1783),
.B(n_1737),
.Y(n_1809)
);

NAND4xp25_ASAP7_75t_L g1810 ( 
.A(n_1759),
.B(n_1700),
.C(n_1727),
.D(n_1684),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1774),
.B(n_1740),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1754),
.B(n_1734),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1764),
.A2(n_1693),
.B1(n_1717),
.B2(n_1753),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1774),
.B(n_1740),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1779),
.B(n_1749),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1762),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1779),
.B(n_1754),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1789),
.B(n_1771),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1816),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1788),
.Y(n_1820)
);

INVxp67_ASAP7_75t_SL g1821 ( 
.A(n_1804),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1789),
.B(n_1771),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1788),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1791),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1786),
.Y(n_1825)
);

OAI21xp33_ASAP7_75t_L g1826 ( 
.A1(n_1804),
.A2(n_1762),
.B(n_1766),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1816),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1796),
.B(n_1754),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1802),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1786),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1796),
.B(n_1771),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1802),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1817),
.B(n_1771),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1785),
.B(n_1793),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1791),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1792),
.Y(n_1836)
);

AOI211xp5_ASAP7_75t_L g1837 ( 
.A1(n_1810),
.A2(n_1770),
.B(n_1765),
.C(n_1766),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1790),
.B(n_1778),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1785),
.B(n_1760),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1786),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1792),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1790),
.B(n_1783),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1797),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1811),
.B(n_1761),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1784),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1802),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1802),
.B(n_1760),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1817),
.B(n_1769),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1811),
.B(n_1761),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1794),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1811),
.B(n_1761),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1793),
.B(n_1769),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1799),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1797),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1798),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1814),
.B(n_1781),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1798),
.Y(n_1857)
);

AOI21xp33_ASAP7_75t_L g1858 ( 
.A1(n_1813),
.A2(n_1770),
.B(n_1765),
.Y(n_1858)
);

INVxp33_ASAP7_75t_L g1859 ( 
.A(n_1810),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1808),
.B(n_1760),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1799),
.B(n_1777),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1808),
.B(n_1812),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1801),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1834),
.B(n_1812),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1820),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1820),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1826),
.B(n_1794),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1856),
.B(n_1799),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1862),
.B(n_1815),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1862),
.B(n_1815),
.Y(n_1870)
);

AOI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1826),
.A2(n_1762),
.B1(n_1758),
.B2(n_1816),
.C(n_1787),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1821),
.B(n_1801),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1819),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1837),
.B(n_1805),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1828),
.B(n_1800),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1856),
.B(n_1814),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1842),
.B(n_1814),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1819),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1850),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1818),
.B(n_1800),
.Y(n_1880)
);

INVx2_ASAP7_75t_SL g1881 ( 
.A(n_1829),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1837),
.B(n_1807),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1823),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1823),
.B(n_1805),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1842),
.B(n_1803),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1827),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1844),
.B(n_1849),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1827),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1824),
.B(n_1806),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1824),
.Y(n_1890)
);

INVxp67_ASAP7_75t_L g1891 ( 
.A(n_1853),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1835),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1833),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1844),
.B(n_1803),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1833),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1849),
.B(n_1803),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1838),
.B(n_1809),
.Y(n_1897)
);

NAND4xp25_ASAP7_75t_L g1898 ( 
.A(n_1858),
.B(n_1787),
.C(n_1700),
.D(n_1727),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1847),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1845),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1874),
.B(n_1859),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1865),
.Y(n_1902)
);

AOI32xp33_ASAP7_75t_L g1903 ( 
.A1(n_1874),
.A2(n_1847),
.A3(n_1839),
.B1(n_1860),
.B2(n_1848),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1865),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1897),
.B(n_1838),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1882),
.A2(n_1847),
.B1(n_1768),
.B2(n_1762),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1866),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1867),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1866),
.Y(n_1909)
);

INVx2_ASAP7_75t_SL g1910 ( 
.A(n_1868),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1897),
.B(n_1851),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1900),
.B(n_1851),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_1900),
.Y(n_1913)
);

NOR4xp25_ASAP7_75t_L g1914 ( 
.A(n_1867),
.B(n_1840),
.C(n_1830),
.D(n_1825),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1883),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1879),
.B(n_1818),
.Y(n_1916)
);

OAI21xp33_ASAP7_75t_L g1917 ( 
.A1(n_1898),
.A2(n_1847),
.B(n_1848),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1869),
.B(n_1822),
.Y(n_1918)
);

AOI211xp5_ASAP7_75t_L g1919 ( 
.A1(n_1871),
.A2(n_1846),
.B(n_1829),
.C(n_1832),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1879),
.B(n_1822),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1883),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1871),
.A2(n_1861),
.B1(n_1846),
.B2(n_1832),
.Y(n_1922)
);

AOI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1898),
.A2(n_1755),
.B1(n_1768),
.B2(n_1807),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1890),
.Y(n_1924)
);

OAI31xp33_ASAP7_75t_L g1925 ( 
.A1(n_1872),
.A2(n_1899),
.A3(n_1893),
.B(n_1895),
.Y(n_1925)
);

AOI221xp5_ASAP7_75t_L g1926 ( 
.A1(n_1872),
.A2(n_1852),
.B1(n_1830),
.B2(n_1825),
.C(n_1840),
.Y(n_1926)
);

AOI21xp33_ASAP7_75t_L g1927 ( 
.A1(n_1893),
.A2(n_1830),
.B(n_1825),
.Y(n_1927)
);

INVxp67_ASAP7_75t_L g1928 ( 
.A(n_1901),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1913),
.B(n_1891),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1901),
.A2(n_1891),
.B(n_1881),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1905),
.B(n_1887),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1902),
.Y(n_1932)
);

O2A1O1Ixp33_ASAP7_75t_L g1933 ( 
.A1(n_1908),
.A2(n_1881),
.B(n_1890),
.C(n_1892),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1904),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1914),
.A2(n_1899),
.B1(n_1893),
.B2(n_1895),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1907),
.Y(n_1936)
);

OAI21xp33_ASAP7_75t_L g1937 ( 
.A1(n_1917),
.A2(n_1899),
.B(n_1868),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1909),
.Y(n_1938)
);

OAI21xp33_ASAP7_75t_L g1939 ( 
.A1(n_1903),
.A2(n_1868),
.B(n_1875),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1915),
.Y(n_1940)
);

OAI311xp33_ASAP7_75t_L g1941 ( 
.A1(n_1906),
.A2(n_1869),
.A3(n_1870),
.B1(n_1875),
.C1(n_1887),
.Y(n_1941)
);

OAI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1923),
.A2(n_1868),
.B1(n_1887),
.B2(n_1885),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1906),
.A2(n_1877),
.B1(n_1885),
.B2(n_1870),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1908),
.A2(n_1768),
.B1(n_1888),
.B2(n_1886),
.Y(n_1944)
);

HB1xp67_ASAP7_75t_L g1945 ( 
.A(n_1916),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1921),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1922),
.A2(n_1895),
.B1(n_1888),
.B2(n_1886),
.Y(n_1947)
);

OAI211xp5_ASAP7_75t_SL g1948 ( 
.A1(n_1925),
.A2(n_1919),
.B(n_1912),
.C(n_1926),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1931),
.Y(n_1949)
);

XOR2x2_ASAP7_75t_L g1950 ( 
.A(n_1930),
.B(n_1661),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1928),
.Y(n_1951)
);

OAI322xp33_ASAP7_75t_L g1952 ( 
.A1(n_1928),
.A2(n_1920),
.A3(n_1918),
.B1(n_1924),
.B2(n_1910),
.C1(n_1881),
.C2(n_1892),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1947),
.A2(n_1910),
.B1(n_1905),
.B2(n_1911),
.Y(n_1953)
);

OAI322xp33_ASAP7_75t_L g1954 ( 
.A1(n_1929),
.A2(n_1935),
.A3(n_1945),
.B1(n_1933),
.B2(n_1932),
.C1(n_1936),
.C2(n_1946),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1945),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1939),
.B(n_1911),
.Y(n_1956)
);

XNOR2x1_ASAP7_75t_L g1957 ( 
.A(n_1943),
.B(n_1733),
.Y(n_1957)
);

XNOR2xp5_ASAP7_75t_L g1958 ( 
.A(n_1942),
.B(n_1706),
.Y(n_1958)
);

OAI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1948),
.A2(n_1927),
.B1(n_1829),
.B2(n_1832),
.C(n_1846),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1937),
.B(n_1602),
.Y(n_1960)
);

INVx2_ASAP7_75t_SL g1961 ( 
.A(n_1934),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1951),
.B(n_1952),
.Y(n_1962)
);

NAND4xp25_ASAP7_75t_L g1963 ( 
.A(n_1956),
.B(n_1940),
.C(n_1938),
.D(n_1941),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1955),
.B(n_1877),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1961),
.Y(n_1965)
);

NAND3xp33_ASAP7_75t_SL g1966 ( 
.A(n_1959),
.B(n_1944),
.C(n_1896),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1950),
.Y(n_1967)
);

NOR3xp33_ASAP7_75t_SL g1968 ( 
.A(n_1954),
.B(n_1706),
.C(n_1884),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1958),
.B(n_1829),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1949),
.B(n_1877),
.Y(n_1970)
);

NOR3xp33_ASAP7_75t_L g1971 ( 
.A(n_1954),
.B(n_1953),
.C(n_1960),
.Y(n_1971)
);

NOR2x1_ASAP7_75t_L g1972 ( 
.A(n_1957),
.B(n_1659),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1964),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1971),
.B(n_1894),
.Y(n_1974)
);

AOI222xp33_ASAP7_75t_L g1975 ( 
.A1(n_1962),
.A2(n_1888),
.B1(n_1873),
.B2(n_1886),
.C1(n_1878),
.C2(n_1840),
.Y(n_1975)
);

OAI211xp5_ASAP7_75t_L g1976 ( 
.A1(n_1963),
.A2(n_1846),
.B(n_1832),
.C(n_1896),
.Y(n_1976)
);

OAI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1968),
.A2(n_1896),
.B(n_1894),
.Y(n_1977)
);

AOI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1966),
.A2(n_1967),
.B1(n_1970),
.B2(n_1965),
.C(n_1873),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1973),
.B(n_1972),
.Y(n_1979)
);

OAI221xp5_ASAP7_75t_L g1980 ( 
.A1(n_1975),
.A2(n_1969),
.B1(n_1873),
.B2(n_1878),
.C(n_1880),
.Y(n_1980)
);

AOI221xp5_ASAP7_75t_L g1981 ( 
.A1(n_1976),
.A2(n_1878),
.B1(n_1889),
.B2(n_1884),
.C(n_1787),
.Y(n_1981)
);

AOI221xp5_ASAP7_75t_L g1982 ( 
.A1(n_1978),
.A2(n_1889),
.B1(n_1876),
.B2(n_1880),
.C(n_1894),
.Y(n_1982)
);

OAI211xp5_ASAP7_75t_L g1983 ( 
.A1(n_1974),
.A2(n_1876),
.B(n_1885),
.C(n_1864),
.Y(n_1983)
);

OAI211xp5_ASAP7_75t_SL g1984 ( 
.A1(n_1977),
.A2(n_1864),
.B(n_1654),
.C(n_1655),
.Y(n_1984)
);

NOR2x1_ASAP7_75t_L g1985 ( 
.A(n_1979),
.B(n_1876),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1983),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1980),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1984),
.A2(n_1735),
.B1(n_1704),
.B2(n_1852),
.Y(n_1988)
);

AOI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1982),
.A2(n_1718),
.B1(n_1831),
.B2(n_1807),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1985),
.B(n_1835),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1986),
.B(n_1831),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_SL g1992 ( 
.A(n_1987),
.B(n_1713),
.Y(n_1992)
);

AOI211xp5_ASAP7_75t_SL g1993 ( 
.A1(n_1991),
.A2(n_1981),
.B(n_1988),
.C(n_1989),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1993),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_1992),
.B1(n_1990),
.B2(n_1672),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1994),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1996),
.Y(n_1997)
);

OAI22x1_ASAP7_75t_L g1998 ( 
.A1(n_1995),
.A2(n_1863),
.B1(n_1857),
.B2(n_1855),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1997),
.A2(n_1863),
.B1(n_1857),
.B2(n_1855),
.Y(n_1999)
);

OAI221xp5_ASAP7_75t_SL g2000 ( 
.A1(n_1998),
.A2(n_1854),
.B1(n_1843),
.B2(n_1841),
.C(n_1836),
.Y(n_2000)
);

OAI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_2000),
.A2(n_1854),
.B(n_1843),
.Y(n_2001)
);

OAI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_2001),
.A2(n_1999),
.B(n_1841),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_2002),
.Y(n_2003)
);

OAI221xp5_ASAP7_75t_R g2004 ( 
.A1(n_2003),
.A2(n_1672),
.B1(n_1836),
.B2(n_1795),
.C(n_1747),
.Y(n_2004)
);

AOI211xp5_ASAP7_75t_L g2005 ( 
.A1(n_2004),
.A2(n_1690),
.B(n_1767),
.C(n_1807),
.Y(n_2005)
);


endmodule