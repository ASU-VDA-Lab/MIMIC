module real_jpeg_5649_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_469;
wire n_98;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_531;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_0),
.A2(n_49),
.B1(n_51),
.B2(n_57),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_0),
.A2(n_57),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_0),
.A2(n_57),
.B1(n_144),
.B2(n_148),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_0),
.A2(n_57),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_1),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_1),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_1),
.Y(n_246)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_1),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_1),
.Y(n_435)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_2),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_2),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_3),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_3),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_3),
.A2(n_77),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_3),
.A2(n_77),
.B1(n_406),
.B2(n_407),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_3),
.A2(n_77),
.B1(n_110),
.B2(n_416),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_4),
.A2(n_210),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_4),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_4),
.A2(n_290),
.B1(n_385),
.B2(n_387),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_4),
.A2(n_277),
.B1(n_290),
.B2(n_414),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_4),
.A2(n_290),
.B1(n_348),
.B2(n_469),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_6),
.A2(n_164),
.B1(n_167),
.B2(n_171),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_6),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_6),
.B(n_181),
.C(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_6),
.B(n_93),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_6),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_6),
.B(n_142),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_6),
.B(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_7),
.Y(n_545)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_8),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_52),
.B1(n_61),
.B2(n_64),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_9),
.A2(n_64),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_9),
.A2(n_64),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_9),
.A2(n_64),
.B1(n_406),
.B2(n_423),
.Y(n_422)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_11),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_11),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_12),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_12),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_12),
.A2(n_194),
.B1(n_219),
.B2(n_241),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_12),
.A2(n_219),
.B1(n_318),
.B2(n_320),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_12),
.A2(n_74),
.B1(n_219),
.B2(n_439),
.Y(n_438)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_14),
.Y(n_548)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_16),
.A2(n_188),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_16),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_16),
.A2(n_179),
.B1(n_192),
.B2(n_267),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_16),
.A2(n_109),
.B1(n_192),
.B2(n_282),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_16),
.A2(n_74),
.B1(n_76),
.B2(n_192),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_17),
.A2(n_62),
.B1(n_79),
.B2(n_81),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_17),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_17),
.A2(n_81),
.B1(n_190),
.B2(n_329),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_17),
.A2(n_81),
.B1(n_148),
.B2(n_410),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_17),
.A2(n_81),
.B1(n_453),
.B2(n_455),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_18),
.A2(n_127),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_18),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_18),
.A2(n_174),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_18),
.A2(n_104),
.B1(n_174),
.B2(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_18),
.A2(n_174),
.B1(n_374),
.B2(n_379),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_544),
.B(n_546),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_66),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_58),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_39),
.B(n_47),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_24),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_24),
.B(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_33),
.B2(n_37),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_28),
.Y(n_352)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_31),
.Y(n_456)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_32),
.Y(n_274)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_32),
.Y(n_283)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_32),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_32),
.Y(n_454)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_36),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_36),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_39),
.A2(n_373),
.B(n_376),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_39),
.B(n_378),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g350 ( 
.A(n_43),
.Y(n_350)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_58)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_56),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_58),
.B(n_69),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_65),
.B1(n_73),
.B2(n_78),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_78),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_59),
.A2(n_377),
.B(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_59),
.A2(n_65),
.B1(n_418),
.B2(n_438),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_59),
.A2(n_65),
.B1(n_73),
.B2(n_516),
.Y(n_515)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_63),
.Y(n_359)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_63),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_65),
.B(n_171),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_65),
.A2(n_438),
.B(n_470),
.Y(n_480)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_153),
.B(n_543),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_149),
.C(n_150),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_70),
.A2(n_71),
.B1(n_539),
.B2(n_540),
.Y(n_538)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_82),
.C(n_112),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_72),
.B(n_531),
.Y(n_530)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_76),
.Y(n_379)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_82),
.A2(n_112),
.B1(n_113),
.B2(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_82),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_101),
.B1(n_106),
.B2(n_107),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_83),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_83),
.A2(n_106),
.B1(n_317),
.B2(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_83),
.A2(n_106),
.B1(n_413),
.B2(n_415),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_83),
.A2(n_101),
.B1(n_106),
.B2(n_520),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_89),
.Y(n_299)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_89),
.Y(n_306)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_93),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

AOI22x1_ASAP7_75t_L g442 ( 
.A1(n_93),
.A2(n_151),
.B1(n_324),
.B2(n_443),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_93),
.A2(n_151),
.B1(n_451),
.B2(n_452),
.Y(n_450)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_99),
.Y(n_93)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_95),
.Y(n_386)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_96),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_96),
.Y(n_267)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx6_ASAP7_75t_L g425 ( 
.A(n_98),
.Y(n_425)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_106),
.B(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_106),
.A2(n_317),
.B(n_323),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g293 ( 
.A1(n_109),
.A2(n_276),
.A3(n_294),
.B1(n_296),
.B2(n_300),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_111),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_112),
.A2(n_113),
.B1(n_518),
.B2(n_519),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_112),
.B(n_515),
.C(n_518),
.Y(n_526)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_141),
.B(n_143),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_114),
.A2(n_163),
.B(n_172),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_114),
.A2(n_141),
.B1(n_217),
.B2(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_114),
.A2(n_172),
.B(n_266),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_114),
.A2(n_141),
.B1(n_384),
.B2(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_115),
.B(n_173),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_115),
.A2(n_142),
.B1(n_405),
.B2(n_409),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_115),
.A2(n_142),
.B1(n_409),
.B2(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_115),
.A2(n_142),
.B1(n_422),
.B2(n_459),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_130),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_120),
.B1(n_123),
.B2(n_127),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_131),
.B1(n_135),
.B2(n_138),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_129),
.Y(n_388)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_130),
.A2(n_217),
.B(n_223),
.Y(n_216)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_133),
.Y(n_330)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_133),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_137),
.Y(n_289)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_141),
.A2(n_223),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_142),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_143),
.Y(n_459)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_149),
.B(n_150),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_151),
.A2(n_270),
.B(n_279),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_151),
.B(n_324),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_151),
.A2(n_279),
.B(n_483),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_537),
.B(n_542),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_509),
.B(n_534),
.Y(n_154)
);

OAI311xp33_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_391),
.A3(n_485),
.B1(n_503),
.C1(n_508),
.Y(n_155)
);

AOI21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_336),
.B(n_390),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_308),
.B(n_335),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_260),
.B(n_307),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_226),
.B(n_259),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_185),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_161),
.B(n_185),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_176),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_162),
.A2(n_176),
.B1(n_177),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_162),
.Y(n_257)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_166),
.Y(n_410)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_170),
.Y(n_295)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_170),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_171),
.A2(n_198),
.B(n_205),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_SL g270 ( 
.A1(n_171),
.A2(n_271),
.B(n_275),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_171),
.B(n_357),
.Y(n_356)
);

OAI21xp33_ASAP7_75t_SL g373 ( 
.A1(n_171),
.A2(n_356),
.B(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_175),
.Y(n_406)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_214),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_186),
.B(n_215),
.C(n_225),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_198),
.B(n_205),
.Y(n_186)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_190),
.Y(n_399)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_198),
.A2(n_362),
.B1(n_363),
.B2(n_365),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_198),
.A2(n_397),
.B1(n_400),
.B2(n_401),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_198),
.A2(n_332),
.B(n_401),
.Y(n_426)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_199),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_199),
.A2(n_287),
.B1(n_328),
.B2(n_331),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_199),
.A2(n_366),
.B1(n_433),
.B2(n_434),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_213),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_224),
.B2(n_225),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_218),
.Y(n_408)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_250),
.B(n_258),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_238),
.B(n_249),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_237),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_236),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_248),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_248),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_244),
.B(n_247),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_286),
.B(n_291),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_256),
.Y(n_258)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_262),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_284),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_268),
.B2(n_269),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_268),
.C(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_293),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_293),
.Y(n_314)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_309),
.B(n_310),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_315),
.B2(n_334),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_314),
.C(n_334),
.Y(n_337)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_315),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_325),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_316),
.B(n_326),
.C(n_327),
.Y(n_367)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_329),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_331),
.Y(n_400)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx8_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_337),
.B(n_338),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_370),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_367),
.B1(n_368),
.B2(n_369),
.Y(n_339)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_340),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_360),
.B2(n_361),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_342),
.B(n_360),
.Y(n_481)
);

OAI32xp33_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_346),
.A3(n_349),
.B1(n_351),
.B2(n_356),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx8_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_367),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_367),
.B(n_368),
.C(n_370),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_380),
.B2(n_389),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_371),
.B(n_381),
.C(n_383),
.Y(n_494)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_380),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_471),
.Y(n_391)
);

A2O1A1Ixp33_ASAP7_75t_SL g503 ( 
.A1(n_392),
.A2(n_471),
.B(n_504),
.C(n_507),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_444),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_393),
.B(n_444),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_419),
.C(n_428),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g484 ( 
.A(n_394),
.B(n_419),
.CI(n_428),
.CON(n_484),
.SN(n_484)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_411),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_395),
.B(n_412),
.C(n_417),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_404),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_396),
.B(n_404),
.Y(n_477)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_397),
.Y(n_433)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_417),
.Y(n_411)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_415),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_426),
.B2(n_427),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_421),
.B(n_426),
.Y(n_463)
);

INVx3_ASAP7_75t_SL g423 ( 
.A(n_424),
.Y(n_423)
);

INVx8_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_426),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_426),
.A2(n_427),
.B1(n_465),
.B2(n_466),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_426),
.A2(n_463),
.B(n_466),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_436),
.C(n_442),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_429),
.B(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_430),
.B(n_432),
.Y(n_493)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_436),
.A2(n_437),
.B1(n_442),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx8_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_442),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_445),
.B(n_448),
.C(n_461),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_461),
.B2(n_462),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_457),
.B(n_460),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_458),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_452),
.Y(n_520)
);

INVx6_ASAP7_75t_SL g453 ( 
.A(n_454),
.Y(n_453)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

FAx1_ASAP7_75t_SL g511 ( 
.A(n_460),
.B(n_512),
.CI(n_513),
.CON(n_511),
.SN(n_511)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_460),
.B(n_512),
.C(n_513),
.Y(n_533)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_468),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_484),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_484),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_477),
.C(n_478),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_473),
.A2(n_474),
.B1(n_477),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_496),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.C(n_482),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_479),
.A2(n_480),
.B1(n_482),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g551 ( 
.A(n_484),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_486),
.B(n_498),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_487),
.A2(n_505),
.B(n_506),
.Y(n_504)
);

NOR2x1_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_495),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_495),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_492),
.C(n_494),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_501),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_492),
.A2(n_493),
.B1(n_494),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_494),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_500),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_523),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_511),
.B(n_522),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_511),
.B(n_522),
.Y(n_535)
);

BUFx24_ASAP7_75t_SL g550 ( 
.A(n_511),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_514),
.A2(n_515),
.B1(n_517),
.B2(n_521),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_514),
.A2(n_515),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_514),
.B(n_525),
.C(n_529),
.Y(n_541)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_517),
.Y(n_521)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_523),
.A2(n_535),
.B(n_536),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_524),
.B(n_533),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_533),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_525),
.A2(n_526),
.B1(n_527),
.B2(n_528),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_541),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_541),
.Y(n_542)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

BUFx12f_ASAP7_75t_L g547 ( 
.A(n_544),
.Y(n_547)
);

INVx13_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_548),
.Y(n_546)
);


endmodule