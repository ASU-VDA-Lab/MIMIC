module real_aes_18259_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_150;
wire n_147;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g816 ( .A(n_0), .B(n_817), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_1), .A2(n_4), .B1(n_194), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_2), .A2(n_43), .B1(n_132), .B2(n_134), .Y(n_131) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_3), .A2(n_23), .B1(n_134), .B2(n_158), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_5), .A2(n_16), .B1(n_175), .B2(n_212), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_6), .A2(n_61), .B1(n_160), .B2(n_232), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_7), .A2(n_17), .B1(n_132), .B2(n_179), .Y(n_505) );
INVx1_ASAP7_75t_L g817 ( .A(n_8), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_9), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_10), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_11), .A2(n_18), .B1(n_177), .B2(n_231), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_12), .A2(n_65), .B1(n_480), .B2(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_12), .Y(n_480) );
OR2x2_ASAP7_75t_L g112 ( .A(n_13), .B(n_38), .Y(n_112) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_14), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_15), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_19), .A2(n_98), .B1(n_175), .B2(n_194), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_20), .A2(n_39), .B1(n_208), .B2(n_209), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_21), .B(n_176), .Y(n_249) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_22), .A2(n_59), .B(n_149), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_24), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_25), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_26), .B(n_138), .Y(n_529) );
INVx4_ASAP7_75t_R g518 ( .A(n_27), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_28), .A2(n_47), .B1(n_140), .B2(n_142), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_29), .A2(n_54), .B1(n_142), .B2(n_175), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_30), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_31), .B(n_208), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_32), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_33), .B(n_134), .Y(n_536) );
INVx1_ASAP7_75t_L g584 ( .A(n_34), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_SL g565 ( .A1(n_35), .A2(n_132), .B(n_144), .C(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_36), .A2(n_55), .B1(n_132), .B2(n_142), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_37), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_40), .A2(n_86), .B1(n_132), .B2(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g116 ( .A1(n_41), .A2(n_53), .B1(n_117), .B2(n_118), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_41), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_42), .A2(n_46), .B1(n_132), .B2(n_179), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_44), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_45), .A2(n_60), .B1(n_175), .B2(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g533 ( .A(n_48), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_49), .B(n_132), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_50), .Y(n_546) );
INVx2_ASAP7_75t_L g470 ( .A(n_51), .Y(n_470) );
INVx1_ASAP7_75t_L g110 ( .A(n_52), .Y(n_110) );
BUFx3_ASAP7_75t_L g477 ( .A(n_52), .Y(n_477) );
INVx1_ASAP7_75t_L g117 ( .A(n_53), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_53), .B(n_831), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_56), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_57), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_58), .A2(n_87), .B1(n_132), .B2(n_142), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_62), .A2(n_75), .B1(n_140), .B2(n_197), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_63), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_64), .A2(n_77), .B1(n_132), .B2(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g481 ( .A(n_65), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_66), .A2(n_97), .B1(n_175), .B2(n_177), .Y(n_174) );
AND2x4_ASAP7_75t_L g128 ( .A(n_67), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g149 ( .A(n_68), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_69), .A2(n_89), .B1(n_140), .B2(n_142), .Y(n_580) );
AO22x1_ASAP7_75t_L g494 ( .A1(n_70), .A2(n_76), .B1(n_209), .B2(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g129 ( .A(n_71), .Y(n_129) );
AND2x2_ASAP7_75t_L g568 ( .A(n_72), .B(n_146), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_73), .B(n_160), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_74), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_78), .B(n_134), .Y(n_547) );
INVx2_ASAP7_75t_L g138 ( .A(n_79), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_80), .B(n_146), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_81), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_82), .A2(n_96), .B1(n_142), .B2(n_160), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_83), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_84), .B(n_167), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_85), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_88), .B(n_146), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_90), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_91), .B(n_146), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_92), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g802 ( .A(n_92), .Y(n_802) );
NAND2xp33_ASAP7_75t_L g252 ( .A(n_93), .B(n_176), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_94), .A2(n_160), .B(n_162), .C(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g520 ( .A(n_95), .B(n_521), .Y(n_520) );
NAND2xp33_ASAP7_75t_L g551 ( .A(n_99), .B(n_141), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_813), .B(n_819), .Y(n_100) );
OAI21xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_466), .B(n_471), .Y(n_101) );
OAI21xp33_ASAP7_75t_L g819 ( .A1(n_102), .A2(n_820), .B(n_830), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_113), .B(n_463), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx4_ASAP7_75t_L g465 ( .A(n_105), .Y(n_465) );
INVx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx8_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx5_ASAP7_75t_L g818 ( .A(n_107), .Y(n_818) );
INVx3_ASAP7_75t_L g829 ( .A(n_107), .Y(n_829) );
AND2x6_ASAP7_75t_SL g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_111), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2x1_ASAP7_75t_L g812 ( .A(n_112), .B(n_477), .Y(n_812) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
XNOR2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_119), .Y(n_115) );
OAI22x1_ASAP7_75t_L g484 ( .A1(n_119), .A2(n_485), .B1(n_799), .B2(n_803), .Y(n_484) );
NOR2x1p5_ASAP7_75t_L g119 ( .A(n_120), .B(n_373), .Y(n_119) );
NAND4xp75_ASAP7_75t_L g120 ( .A(n_121), .B(n_318), .C(n_338), .D(n_354), .Y(n_120) );
NOR2x1p5_ASAP7_75t_SL g121 ( .A(n_122), .B(n_288), .Y(n_121) );
NAND4xp75_ASAP7_75t_L g122 ( .A(n_123), .B(n_224), .C(n_265), .D(n_274), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_185), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_152), .Y(n_124) );
AND2x4_ASAP7_75t_L g398 ( .A(n_125), .B(n_325), .Y(n_398) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_126), .Y(n_241) );
INVx2_ASAP7_75t_L g259 ( .A(n_126), .Y(n_259) );
AND2x2_ASAP7_75t_L g282 ( .A(n_126), .B(n_244), .Y(n_282) );
OR2x2_ASAP7_75t_L g337 ( .A(n_126), .B(n_153), .Y(n_337) );
AO31x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .A3(n_145), .B(n_150), .Y(n_126) );
INVx2_ASAP7_75t_L g182 ( .A(n_127), .Y(n_182) );
AO31x2_ASAP7_75t_L g205 ( .A1(n_127), .A2(n_154), .A3(n_206), .B(n_214), .Y(n_205) );
AO31x2_ASAP7_75t_L g228 ( .A1(n_127), .A2(n_171), .A3(n_229), .B(n_235), .Y(n_228) );
AO31x2_ASAP7_75t_L g503 ( .A1(n_127), .A2(n_202), .A3(n_504), .B(n_507), .Y(n_503) );
BUFx10_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g164 ( .A(n_128), .Y(n_164) );
INVx1_ASAP7_75t_L g501 ( .A(n_128), .Y(n_501) );
BUFx10_ASAP7_75t_L g538 ( .A(n_128), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_135), .B1(n_139), .B2(n_143), .Y(n_130) );
INVx1_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
INVx4_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
INVx1_ASAP7_75t_L g197 ( .A(n_132), .Y(n_197) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_133), .Y(n_134) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_133), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_133), .Y(n_142) );
INVx2_ASAP7_75t_L g158 ( .A(n_133), .Y(n_158) );
INVx1_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
INVx1_ASAP7_75t_L g195 ( .A(n_133), .Y(n_195) );
INVx1_ASAP7_75t_L g210 ( .A(n_133), .Y(n_210) );
INVx1_ASAP7_75t_L g213 ( .A(n_133), .Y(n_213) );
INVx1_ASAP7_75t_L g233 ( .A(n_133), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_134), .B(n_561), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_135), .A2(n_143), .B1(n_193), .B2(n_196), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_135), .A2(n_143), .B1(n_207), .B2(n_211), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_135), .A2(n_143), .B1(n_220), .B2(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g497 ( .A(n_136), .Y(n_497) );
BUFx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g549 ( .A(n_137), .Y(n_549) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx8_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx1_ASAP7_75t_L g162 ( .A(n_138), .Y(n_162) );
INVx1_ASAP7_75t_L g532 ( .A(n_138), .Y(n_532) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g208 ( .A(n_141), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g517 ( .A1(n_141), .A2(n_213), .B1(n_518), .B2(n_519), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_142), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g582 ( .A(n_142), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g155 ( .A1(n_143), .A2(n_156), .B1(n_159), .B2(n_161), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_143), .A2(n_174), .B1(n_178), .B2(n_180), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_143), .A2(n_180), .B1(n_230), .B2(n_234), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_143), .A2(n_251), .B(n_252), .Y(n_250) );
OAI22x1_ASAP7_75t_L g504 ( .A1(n_143), .A2(n_161), .B1(n_505), .B2(n_506), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_143), .A2(n_497), .B1(n_572), .B2(n_573), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_143), .A2(n_161), .B1(n_580), .B2(n_581), .Y(n_579) );
INVx6_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
O2A1O1Ixp5_ASAP7_75t_L g247 ( .A1(n_144), .A2(n_179), .B(n_248), .C(n_249), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_144), .A2(n_494), .B(n_496), .C(n_500), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_144), .A2(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_144), .B(n_494), .Y(n_596) );
AO31x2_ASAP7_75t_L g570 ( .A1(n_145), .A2(n_538), .A3(n_571), .B(n_574), .Y(n_570) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_146), .B(n_554), .Y(n_553) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_147), .B(n_151), .Y(n_150) );
BUFx3_ASAP7_75t_L g154 ( .A(n_147), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_147), .B(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_147), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_SL g245 ( .A(n_147), .Y(n_245) );
AND2x2_ASAP7_75t_L g537 ( .A(n_147), .B(n_538), .Y(n_537) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
AND2x2_ASAP7_75t_L g255 ( .A(n_152), .B(n_256), .Y(n_255) );
AND2x4_ASAP7_75t_L g405 ( .A(n_152), .B(n_282), .Y(n_405) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_169), .Y(n_152) );
OR2x2_ASAP7_75t_L g242 ( .A(n_153), .B(n_243), .Y(n_242) );
BUFx2_ASAP7_75t_L g273 ( .A(n_153), .Y(n_273) );
AND2x2_ASAP7_75t_L g279 ( .A(n_153), .B(n_170), .Y(n_279) );
INVx1_ASAP7_75t_L g297 ( .A(n_153), .Y(n_297) );
INVx2_ASAP7_75t_L g326 ( .A(n_153), .Y(n_326) );
AO31x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .A3(n_163), .B(n_165), .Y(n_153) );
INVx2_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_158), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_161), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_SL g180 ( .A(n_162), .Y(n_180) );
AO31x2_ASAP7_75t_L g218 ( .A1(n_163), .A2(n_198), .A3(n_219), .B(n_222), .Y(n_218) );
AO31x2_ASAP7_75t_L g578 ( .A1(n_163), .A2(n_171), .A3(n_579), .B(n_583), .Y(n_578) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_SL g253 ( .A(n_164), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_168), .Y(n_165) );
INVx2_ASAP7_75t_L g199 ( .A(n_166), .Y(n_199) );
NOR2xp33_ASAP7_75t_SL g235 ( .A(n_166), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g172 ( .A(n_167), .Y(n_172) );
INVx2_ASAP7_75t_L g202 ( .A(n_167), .Y(n_202) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_167), .A2(n_499), .B(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g302 ( .A(n_169), .Y(n_302) );
INVx2_ASAP7_75t_L g307 ( .A(n_169), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_169), .B(n_258), .Y(n_312) );
AND2x2_ASAP7_75t_L g335 ( .A(n_169), .B(n_314), .Y(n_335) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_169), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_169), .B(n_390), .Y(n_389) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx2_ASAP7_75t_L g324 ( .A(n_170), .Y(n_324) );
AND2x2_ASAP7_75t_L g372 ( .A(n_170), .B(n_326), .Y(n_372) );
AO31x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .A3(n_181), .B(n_183), .Y(n_170) );
AOI21x1_ASAP7_75t_L g557 ( .A1(n_171), .A2(n_558), .B(n_568), .Y(n_557) );
BUFx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_172), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g521 ( .A(n_172), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_172), .B(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_172), .B(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_176), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_179), .A2(n_546), .B(n_547), .C(n_548), .Y(n_545) );
AO31x2_ASAP7_75t_L g191 ( .A1(n_181), .A2(n_192), .A3(n_198), .B(n_200), .Y(n_191) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_182), .A2(n_513), .B(n_516), .Y(n_512) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_203), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_187), .B(n_316), .Y(n_363) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2x1p5_ASAP7_75t_L g360 ( .A(n_188), .B(n_316), .Y(n_360) );
INVx1_ASAP7_75t_L g461 ( .A(n_188), .Y(n_461) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g411 ( .A(n_189), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g264 ( .A(n_190), .Y(n_264) );
OR2x2_ASAP7_75t_L g345 ( .A(n_190), .B(n_217), .Y(n_345) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g287 ( .A(n_191), .Y(n_287) );
AND2x4_ASAP7_75t_L g293 ( .A(n_191), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_195), .B(n_563), .Y(n_562) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_198), .A2(n_512), .B(n_520), .Y(n_511) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_202), .B(n_223), .Y(n_222) );
AOI32xp33_ASAP7_75t_L g431 ( .A1(n_203), .A2(n_334), .A3(n_432), .B1(n_434), .B2(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g380 ( .A(n_204), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_216), .Y(n_204) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_205), .Y(n_226) );
OR2x2_ASAP7_75t_L g262 ( .A(n_205), .B(n_218), .Y(n_262) );
INVx1_ASAP7_75t_L g277 ( .A(n_205), .Y(n_277) );
AND2x2_ASAP7_75t_L g286 ( .A(n_205), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g292 ( .A(n_205), .Y(n_292) );
INVx2_ASAP7_75t_L g317 ( .A(n_205), .Y(n_317) );
AND2x2_ASAP7_75t_L g436 ( .A(n_205), .B(n_228), .Y(n_436) );
OAI21xp33_ASAP7_75t_SL g528 ( .A1(n_209), .A2(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_216), .B(n_269), .Y(n_356) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g227 ( .A(n_218), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g285 ( .A(n_218), .Y(n_285) );
INVx2_ASAP7_75t_L g294 ( .A(n_218), .Y(n_294) );
AND2x4_ASAP7_75t_L g316 ( .A(n_218), .B(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_218), .Y(n_408) );
AOI22x1_ASAP7_75t_SL g224 ( .A1(n_225), .A2(n_237), .B1(n_255), .B2(n_260), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NAND4xp25_ASAP7_75t_L g385 ( .A(n_227), .B(n_386), .C(n_387), .D(n_388), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_227), .B(n_286), .Y(n_416) );
INVx4_ASAP7_75t_SL g269 ( .A(n_228), .Y(n_269) );
BUFx2_ASAP7_75t_L g332 ( .A(n_228), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_228), .B(n_277), .Y(n_395) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_233), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g357 ( .A(n_239), .B(n_306), .Y(n_357) );
NOR2x1_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x4_ASAP7_75t_L g280 ( .A(n_243), .B(n_258), .Y(n_280) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_244), .B(n_259), .Y(n_304) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_254), .Y(n_244) );
OAI21x1_ASAP7_75t_L g299 ( .A1(n_245), .A2(n_246), .B(n_254), .Y(n_299) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_250), .B(n_253), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_256), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g322 ( .A(n_256), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g361 ( .A(n_257), .B(n_279), .Y(n_361) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g404 ( .A(n_259), .B(n_314), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_260), .A2(n_377), .B1(n_379), .B2(n_382), .C(n_384), .Y(n_376) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g270 ( .A(n_262), .Y(n_270) );
OR2x2_ASAP7_75t_L g370 ( .A(n_262), .B(n_309), .Y(n_370) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_271), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_266), .A2(n_392), .B1(n_396), .B2(n_399), .Y(n_391) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_270), .Y(n_266) );
AND2x4_ASAP7_75t_L g315 ( .A(n_267), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g427 ( .A(n_267), .B(n_345), .Y(n_427) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g275 ( .A(n_269), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g291 ( .A(n_269), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g350 ( .A(n_269), .B(n_287), .Y(n_350) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_269), .Y(n_367) );
INVx1_ASAP7_75t_L g381 ( .A(n_269), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_269), .B(n_294), .Y(n_424) );
AND2x4_ASAP7_75t_L g331 ( .A(n_270), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g329 ( .A(n_272), .Y(n_329) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_273), .B(n_314), .Y(n_313) );
NAND2x1_ASAP7_75t_L g433 ( .A(n_273), .B(n_335), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_278), .B1(n_281), .B2(n_283), .Y(n_274) );
AND2x2_ASAP7_75t_L g300 ( .A(n_275), .B(n_293), .Y(n_300) );
INVx1_ASAP7_75t_L g341 ( .A(n_275), .Y(n_341) );
AND2x2_ASAP7_75t_L g448 ( .A(n_275), .B(n_309), .Y(n_448) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_SL g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g281 ( .A(n_279), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g421 ( .A(n_279), .Y(n_421) );
AND2x2_ASAP7_75t_L g438 ( .A(n_279), .B(n_298), .Y(n_438) );
AND2x2_ASAP7_75t_L g454 ( .A(n_279), .B(n_404), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_280), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g377 ( .A(n_280), .B(n_378), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_280), .A2(n_370), .B1(n_385), .B2(n_389), .Y(n_384) );
INVx1_ASAP7_75t_L g340 ( .A(n_282), .Y(n_340) );
AND2x2_ASAP7_75t_L g371 ( .A(n_282), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_282), .B(n_378), .Y(n_400) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g406 ( .A(n_286), .B(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_286), .A2(n_310), .B1(n_415), .B2(n_417), .Y(n_414) );
INVx3_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
AND2x2_ASAP7_75t_L g441 ( .A(n_287), .B(n_294), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_305), .Y(n_288) );
AOI32xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_295), .A3(n_298), .B1(n_300), .B2(n_301), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_292), .Y(n_387) );
INVx1_ASAP7_75t_L g412 ( .A(n_292), .Y(n_412) );
INVx3_ASAP7_75t_L g368 ( .A(n_293), .Y(n_368) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OAI221xp5_ASAP7_75t_L g443 ( .A1(n_296), .A2(n_444), .B1(n_445), .B2(n_446), .C(n_447), .Y(n_443) );
BUFx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g420 ( .A(n_298), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g456 ( .A(n_298), .B(n_417), .Y(n_456) );
BUFx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g314 ( .A(n_299), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_301), .B(n_329), .Y(n_328) );
AO22x1_ASAP7_75t_L g358 ( .A1(n_301), .A2(n_359), .B1(n_361), .B2(n_362), .Y(n_358) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_301), .B(n_329), .Y(n_462) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g378 ( .A(n_302), .Y(n_378) );
INVx1_ASAP7_75t_L g388 ( .A(n_302), .Y(n_388) );
AND2x2_ASAP7_75t_L g308 ( .A(n_303), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_304), .Y(n_390) );
INVx1_ASAP7_75t_L g430 ( .A(n_304), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_308), .B(n_310), .C(n_315), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2x1p5_ASAP7_75t_L g417 ( .A(n_307), .B(n_337), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_308), .B(n_367), .Y(n_444) );
AOI31xp33_ASAP7_75t_L g327 ( .A1(n_309), .A2(n_328), .A3(n_330), .B(n_333), .Y(n_327) );
INVx4_ASAP7_75t_L g386 ( .A(n_309), .Y(n_386) );
OR2x2_ASAP7_75t_L g423 ( .A(n_309), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x4_ASAP7_75t_L g325 ( .A(n_314), .B(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_316), .Y(n_321) );
AND2x2_ASAP7_75t_L g352 ( .A(n_316), .B(n_350), .Y(n_352) );
NOR2xp67_ASAP7_75t_L g318 ( .A(n_319), .B(n_327), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g445 ( .A(n_322), .Y(n_445) );
INVx1_ASAP7_75t_L g353 ( .A(n_323), .Y(n_353) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g383 ( .A(n_324), .Y(n_383) );
AND2x2_ASAP7_75t_L g382 ( .A(n_325), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI322xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .A3(n_342), .B1(n_346), .B2(n_349), .C1(n_351), .C2(n_353), .Y(n_339) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI211x1_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B(n_358), .C(n_364), .Y(n_354) );
INVx1_ASAP7_75t_L g459 ( .A(n_355), .Y(n_459) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g413 ( .A(n_357), .Y(n_413) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OA21x2_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_369), .B(n_371), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx2_ASAP7_75t_L g434 ( .A(n_368), .Y(n_434) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp33_ASAP7_75t_L g429 ( .A(n_372), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_442), .Y(n_373) );
NOR3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_409), .C(n_425), .Y(n_374) );
NAND3xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_391), .C(n_401), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_378), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI21xp33_ASAP7_75t_L g437 ( .A1(n_382), .A2(n_438), .B(n_439), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_386), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_386), .B(n_436), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_387), .B(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_388), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_398), .A2(n_448), .B(n_449), .Y(n_447) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B(n_406), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_413), .B(n_414), .C(n_418), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_SL g428 ( .A(n_420), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_424), .Y(n_446) );
OAI211xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B(n_431), .C(n_437), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_436), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g457 ( .A(n_436), .Y(n_457) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g453 ( .A(n_441), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_451), .C(n_458), .Y(n_442) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI21xp33_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_455), .B(n_457), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI21xp33_ASAP7_75t_R g458 ( .A1(n_459), .A2(n_460), .B(n_462), .Y(n_458) );
NOR2x1_ASAP7_75t_R g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVxp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_469), .B(n_827), .Y(n_826) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g474 ( .A(n_470), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_470), .B(n_810), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_470), .B(n_829), .Y(n_833) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_478), .B(n_805), .Y(n_471) );
BUFx12f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x6_ASAP7_75t_SL g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI22xp33_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_482), .B1(n_483), .B2(n_804), .Y(n_478) );
INVx1_ASAP7_75t_L g804 ( .A(n_479), .Y(n_804) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_709), .Y(n_485) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_638), .C(n_680), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_612), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_522), .B1(n_587), .B2(n_598), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_509), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_491), .A2(n_632), .B(n_634), .Y(n_631) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_491), .A2(n_705), .B(n_706), .Y(n_704) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_502), .Y(n_491) );
INVx2_ASAP7_75t_L g624 ( .A(n_492), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_492), .B(n_503), .Y(n_654) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g595 ( .A(n_496), .Y(n_595) );
OAI21x1_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_499), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_497), .A2(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g597 ( .A(n_500), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_501), .A2(n_559), .B(n_565), .Y(n_558) );
AND2x2_ASAP7_75t_L g694 ( .A(n_502), .B(n_541), .Y(n_694) );
INVx1_ASAP7_75t_L g727 ( .A(n_502), .Y(n_727) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g589 ( .A(n_503), .B(n_542), .Y(n_589) );
AND2x2_ASAP7_75t_L g620 ( .A(n_503), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g629 ( .A(n_503), .Y(n_629) );
OR2x2_ASAP7_75t_L g648 ( .A(n_503), .B(n_511), .Y(n_648) );
AND2x2_ASAP7_75t_L g663 ( .A(n_503), .B(n_511), .Y(n_663) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_510), .B(n_662), .Y(n_705) );
OR2x2_ASAP7_75t_L g793 ( .A(n_510), .B(n_654), .Y(n_793) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g621 ( .A(n_511), .Y(n_621) );
AND2x2_ASAP7_75t_L g630 ( .A(n_511), .B(n_593), .Y(n_630) );
AND2x2_ASAP7_75t_L g633 ( .A(n_511), .B(n_542), .Y(n_633) );
AND2x2_ASAP7_75t_L g652 ( .A(n_511), .B(n_541), .Y(n_652) );
AND2x4_ASAP7_75t_L g671 ( .A(n_511), .B(n_594), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_539), .B(n_576), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_523), .B(n_666), .Y(n_769) );
CKINVDCx14_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_525), .B(n_586), .Y(n_585) );
INVx3_ASAP7_75t_L g602 ( .A(n_525), .Y(n_602) );
OR2x2_ASAP7_75t_L g610 ( .A(n_525), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_525), .B(n_603), .Y(n_635) );
AND2x2_ASAP7_75t_L g660 ( .A(n_525), .B(n_578), .Y(n_660) );
AND2x2_ASAP7_75t_L g678 ( .A(n_525), .B(n_608), .Y(n_678) );
INVx1_ASAP7_75t_L g717 ( .A(n_525), .Y(n_717) );
AND2x2_ASAP7_75t_L g719 ( .A(n_525), .B(n_720), .Y(n_719) );
NAND2x1p5_ASAP7_75t_SL g738 ( .A(n_525), .B(n_659), .Y(n_738) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_534), .B(n_537), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
BUFx4f_ASAP7_75t_L g564 ( .A(n_532), .Y(n_564) );
INVx1_ASAP7_75t_L g554 ( .A(n_538), .Y(n_554) );
OAI32xp33_ASAP7_75t_L g622 ( .A1(n_539), .A2(n_614), .A3(n_623), .B1(n_625), .B2(n_627), .Y(n_622) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_555), .Y(n_539) );
INVx1_ASAP7_75t_L g662 ( .A(n_540), .Y(n_662) );
AND2x2_ASAP7_75t_L g670 ( .A(n_540), .B(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g669 ( .A(n_541), .B(n_593), .Y(n_669) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g619 ( .A(n_542), .Y(n_619) );
AND2x2_ASAP7_75t_L g628 ( .A(n_542), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g734 ( .A(n_542), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
OAI21x1_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_550), .B(n_553), .Y(n_544) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g604 ( .A(n_555), .Y(n_604) );
OR2x2_ASAP7_75t_L g614 ( .A(n_555), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g736 ( .A(n_555), .Y(n_736) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_569), .Y(n_555) );
AND2x2_ASAP7_75t_L g637 ( .A(n_556), .B(n_570), .Y(n_637) );
INVx2_ASAP7_75t_L g659 ( .A(n_556), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_556), .B(n_578), .Y(n_679) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g586 ( .A(n_557), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_562), .B(n_564), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_569), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g668 ( .A(n_569), .Y(n_668) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
BUFx2_ASAP7_75t_L g608 ( .A(n_570), .Y(n_608) );
OR2x2_ASAP7_75t_L g674 ( .A(n_570), .B(n_578), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_570), .B(n_578), .Y(n_707) );
INVx2_ASAP7_75t_L g655 ( .A(n_576), .Y(n_655) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_585), .Y(n_576) );
OR2x2_ASAP7_75t_L g642 ( .A(n_577), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g720 ( .A(n_577), .Y(n_720) );
INVx1_ASAP7_75t_L g603 ( .A(n_578), .Y(n_603) );
INVx1_ASAP7_75t_L g611 ( .A(n_578), .Y(n_611) );
INVx1_ASAP7_75t_L g626 ( .A(n_578), .Y(n_626) );
OR2x2_ASAP7_75t_L g730 ( .A(n_585), .B(n_707), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_586), .B(n_602), .Y(n_643) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_586), .Y(n_645) );
OR2x2_ASAP7_75t_L g744 ( .A(n_586), .B(n_668), .Y(n_744) );
INVxp67_ASAP7_75t_L g768 ( .A(n_586), .Y(n_768) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
NAND2x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_589), .B(n_630), .Y(n_697) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g646 ( .A(n_591), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g759 ( .A(n_592), .Y(n_759) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g788 ( .A(n_593), .B(n_621), .Y(n_788) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g714 ( .A(n_594), .B(n_621), .Y(n_714) );
AOI21x1_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_597), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_605), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_601), .B(n_637), .Y(n_751) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx2_ASAP7_75t_L g615 ( .A(n_602), .Y(n_615) );
AND2x2_ASAP7_75t_L g665 ( .A(n_602), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_602), .B(n_659), .Y(n_708) );
OR2x2_ASAP7_75t_L g780 ( .A(n_602), .B(n_667), .Y(n_780) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g700 ( .A(n_606), .B(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx2_ASAP7_75t_L g691 ( .A(n_607), .Y(n_691) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g681 ( .A(n_610), .B(n_682), .Y(n_681) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_610), .Y(n_692) );
OR2x2_ASAP7_75t_L g743 ( .A(n_610), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g798 ( .A(n_610), .Y(n_798) );
AOI211xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_616), .B(n_622), .C(n_631), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g687 ( .A(n_615), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_615), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g760 ( .A(n_615), .B(n_637), .Y(n_760) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_618), .B(n_663), .Y(n_685) );
NAND2x1p5_ASAP7_75t_L g702 ( .A(n_618), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g770 ( .A(n_618), .B(n_771), .Y(n_770) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g713 ( .A(n_619), .Y(n_713) );
AND2x2_ASAP7_75t_L g741 ( .A(n_620), .B(n_669), .Y(n_741) );
INVx2_ASAP7_75t_L g764 ( .A(n_620), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_620), .B(n_662), .Y(n_796) );
AND2x4_ASAP7_75t_SL g750 ( .A(n_623), .B(n_628), .Y(n_750) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g703 ( .A(n_624), .B(n_629), .Y(n_703) );
OR2x2_ASAP7_75t_L g755 ( .A(n_624), .B(n_648), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_625), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_625), .B(n_637), .Y(n_791) );
BUFx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g739 ( .A(n_626), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g722 ( .A(n_628), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_628), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g772 ( .A(n_629), .Y(n_772) );
BUFx2_ASAP7_75t_L g640 ( .A(n_630), .Y(n_640) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g758 ( .A(n_633), .B(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g682 ( .A(n_637), .Y(n_682) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_637), .Y(n_699) );
NAND3xp33_ASAP7_75t_SL g638 ( .A(n_639), .B(n_649), .C(n_664), .Y(n_638) );
AOI22xp33_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_641), .B1(n_644), .B2(n_646), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI222xp33_ASAP7_75t_L g752 ( .A1(n_646), .A2(n_672), .B1(n_753), .B2(n_756), .C1(n_758), .C2(n_760), .Y(n_752) );
AND2x2_ASAP7_75t_L g784 ( .A(n_647), .B(n_733), .Y(n_784) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g732 ( .A(n_648), .B(n_733), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_655), .B1(n_656), .B2(n_661), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx2_ASAP7_75t_SL g728 ( .A(n_652), .Y(n_728) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_660), .Y(n_656) );
AND2x2_ASAP7_75t_L g715 ( .A(n_657), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g673 ( .A(n_658), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g667 ( .A(n_659), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g782 ( .A(n_660), .Y(n_782) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_663), .B(n_759), .Y(n_778) );
INVx1_ASAP7_75t_L g795 ( .A(n_663), .Y(n_795) );
AOI222xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_669), .B1(n_670), .B2(n_672), .C1(n_675), .C2(n_676), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_671), .Y(n_675) );
AND2x2_ASAP7_75t_L g693 ( .A(n_671), .B(n_694), .Y(n_693) );
INVx3_ASAP7_75t_L g724 ( .A(n_671), .Y(n_724) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g688 ( .A(n_674), .Y(n_688) );
OR2x2_ASAP7_75t_L g757 ( .A(n_674), .B(n_738), .Y(n_757) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OAI211xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B(n_686), .C(n_695), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_693), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_687), .A2(n_725), .B1(n_774), .B2(n_777), .C(n_779), .Y(n_773) );
AND2x4_ASAP7_75t_L g716 ( .A(n_688), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g747 ( .A(n_694), .Y(n_747) );
AOI211x1_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B(n_700), .C(n_704), .Y(n_695) );
INVxp67_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g765 ( .A(n_703), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g753 ( .A(n_706), .B(n_754), .C(n_755), .Y(n_753) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g789 ( .A(n_707), .Y(n_789) );
NOR2x1_ASAP7_75t_L g709 ( .A(n_710), .B(n_761), .Y(n_709) );
NAND4xp25_ASAP7_75t_L g710 ( .A(n_711), .B(n_718), .C(n_740), .D(n_752), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_715), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
AND2x2_ASAP7_75t_L g771 ( .A(n_714), .B(n_772), .Y(n_771) );
AOI221x1_ASAP7_75t_L g740 ( .A1(n_716), .A2(n_741), .B1(n_742), .B2(n_745), .C(n_748), .Y(n_740) );
AND2x2_ASAP7_75t_L g766 ( .A(n_716), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g776 ( .A(n_717), .Y(n_776) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B1(n_725), .B2(n_729), .C(n_731), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_723), .B(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_728), .A2(n_732), .B1(n_735), .B2(n_737), .Y(n_731) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_732), .A2(n_749), .B(n_751), .Y(n_748) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g754 ( .A(n_734), .Y(n_754) );
OR2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVxp67_ASAP7_75t_L g775 ( .A(n_744), .Y(n_775) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_757), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_794) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_773), .C(n_785), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_766), .B1(n_769), .B2(n_770), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVxp67_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g781 ( .A(n_768), .B(n_782), .Y(n_781) );
NAND2x1_ASAP7_75t_L g797 ( .A(n_768), .B(n_798), .Y(n_797) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx2_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B(n_783), .Y(n_779) );
INVx1_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_789), .B1(n_790), .B2(n_792), .C(n_794), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx3_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
INVx4_ASAP7_75t_L g803 ( .A(n_799), .Y(n_803) );
BUFx12f_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
AND2x2_ASAP7_75t_L g811 ( .A(n_801), .B(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx6_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx10_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
CKINVDCx16_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_818), .Y(n_815) );
INVx2_ASAP7_75t_SL g828 ( .A(n_816), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_823), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
OR2x6_ASAP7_75t_L g824 ( .A(n_825), .B(n_829), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
OR2x4_ASAP7_75t_L g832 ( .A(n_827), .B(n_833), .Y(n_832) );
BUFx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
BUFx3_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
endmodule