module real_jpeg_27034_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_150;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g46 ( 
.A(n_0),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_50),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_5),
.A2(n_24),
.B1(n_26),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_8),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_8),
.A2(n_11),
.B(n_45),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_9),
.A2(n_24),
.B1(n_26),
.B2(n_33),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_9),
.A2(n_33),
.B1(n_70),
.B2(n_71),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_9),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_11),
.A2(n_24),
.B1(n_26),
.B2(n_36),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_11),
.A2(n_36),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_11),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_11),
.A2(n_28),
.B(n_75),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_11),
.B(n_73),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_11),
.A2(n_24),
.B(n_30),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_11),
.B(n_23),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_120),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_119),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_93),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_16),
.B(n_93),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_79),
.B2(n_92),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_52),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_38),
.B(n_51),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_20),
.A2(n_86),
.B1(n_97),
.B2(n_126),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_20),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_20),
.B(n_150),
.C(n_151),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_20),
.A2(n_126),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_32),
.B1(n_34),
.B2(n_37),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_22),
.B(n_23),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_24),
.A2(n_26),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_24),
.A2(n_36),
.B(n_42),
.C(n_180),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_28),
.A2(n_29),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_31),
.B(n_36),
.C(n_160),
.Y(n_159)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_32),
.A2(n_37),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_34),
.B(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_36),
.A2(n_70),
.B(n_74),
.C(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_36),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_36),
.B(n_43),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_39),
.A2(n_43),
.B1(n_64),
.B2(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_39),
.B(n_43),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_47),
.B(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_44),
.B(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_59),
.Y(n_58)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_65),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_66),
.B1(n_67),
.B2(n_78),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_54),
.A2(n_61),
.B1(n_78),
.B2(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_58),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_57),
.B(n_106),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_58),
.A2(n_83),
.B1(n_107),
.B2(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_73),
.B1(n_76),
.B2(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_76),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_70),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.C(n_89),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_81),
.A2(n_84),
.B1(n_174),
.B2(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_81),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_83),
.A2(n_104),
.B(n_132),
.Y(n_150)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_83),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_84),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_84),
.A2(n_174),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_84),
.B(n_131),
.C(n_184),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_84),
.B(n_165),
.C(n_173),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_86),
.B(n_126),
.C(n_127),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_89),
.A2(n_90),
.B1(n_136),
.B2(n_137),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_89),
.B(n_109),
.C(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_89),
.A2(n_90),
.B1(n_108),
.B2(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_116),
.C(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_100),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_98),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_100),
.B(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_112),
.C(n_115),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_101),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_108),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_108),
.B1(n_109),
.B2(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_108),
.A2(n_109),
.B1(n_179),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_109),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_116),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_225),
.B(n_230),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_153),
.B(n_213),
.C(n_224),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_143),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_123),
.B(n_143),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_133),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_124),
.B(n_134),
.C(n_141),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_131),
.A2(n_148),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_131),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_197),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_140),
.B2(n_141),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_149),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_144),
.B(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_147),
.B(n_149),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_150),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_212),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_207),
.B(n_211),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_175),
.B(n_206),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_164),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_164),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_159),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_163),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_171),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_168),
.B(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_172),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_201),
.B(n_205),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_186),
.B(n_200),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_181),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_179),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_182),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_183),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B(n_199),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_196),
.B(n_198),
.Y(n_190)
);

INVx5_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_209),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_215),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_222),
.B2(n_223),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_220),
.C(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_222),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_226),
.B(n_227),
.Y(n_230)
);


endmodule