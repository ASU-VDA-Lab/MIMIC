module fake_jpeg_9885_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_41),
.Y(n_68)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_44),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_14),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_16),
.B(n_1),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_57),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_48),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_59),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_80),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_35),
.B1(n_28),
.B2(n_20),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_63),
.A2(n_72),
.B1(n_77),
.B2(n_30),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_70),
.Y(n_99)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_36),
.A2(n_35),
.B1(n_16),
.B2(n_30),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_77),
.B1(n_30),
.B2(n_33),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_39),
.A2(n_35),
.B1(n_20),
.B2(n_28),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_62),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_39),
.A2(n_28),
.B1(n_26),
.B2(n_25),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_33),
.C(n_27),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_85),
.B(n_97),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_87),
.B(n_98),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_89),
.A2(n_102),
.B1(n_112),
.B2(n_115),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_50),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_113),
.C(n_100),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_57),
.B(n_40),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_21),
.B(n_19),
.C(n_46),
.Y(n_103)
);

XOR2x2_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_34),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_106),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_107),
.B1(n_122),
.B2(n_123),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_75),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_113),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_55),
.A2(n_27),
.B1(n_33),
.B2(n_21),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_12),
.B1(n_11),
.B2(n_13),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_45),
.B1(n_38),
.B2(n_27),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_26),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_64),
.A2(n_25),
.B1(n_26),
.B2(n_18),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_68),
.B(n_29),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_75),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_69),
.A2(n_25),
.B1(n_26),
.B2(n_18),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_24),
.B1(n_23),
.B2(n_31),
.Y(n_146)
);

AOI22x1_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_69),
.B1(n_54),
.B2(n_67),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_131),
.B(n_138),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_130),
.B(n_2),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g131 ( 
.A1(n_85),
.A2(n_56),
.B(n_18),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_86),
.A2(n_70),
.B1(n_78),
.B2(n_58),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_136),
.A2(n_140),
.B1(n_119),
.B2(n_107),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_150),
.C(n_151),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_1),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_86),
.A2(n_18),
.B1(n_31),
.B2(n_29),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_92),
.A2(n_90),
.B1(n_89),
.B2(n_104),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_146),
.B1(n_149),
.B2(n_98),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_24),
.B1(n_31),
.B2(n_34),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_116),
.B(n_121),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_109),
.A2(n_59),
.B1(n_84),
.B2(n_13),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_86),
.C(n_92),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_90),
.B(n_2),
.C(n_3),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_87),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_2),
.C(n_3),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_151),
.C(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_156),
.B(n_157),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_101),
.B1(n_108),
.B2(n_119),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_165),
.B1(n_177),
.B2(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_103),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_161),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_87),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_146),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_99),
.B1(n_112),
.B2(n_115),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_117),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_164),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_120),
.B1(n_114),
.B2(n_124),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_95),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_167),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_168),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_11),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_172),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_12),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_118),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_94),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_176),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_135),
.B(n_12),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_88),
.B1(n_91),
.B2(n_116),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_181),
.B(n_135),
.CI(n_4),
.CON(n_200),
.SN(n_200)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_153),
.B1(n_142),
.B2(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_183),
.A2(n_185),
.B(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_94),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_127),
.A2(n_88),
.B1(n_116),
.B2(n_94),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_134),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_189),
.A2(n_190),
.B(n_162),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_131),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_169),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_138),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_194),
.B(n_196),
.C(n_216),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_183),
.A2(n_131),
.B1(n_147),
.B2(n_155),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_200),
.B(n_157),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_161),
.C(n_160),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_202),
.A2(n_221),
.B1(n_5),
.B2(n_6),
.Y(n_241)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_204),
.Y(n_246)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_159),
.A2(n_128),
.B1(n_142),
.B2(n_154),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_211),
.B(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_163),
.A2(n_128),
.B1(n_153),
.B2(n_116),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_168),
.B1(n_4),
.B2(n_5),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_184),
.A2(n_3),
.B(n_4),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_217),
.A2(n_166),
.B(n_185),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_168),
.B(n_6),
.Y(n_239)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_226),
.B1(n_227),
.B2(n_229),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_SL g262 ( 
.A(n_224),
.B(n_225),
.C(n_242),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_175),
.B1(n_156),
.B2(n_177),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_181),
.B1(n_170),
.B2(n_173),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_171),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_231),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_170),
.B1(n_176),
.B2(n_172),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_241),
.B1(n_247),
.B2(n_249),
.Y(n_251)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_233),
.B(n_238),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_96),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_197),
.C(n_196),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_237),
.B(n_239),
.C(n_244),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_3),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_245),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_201),
.A2(n_5),
.B(n_7),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_198),
.B(n_5),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_243),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_192),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_249)
);

XOR2x1_ASAP7_75t_SL g255 ( 
.A(n_239),
.B(n_200),
.Y(n_255)
);

FAx1_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_217),
.CI(n_224),
.CON(n_273),
.SN(n_273)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_211),
.B1(n_221),
.B2(n_206),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_256),
.A2(n_258),
.B1(n_237),
.B2(n_210),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_216),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_260),
.C(n_263),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_215),
.B1(n_205),
.B2(n_213),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_243),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_197),
.C(n_209),
.Y(n_263)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_264),
.B(n_210),
.Y(n_286)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_219),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_267),
.C(n_270),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_219),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_195),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_271),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_193),
.C(n_191),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_225),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_237),
.Y(n_272)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_277),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_235),
.B(n_246),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_278),
.B1(n_282),
.B2(n_253),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_269),
.A2(n_231),
.B(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_276),
.Y(n_301)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_266),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_240),
.B1(n_238),
.B2(n_244),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_285),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_250),
.A2(n_223),
.B1(n_249),
.B2(n_205),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_236),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_242),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_191),
.C(n_222),
.Y(n_285)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_253),
.B1(n_265),
.B2(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_289),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_251),
.B(n_267),
.C(n_253),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_282),
.B1(n_273),
.B2(n_277),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_293),
.A2(n_295),
.B1(n_200),
.B2(n_8),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_253),
.B1(n_252),
.B2(n_263),
.Y(n_295)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVx11_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_284),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_283),
.C(n_280),
.Y(n_314)
);

INVx13_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_273),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_199),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_279),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_305),
.A2(n_309),
.B(n_7),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_308),
.B1(n_311),
.B2(n_312),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_290),
.B1(n_301),
.B2(n_293),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_199),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_315),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_304),
.A2(n_300),
.B1(n_294),
.B2(n_298),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_283),
.B1(n_285),
.B2(n_279),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_313),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_280),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_291),
.B1(n_303),
.B2(n_295),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_315),
.A2(n_292),
.B(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_320),
.C(n_321),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_299),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_296),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_324),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_316),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_311),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_313),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_330),
.B(n_314),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_306),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_319),
.B(n_318),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_327),
.C(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

AOI21x1_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_335),
.B(n_320),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_321),
.B(n_8),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_9),
.C(n_324),
.Y(n_341)
);


endmodule