module fake_jpeg_7707_n_334 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_24),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_17),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_22),
.B1(n_30),
.B2(n_21),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_46),
.A2(n_62),
.B1(n_65),
.B2(n_23),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_47),
.B(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_58),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_22),
.B1(n_30),
.B2(n_21),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_64),
.B1(n_70),
.B2(n_25),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_22),
.B1(n_21),
.B2(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_22),
.B1(n_25),
.B2(n_17),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_25),
.B1(n_17),
.B2(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_25),
.B1(n_29),
.B2(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_72),
.B(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_29),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_82),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_28),
.B(n_27),
.C(n_34),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_79),
.B(n_93),
.Y(n_117)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_19),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_90),
.Y(n_125)
);

AO22x2_ASAP7_75t_SL g84 ( 
.A1(n_60),
.A2(n_18),
.B1(n_19),
.B2(n_44),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_52),
.B(n_54),
.C(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_56),
.B1(n_26),
.B2(n_20),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_23),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_51),
.A2(n_34),
.B1(n_27),
.B2(n_28),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_27),
.B1(n_51),
.B2(n_63),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_98),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_46),
.B1(n_62),
.B2(n_48),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_101),
.B1(n_103),
.B2(n_110),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_66),
.B1(n_55),
.B2(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_120),
.Y(n_134)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_82),
.C(n_83),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_107),
.Y(n_127)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_118),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_58),
.C(n_69),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_92),
.B1(n_91),
.B2(n_85),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_0),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_109),
.A2(n_114),
.B(n_102),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_56),
.B1(n_70),
.B2(n_59),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_84),
.B(n_90),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_57),
.B1(n_56),
.B2(n_68),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_95),
.B1(n_74),
.B2(n_85),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_26),
.B(n_20),
.Y(n_114)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_57),
.C(n_36),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_SL g182 ( 
.A(n_130),
.B(n_132),
.C(n_152),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_121),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_133),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_97),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_144),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_81),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_93),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_99),
.A2(n_94),
.B1(n_87),
.B2(n_85),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_94),
.B1(n_87),
.B2(n_95),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_110),
.B1(n_101),
.B2(n_119),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_153),
.A2(n_125),
.B(n_117),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_128),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_114),
.B(n_117),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_157),
.A2(n_174),
.B(n_179),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_105),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_169),
.C(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_152),
.B(n_109),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_177),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_127),
.C(n_153),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_103),
.B1(n_100),
.B2(n_112),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_171),
.B1(n_181),
.B2(n_128),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_103),
.B1(n_120),
.B2(n_98),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_107),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_103),
.B(n_109),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_175),
.B(n_147),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_141),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_59),
.C(n_49),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_133),
.C(n_131),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_79),
.B(n_103),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_79),
.B(n_20),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_104),
.B1(n_49),
.B2(n_44),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_192),
.B1(n_182),
.B2(n_175),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_185),
.B(n_189),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_135),
.B1(n_129),
.B2(n_127),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_186),
.A2(n_179),
.B1(n_174),
.B2(n_164),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_193),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_191),
.A2(n_203),
.B(n_205),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_171),
.A2(n_126),
.B1(n_146),
.B2(n_139),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_139),
.C(n_13),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_208),
.B1(n_26),
.B2(n_9),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_131),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_169),
.C(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_210),
.A2(n_219),
.B1(n_229),
.B2(n_235),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_218),
.C(n_222),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_170),
.B1(n_182),
.B2(n_165),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_227),
.B1(n_234),
.B2(n_191),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_217),
.A2(n_230),
.B(n_201),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_172),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_165),
.B1(n_168),
.B2(n_157),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_36),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_187),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_18),
.B1(n_26),
.B2(n_2),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_199),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_232),
.C(n_208),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_18),
.B1(n_26),
.B2(n_43),
.Y(n_229)
);

AND3x1_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_26),
.C(n_44),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_36),
.C(n_43),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_187),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_231),
.Y(n_238)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_239),
.B(n_254),
.Y(n_259)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_240),
.A2(n_243),
.B(n_244),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_203),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_246),
.Y(n_270)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_250),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_249),
.C(n_251),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_202),
.C(n_188),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_188),
.C(n_197),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_190),
.C(n_196),
.Y(n_252)
);

OAI322xp33_ASAP7_75t_L g265 ( 
.A1(n_252),
.A2(n_245),
.A3(n_240),
.B1(n_244),
.B2(n_258),
.C1(n_255),
.C2(n_236),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_255),
.Y(n_266)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_224),
.B(n_195),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_201),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_212),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_214),
.B1(n_210),
.B2(n_219),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_260),
.A2(n_266),
.B1(n_263),
.B2(n_267),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_224),
.B1(n_215),
.B2(n_217),
.Y(n_261)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

NOR4xp25_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_10),
.C(n_15),
.D(n_14),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_7),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_222),
.C(n_226),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_269),
.C(n_271),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_228),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_232),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_197),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_274),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_229),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_206),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_8),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_250),
.B(n_247),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_286),
.C(n_288),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_246),
.B(n_236),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_261),
.B(n_241),
.CI(n_235),
.CON(n_279),
.SN(n_279)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_289),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_272),
.A2(n_10),
.B(n_15),
.Y(n_281)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_287),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_8),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_264),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_16),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_285),
.C(n_280),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_263),
.A2(n_7),
.B(n_13),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_291),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_11),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_275),
.B1(n_274),
.B2(n_273),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_293),
.B(n_297),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_268),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_14),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_302),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_303),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_282),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_310),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_288),
.B1(n_280),
.B2(n_290),
.Y(n_309)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_282),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_12),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_313),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_12),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_4),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_5),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_299),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_321),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

NOR2x1p5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_293),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_323),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_301),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_316),
.B(n_322),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_327),
.B(n_5),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_306),
.Y(n_326)
);

XOR2x2_ASAP7_75t_SL g329 ( 
.A(n_326),
.B(n_304),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_304),
.B(n_5),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_324),
.B(n_328),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_5),
.B(n_6),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_6),
.B(n_305),
.Y(n_334)
);


endmodule