module fake_ariane_62_n_790 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_790);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_790;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_745;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_56),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_55),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

BUFx2_ASAP7_75t_SL g164 ( 
.A(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_26),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_101),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_47),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_34),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_32),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_109),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_17),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_4),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_57),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_92),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_11),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_74),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_69),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_43),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_95),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_124),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_133),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_27),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_20),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_94),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_41),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_127),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_149),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_40),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_24),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_118),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_60),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_15),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_23),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_84),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_122),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_107),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_90),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_29),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_9),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_148),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_110),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_0),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

AOI22x1_ASAP7_75t_SL g225 ( 
.A1(n_186),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_2),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_172),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_3),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_160),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_3),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_186),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_161),
.B(n_5),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_163),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_175),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_208),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_162),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_162),
.B(n_7),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_166),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_171),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_194),
.B(n_8),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_181),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_209),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_251),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_191),
.B1(n_165),
.B2(n_199),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_195),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_197),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_202),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_209),
.C(n_198),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_219),
.B(n_206),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_182),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_187),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_210),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_221),
.B(n_187),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_251),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_221),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_221),
.B(n_198),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_221),
.B(n_201),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_245),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_221),
.B(n_201),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_254),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_229),
.B(n_204),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_229),
.B(n_204),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_232),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_220),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_L g300 ( 
.A(n_230),
.B(n_214),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_229),
.B(n_215),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_236),
.B(n_200),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_232),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_234),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_228),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_L g307 ( 
.A(n_230),
.B(n_215),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_229),
.B(n_159),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_306),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_298),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_267),
.B(n_253),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_272),
.B(n_216),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_253),
.Y(n_315)
);

NAND3xp33_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_227),
.C(n_224),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_L g317 ( 
.A1(n_262),
.A2(n_239),
.B1(n_302),
.B2(n_240),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_274),
.B(n_223),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_223),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_300),
.A2(n_250),
.B1(n_255),
.B2(n_238),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_292),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_299),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_307),
.A2(n_238),
.B1(n_255),
.B2(n_246),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_273),
.B(n_238),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_286),
.B(n_241),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_249),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_305),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_274),
.B(n_241),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_274),
.A2(n_246),
.B1(n_243),
.B2(n_252),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_261),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_L g341 ( 
.A(n_292),
.B(n_237),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_274),
.B(n_174),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_260),
.B(n_225),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_306),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_176),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_286),
.B(n_244),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_289),
.B(n_297),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_288),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_266),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_L g350 ( 
.A(n_295),
.B(n_183),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_288),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_289),
.B(n_256),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_259),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_293),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_283),
.B(n_308),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_292),
.B(n_217),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_293),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_283),
.B(n_220),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_291),
.B(n_220),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_291),
.B(n_231),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_291),
.B(n_294),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_269),
.A2(n_290),
.B1(n_307),
.B2(n_279),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_294),
.B(n_218),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_264),
.B(n_242),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_282),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_271),
.B(n_231),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_265),
.B(n_242),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_285),
.A2(n_301),
.B1(n_296),
.B2(n_260),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_266),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_271),
.B(n_231),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_276),
.B(n_231),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_276),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_270),
.B(n_242),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_281),
.B(n_235),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_327),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_347),
.A2(n_281),
.B(n_287),
.Y(n_376)
);

NAND3xp33_ASAP7_75t_L g377 ( 
.A(n_311),
.B(n_287),
.C(n_299),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_309),
.B(n_299),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_311),
.B(n_268),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_315),
.A2(n_284),
.B(n_280),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_222),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_SL g382 ( 
.A(n_318),
.B(n_164),
.Y(n_382)
);

OAI21xp33_ASAP7_75t_L g383 ( 
.A1(n_321),
.A2(n_226),
.B(n_233),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_322),
.B(n_268),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_312),
.B(n_235),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_355),
.A2(n_284),
.B(n_280),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_329),
.A2(n_211),
.B1(n_192),
.B2(n_193),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_319),
.A2(n_277),
.B(n_275),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_330),
.A2(n_277),
.B(n_275),
.Y(n_390)
);

O2A1O1Ixp5_ASAP7_75t_L g391 ( 
.A1(n_318),
.A2(n_299),
.B(n_263),
.C(n_207),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_334),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_235),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_321),
.B(n_235),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_317),
.A2(n_190),
.B1(n_10),
.B2(n_11),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_317),
.A2(n_263),
.B1(n_10),
.B2(n_12),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

AOI21x1_ASAP7_75t_L g400 ( 
.A1(n_361),
.A2(n_263),
.B(n_80),
.Y(n_400)
);

AOI21x1_ASAP7_75t_L g401 ( 
.A1(n_359),
.A2(n_263),
.B(n_81),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_353),
.B(n_263),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_360),
.A2(n_350),
.B(n_345),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_316),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_14),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_L g406 ( 
.A1(n_342),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_358),
.A2(n_83),
.B(n_157),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_348),
.Y(n_408)
);

AOI21x1_ASAP7_75t_L g409 ( 
.A1(n_351),
.A2(n_82),
.B(n_155),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_354),
.B(n_16),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_362),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

OAI21xp33_ASAP7_75t_L g413 ( 
.A1(n_338),
.A2(n_18),
.B(n_19),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_352),
.B(n_158),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_328),
.A2(n_21),
.B(n_22),
.Y(n_415)
);

AOI21x1_ASAP7_75t_L g416 ( 
.A1(n_357),
.A2(n_310),
.B(n_313),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_342),
.A2(n_25),
.B(n_28),
.C(n_30),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

AND2x6_ASAP7_75t_SL g419 ( 
.A(n_343),
.B(n_31),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_320),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_314),
.B(n_33),
.Y(n_421)
);

O2A1O1Ixp33_ASAP7_75t_L g422 ( 
.A1(n_336),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_363),
.B(n_38),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_372),
.A2(n_39),
.B(n_42),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_363),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_341),
.A2(n_44),
.B(n_45),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_323),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_344),
.B(n_50),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_336),
.B(n_51),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_368),
.A2(n_331),
.B1(n_373),
.B2(n_364),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_328),
.A2(n_52),
.B(n_53),
.Y(n_433)
);

OAI21xp33_ASAP7_75t_SL g434 ( 
.A1(n_356),
.A2(n_54),
.B(n_58),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_364),
.B(n_59),
.Y(n_435)
);

OAI21xp33_ASAP7_75t_L g436 ( 
.A1(n_374),
.A2(n_61),
.B(n_62),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_369),
.Y(n_437)
);

BUFx4f_ASAP7_75t_L g438 ( 
.A(n_335),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_374),
.A2(n_63),
.B(n_65),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_367),
.B(n_154),
.Y(n_440)
);

O2A1O1Ixp5_ASAP7_75t_L g441 ( 
.A1(n_324),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_367),
.B(n_373),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_326),
.A2(n_71),
.B(n_72),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_365),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_399),
.Y(n_445)
);

AOI221x1_ASAP7_75t_L g446 ( 
.A1(n_411),
.A2(n_371),
.B1(n_370),
.B2(n_366),
.C(n_337),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_379),
.A2(n_337),
.B(n_75),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_387),
.B(n_73),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_76),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_77),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_375),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_420),
.B(n_78),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_416),
.A2(n_79),
.B(n_85),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_398),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_455)
);

A2O1A1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_413),
.A2(n_89),
.B(n_91),
.C(n_93),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_386),
.A2(n_97),
.B(n_98),
.Y(n_457)
);

A2O1A1Ixp33_ASAP7_75t_L g458 ( 
.A1(n_438),
.A2(n_395),
.B(n_439),
.C(n_432),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_390),
.A2(n_99),
.B(n_100),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_403),
.A2(n_102),
.B(n_104),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_381),
.B(n_106),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_383),
.B(n_108),
.Y(n_462)
);

NAND2x1p5_ASAP7_75t_L g463 ( 
.A(n_426),
.B(n_111),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_393),
.B(n_112),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_390),
.A2(n_113),
.B(n_114),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_395),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_392),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_410),
.Y(n_468)
);

AOI21x1_ASAP7_75t_L g469 ( 
.A1(n_414),
.A2(n_119),
.B(n_120),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_438),
.A2(n_125),
.B(n_128),
.C(n_130),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_394),
.B(n_131),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_388),
.B(n_132),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_389),
.A2(n_135),
.B(n_136),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_399),
.Y(n_475)
);

OAI21x1_ASAP7_75t_L g476 ( 
.A1(n_380),
.A2(n_376),
.B(n_400),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_405),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_410),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_402),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_391),
.A2(n_137),
.B(n_139),
.Y(n_480)
);

AO22x2_ASAP7_75t_L g481 ( 
.A1(n_411),
.A2(n_430),
.B1(n_427),
.B2(n_439),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_415),
.A2(n_140),
.B(n_141),
.Y(n_482)
);

AOI221x1_ASAP7_75t_L g483 ( 
.A1(n_436),
.A2(n_142),
.B1(n_144),
.B2(n_146),
.C(n_147),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_434),
.A2(n_151),
.B(n_153),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_424),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_401),
.A2(n_435),
.B(n_440),
.Y(n_486)
);

AO31x2_ASAP7_75t_L g487 ( 
.A1(n_417),
.A2(n_406),
.A3(n_423),
.B(n_385),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_424),
.B(n_404),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_409),
.A2(n_427),
.B(n_384),
.Y(n_489)
);

NOR4xp25_ASAP7_75t_L g490 ( 
.A(n_422),
.B(n_421),
.C(n_429),
.D(n_377),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_441),
.A2(n_407),
.B(n_425),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

AOI21x1_ASAP7_75t_SL g493 ( 
.A1(n_382),
.A2(n_378),
.B(n_428),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_397),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_418),
.B(n_437),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_424),
.B(n_433),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_443),
.A2(n_379),
.B(n_442),
.Y(n_497)
);

OA21x2_ASAP7_75t_L g498 ( 
.A1(n_419),
.A2(n_390),
.B(n_427),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_375),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g500 ( 
.A1(n_390),
.A2(n_427),
.B(n_439),
.Y(n_500)
);

AOI21x1_ASAP7_75t_L g501 ( 
.A1(n_416),
.A2(n_414),
.B(n_389),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_445),
.Y(n_502)
);

AO21x2_ASAP7_75t_L g503 ( 
.A1(n_480),
.A2(n_486),
.B(n_489),
.Y(n_503)
);

AO21x2_ASAP7_75t_L g504 ( 
.A1(n_480),
.A2(n_501),
.B(n_472),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_444),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_498),
.A2(n_481),
.B1(n_466),
.B2(n_455),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_458),
.B(n_468),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_453),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_494),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_497),
.A2(n_449),
.B(n_478),
.Y(n_510)
);

AO31x2_ASAP7_75t_L g511 ( 
.A1(n_446),
.A2(n_483),
.A3(n_455),
.B(n_456),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_498),
.A2(n_481),
.B1(n_466),
.B2(n_479),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_445),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_500),
.A2(n_492),
.B1(n_477),
.B2(n_467),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_499),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_445),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_495),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_475),
.B(n_463),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_476),
.A2(n_491),
.B(n_465),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_459),
.A2(n_482),
.B(n_457),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_495),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_470),
.B(n_464),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_474),
.A2(n_454),
.B(n_493),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_475),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_470),
.B(n_461),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_450),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_450),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_496),
.A2(n_460),
.B(n_447),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_470),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_449),
.B(n_488),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_485),
.B(n_500),
.Y(n_533)
);

AO31x2_ASAP7_75t_L g534 ( 
.A1(n_462),
.A2(n_452),
.A3(n_448),
.B(n_471),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_473),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_487),
.B(n_490),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_490),
.A2(n_484),
.B(n_469),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_484),
.B(n_487),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_L g539 ( 
.A1(n_487),
.A2(n_395),
.B1(n_411),
.B2(n_317),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_444),
.B(n_412),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_476),
.A2(n_501),
.B(n_491),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_470),
.Y(n_542)
);

OA21x2_ASAP7_75t_L g543 ( 
.A1(n_489),
.A2(n_476),
.B(n_446),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_453),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_453),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_453),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_445),
.B(n_475),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_445),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_444),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_532),
.A2(n_507),
.B(n_539),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_518),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_549),
.B(n_505),
.Y(n_552)
);

NAND2x1_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_527),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_522),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_547),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_536),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_508),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_544),
.B(n_546),
.Y(n_558)
);

OA21x2_ASAP7_75t_L g559 ( 
.A1(n_541),
.A2(n_537),
.B(n_510),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_540),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_545),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_512),
.B(n_506),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_533),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_523),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_524),
.A2(n_521),
.B(n_530),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_513),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_509),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_547),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_513),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_547),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_515),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_524),
.A2(n_521),
.B(n_530),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_539),
.B(n_512),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_514),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_531),
.B(n_548),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_523),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_514),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_506),
.B(n_523),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_528),
.Y(n_579)
);

BUFx2_ASAP7_75t_SL g580 ( 
.A(n_542),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_525),
.B(n_502),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_529),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_538),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_538),
.B(n_542),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_542),
.B(n_502),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_526),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_516),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_543),
.A2(n_520),
.B(n_503),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_535),
.A2(n_519),
.B1(n_516),
.B2(n_548),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_543),
.Y(n_590)
);

AO21x1_ASAP7_75t_L g591 ( 
.A1(n_535),
.A2(n_511),
.B(n_534),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_583),
.B(n_550),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_560),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_583),
.B(n_543),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_511),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_590),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_590),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_556),
.Y(n_598)
);

INVxp67_ASAP7_75t_SL g599 ( 
.A(n_553),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_584),
.B(n_511),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_567),
.Y(n_602)
);

NOR2x1_ASAP7_75t_L g603 ( 
.A(n_553),
.B(n_503),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_573),
.B(n_520),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_558),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_578),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_573),
.B(n_542),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_562),
.B(n_520),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_562),
.B(n_517),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_578),
.B(n_517),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_586),
.B(n_517),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_558),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_588),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_586),
.B(n_554),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_564),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_552),
.B(n_554),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_563),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_551),
.B(n_517),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_551),
.B(n_504),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_582),
.B(n_534),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_564),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_582),
.B(n_534),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_557),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_557),
.B(n_504),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_568),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_561),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_559),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_574),
.A2(n_534),
.B1(n_577),
.B2(n_571),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_561),
.B(n_579),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_569),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_555),
.B(n_570),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_579),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_591),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_575),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_566),
.B(n_555),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_591),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_559),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_605),
.B(n_587),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_612),
.B(n_576),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_599),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_602),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_616),
.B(n_576),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_608),
.B(n_559),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_623),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_598),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_629),
.B(n_555),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_634),
.B(n_593),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_598),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_608),
.B(n_559),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_630),
.B(n_581),
.Y(n_650)
);

OAI31xp33_ASAP7_75t_L g651 ( 
.A1(n_592),
.A2(n_607),
.A3(n_636),
.B(n_589),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_601),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_595),
.B(n_572),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_626),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_614),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_604),
.B(n_572),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_614),
.B(n_555),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_629),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_595),
.B(n_565),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_600),
.B(n_565),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_600),
.B(n_570),
.Y(n_661)
);

NOR2x1p5_ASAP7_75t_L g662 ( 
.A(n_635),
.B(n_570),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_632),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_615),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_604),
.B(n_570),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_601),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_617),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_624),
.B(n_585),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_619),
.B(n_585),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_631),
.B(n_585),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_619),
.B(n_585),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_632),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_617),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_603),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_645),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_645),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_648),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_653),
.B(n_606),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_653),
.B(n_606),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_659),
.B(n_636),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_659),
.B(n_597),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_668),
.B(n_610),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_641),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_640),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_668),
.B(n_610),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_SL g686 ( 
.A(n_650),
.B(n_621),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_648),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_660),
.B(n_596),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_664),
.B(n_655),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_647),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_644),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_652),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_660),
.B(n_597),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_661),
.B(n_597),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_661),
.B(n_637),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_656),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_642),
.B(n_618),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_640),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_652),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_643),
.B(n_649),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_643),
.B(n_649),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_654),
.B(n_618),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_669),
.B(n_637),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_638),
.B(n_609),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_669),
.B(n_637),
.Y(n_705)
);

NOR2x1_ASAP7_75t_L g706 ( 
.A(n_674),
.B(n_603),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_700),
.B(n_671),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_683),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_691),
.Y(n_709)
);

NAND2xp67_ASAP7_75t_L g710 ( 
.A(n_680),
.B(n_611),
.Y(n_710)
);

NAND2x2_ASAP7_75t_L g711 ( 
.A(n_689),
.B(n_662),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_675),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_675),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_676),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_700),
.B(n_671),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_686),
.A2(n_607),
.B1(n_609),
.B2(n_611),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_676),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_680),
.B(n_667),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_684),
.B(n_667),
.Y(n_719)
);

AND3x2_ASAP7_75t_L g720 ( 
.A(n_684),
.B(n_651),
.C(n_674),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_682),
.B(n_658),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_681),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_701),
.B(n_646),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_701),
.B(n_665),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_678),
.B(n_679),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_698),
.Y(n_726)
);

OR2x6_ASAP7_75t_L g727 ( 
.A(n_698),
.B(n_665),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_704),
.B(n_656),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_708),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_709),
.B(n_690),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_724),
.B(n_697),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_712),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_718),
.B(n_696),
.Y(n_733)
);

XOR2x2_ASAP7_75t_L g734 ( 
.A(n_720),
.B(n_716),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_711),
.A2(n_678),
.B1(n_679),
.B2(n_702),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_716),
.A2(n_657),
.B1(n_696),
.B2(n_685),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_726),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_718),
.B(n_696),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_713),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_719),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_740),
.B(n_719),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_734),
.A2(n_727),
.B(n_706),
.Y(n_742)
);

OAI322xp33_ASAP7_75t_L g743 ( 
.A1(n_730),
.A2(n_728),
.A3(n_714),
.B1(n_717),
.B2(n_687),
.C1(n_699),
.C2(n_692),
.Y(n_743)
);

OAI321xp33_ASAP7_75t_L g744 ( 
.A1(n_735),
.A2(n_720),
.A3(n_727),
.B1(n_633),
.B2(n_699),
.C(n_677),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_729),
.B(n_723),
.Y(n_745)
);

NOR2x1_ASAP7_75t_L g746 ( 
.A(n_732),
.B(n_726),
.Y(n_746)
);

AOI221xp5_ASAP7_75t_L g747 ( 
.A1(n_744),
.A2(n_735),
.B1(n_736),
.B2(n_739),
.C(n_738),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_741),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_743),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_L g750 ( 
.A(n_742),
.B(n_733),
.C(n_737),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_745),
.B(n_707),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_746),
.A2(n_693),
.B1(n_688),
.B2(n_681),
.Y(n_752)
);

NAND4xp25_ASAP7_75t_L g753 ( 
.A(n_749),
.B(n_725),
.C(n_687),
.D(n_677),
.Y(n_753)
);

OAI211xp5_ASAP7_75t_L g754 ( 
.A1(n_747),
.A2(n_750),
.B(n_748),
.C(n_752),
.Y(n_754)
);

NOR3x1_ASAP7_75t_L g755 ( 
.A(n_751),
.B(n_731),
.C(n_692),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_748),
.Y(n_756)
);

NAND2x1p5_ASAP7_75t_L g757 ( 
.A(n_751),
.B(n_721),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_754),
.B(n_639),
.C(n_706),
.Y(n_758)
);

AND3x1_ASAP7_75t_L g759 ( 
.A(n_756),
.B(n_715),
.C(n_722),
.Y(n_759)
);

XOR2x1_ASAP7_75t_L g760 ( 
.A(n_759),
.B(n_757),
.Y(n_760)
);

NOR2x1_ASAP7_75t_L g761 ( 
.A(n_758),
.B(n_753),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_758),
.B(n_755),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_761),
.B(n_721),
.Y(n_763)
);

NOR2x1p5_ASAP7_75t_L g764 ( 
.A(n_760),
.B(n_637),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_762),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_761),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_761),
.Y(n_767)
);

XNOR2x1_ASAP7_75t_L g768 ( 
.A(n_767),
.B(n_765),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_766),
.Y(n_769)
);

NAND4xp75_ASAP7_75t_L g770 ( 
.A(n_764),
.B(n_633),
.C(n_625),
.D(n_688),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_L g771 ( 
.A(n_763),
.B(n_622),
.C(n_620),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_SL g772 ( 
.A1(n_763),
.A2(n_727),
.B1(n_580),
.B2(n_625),
.Y(n_772)
);

OAI31xp33_ASAP7_75t_SL g773 ( 
.A1(n_767),
.A2(n_695),
.A3(n_705),
.B(n_703),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_769),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_768),
.B(n_705),
.Y(n_775)
);

NOR2xp67_ASAP7_75t_L g776 ( 
.A(n_772),
.B(n_666),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_771),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_773),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_774),
.B(n_770),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_778),
.A2(n_627),
.B1(n_666),
.B2(n_673),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_775),
.B(n_710),
.Y(n_781)
);

AO21x2_ASAP7_75t_L g782 ( 
.A1(n_776),
.A2(n_695),
.B(n_703),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_779),
.A2(n_776),
.B(n_777),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_780),
.A2(n_663),
.B(n_672),
.Y(n_784)
);

NAND2x1_ASAP7_75t_L g785 ( 
.A(n_781),
.B(n_627),
.Y(n_785)
);

AOI322xp5_ASAP7_75t_SL g786 ( 
.A1(n_783),
.A2(n_782),
.A3(n_621),
.B1(n_615),
.B2(n_670),
.C1(n_580),
.C2(n_694),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_784),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_787),
.A2(n_785),
.B1(n_627),
.B2(n_594),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_788),
.A2(n_786),
.B1(n_693),
.B2(n_627),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_789),
.A2(n_628),
.B1(n_594),
.B2(n_613),
.Y(n_790)
);


endmodule