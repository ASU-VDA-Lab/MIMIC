module fake_aes_8354_n_1280 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1280);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1280;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_411;
wire n_860;
wire n_1208;
wire n_1201;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_659;
wire n_432;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g350 ( .A(n_178), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_85), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_39), .Y(n_352) );
BUFx10_ASAP7_75t_L g353 ( .A(n_256), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_171), .B(n_183), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_189), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_28), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_242), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_54), .Y(n_358) );
NOR2xp67_ASAP7_75t_L g359 ( .A(n_209), .B(n_347), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_329), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_158), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_336), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_167), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_145), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_164), .Y(n_365) );
CKINVDCx16_ASAP7_75t_R g366 ( .A(n_160), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_35), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_332), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_226), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_44), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_131), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_341), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_198), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_205), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_249), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_240), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_308), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_12), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_63), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_293), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_126), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_82), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_138), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_105), .Y(n_384) );
CKINVDCx16_ASAP7_75t_R g385 ( .A(n_5), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_174), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_322), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_12), .Y(n_388) );
INVx4_ASAP7_75t_R g389 ( .A(n_140), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_142), .B(n_194), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_220), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_125), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_241), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_100), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_263), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_116), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_228), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_335), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_13), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_219), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_73), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_342), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_97), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_207), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_104), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_102), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_37), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_204), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_294), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_115), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_326), .Y(n_411) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_301), .B(n_309), .Y(n_412) );
NOR2xp67_ASAP7_75t_L g413 ( .A(n_258), .B(n_290), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_299), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_296), .Y(n_415) );
NOR2xp67_ASAP7_75t_L g416 ( .A(n_298), .B(n_225), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_41), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_330), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_268), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_344), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_208), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_187), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_87), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_34), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_285), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_191), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_80), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_90), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_265), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_143), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_147), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_4), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_118), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_89), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g435 ( .A(n_154), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_17), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_161), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_257), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_21), .Y(n_439) );
CKINVDCx16_ASAP7_75t_R g440 ( .A(n_1), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_182), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_278), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_323), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_23), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_292), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_37), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_151), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_98), .Y(n_448) );
INVxp33_ASAP7_75t_L g449 ( .A(n_244), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_114), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_233), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_180), .Y(n_452) );
INVxp67_ASAP7_75t_SL g453 ( .A(n_331), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_130), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_52), .Y(n_455) );
NOR2xp67_ASAP7_75t_L g456 ( .A(n_62), .B(n_181), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_314), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_259), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_138), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_311), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_26), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_130), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_221), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_327), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_264), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_253), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_246), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_173), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_312), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_98), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_255), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_224), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_67), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_169), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_125), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_109), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_109), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_230), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_105), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_126), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_150), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_176), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_261), .Y(n_483) );
NOR2xp67_ASAP7_75t_L g484 ( .A(n_124), .B(n_243), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_132), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_61), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_319), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_99), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_206), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_156), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_211), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_190), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_193), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_93), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_63), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_271), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_277), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_282), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_92), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_73), .Y(n_500) );
BUFx5_ASAP7_75t_L g501 ( .A(n_252), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_55), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_132), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_229), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_313), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_349), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_119), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_337), .Y(n_508) );
INVxp33_ASAP7_75t_SL g509 ( .A(n_234), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_43), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_120), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_78), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_5), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_76), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_55), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_338), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_273), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_272), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_86), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_197), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_284), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_33), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_210), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_157), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_280), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_15), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_320), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_289), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_339), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_212), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_67), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_175), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_64), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_152), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_162), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_46), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_163), .Y(n_537) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_279), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_172), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_25), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_288), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_19), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_72), .Y(n_543) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_227), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_501), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_503), .B(n_0), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_501), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_503), .B(n_0), .Y(n_548) );
AND2x6_ASAP7_75t_L g549 ( .A(n_517), .B(n_141), .Y(n_549) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_372), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_403), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_403), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_405), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_372), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_449), .B(n_2), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_385), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_556) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_372), .Y(n_557) );
BUFx3_ASAP7_75t_L g558 ( .A(n_517), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_478), .B(n_3), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_384), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_501), .Y(n_561) );
OAI21x1_ASAP7_75t_L g562 ( .A1(n_364), .A2(n_146), .B(n_144), .Y(n_562) );
INVx3_ASAP7_75t_L g563 ( .A(n_353), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_405), .Y(n_564) );
AOI22x1_ASAP7_75t_SL g565 ( .A1(n_358), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_356), .B(n_6), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_365), .B(n_7), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_501), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_440), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_569) );
NAND2xp33_ASAP7_75t_L g570 ( .A(n_501), .B(n_148), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_501), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_353), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_356), .B(n_9), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_366), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_455), .B(n_10), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_406), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_435), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_501), .Y(n_578) );
BUFx3_ASAP7_75t_L g579 ( .A(n_364), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_538), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_382), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_372), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_361), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_455), .Y(n_584) );
AND2x6_ASAP7_75t_L g585 ( .A(n_368), .B(n_149), .Y(n_585) );
BUFx12f_ASAP7_75t_L g586 ( .A(n_353), .Y(n_586) );
AND2x4_ASAP7_75t_L g587 ( .A(n_500), .B(n_11), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_550), .Y(n_588) );
BUFx3_ASAP7_75t_L g589 ( .A(n_558), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_558), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_563), .B(n_544), .Y(n_591) );
AO22x2_ASAP7_75t_L g592 ( .A1(n_565), .A2(n_376), .B1(n_380), .B2(n_368), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_550), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_563), .B(n_449), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_550), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_563), .B(n_500), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_545), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_545), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_546), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_550), .Y(n_600) );
AND3x2_ASAP7_75t_L g601 ( .A(n_560), .B(n_453), .C(n_391), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_547), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_563), .B(n_363), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_572), .B(n_502), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_576), .B(n_461), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_572), .B(n_376), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_572), .B(n_380), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_547), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_572), .B(n_558), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_547), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_561), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_546), .B(n_429), .Y(n_612) );
INVx2_ASAP7_75t_SL g613 ( .A(n_549), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_555), .A2(n_488), .B1(n_386), .B2(n_419), .Y(n_614) );
BUFx3_ASAP7_75t_L g615 ( .A(n_549), .Y(n_615) );
INVx3_ASAP7_75t_L g616 ( .A(n_546), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_550), .Y(n_617) );
INVx6_ASAP7_75t_L g618 ( .A(n_546), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_561), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_555), .B(n_429), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_579), .B(n_441), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_575), .A2(n_367), .B1(n_370), .B2(n_351), .Y(n_622) );
BUFx3_ASAP7_75t_L g623 ( .A(n_549), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_550), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_587), .A2(n_392), .B1(n_394), .B2(n_378), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_587), .A2(n_401), .B1(n_417), .B2(n_399), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_554), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_561), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_594), .B(n_586), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_620), .B(n_581), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_620), .B(n_586), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_615), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_596), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_591), .B(n_586), .Y(n_634) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_615), .Y(n_635) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_605), .B(n_556), .C(n_559), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_605), .Y(n_637) );
BUFx12f_ASAP7_75t_L g638 ( .A(n_605), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_597), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_599), .B(n_566), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_603), .B(n_559), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_597), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g643 ( .A(n_614), .B(n_556), .C(n_569), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_596), .Y(n_644) );
INVxp67_ASAP7_75t_L g645 ( .A(n_614), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_603), .B(n_596), .Y(n_646) );
NOR2xp33_ASAP7_75t_SL g647 ( .A(n_615), .B(n_361), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_604), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_599), .B(n_566), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_613), .A2(n_562), .B(n_568), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_618), .A2(n_566), .B1(n_573), .B2(n_548), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_618), .A2(n_575), .B1(n_587), .B2(n_566), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_604), .B(n_548), .Y(n_653) );
OR2x6_ASAP7_75t_L g654 ( .A(n_592), .B(n_567), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_604), .B(n_567), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_589), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_599), .B(n_573), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_612), .A2(n_587), .B(n_575), .C(n_552), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_606), .B(n_607), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_618), .Y(n_660) );
NOR2xp67_ASAP7_75t_L g661 ( .A(n_606), .B(n_574), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_618), .B(n_548), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_607), .B(n_548), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_618), .A2(n_573), .B1(n_580), .B2(n_577), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_590), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_622), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_609), .B(n_573), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_599), .B(n_575), .Y(n_668) );
BUFx8_ASAP7_75t_L g669 ( .A(n_592), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_609), .B(n_579), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_622), .B(n_583), .Y(n_671) );
HB1xp67_ASAP7_75t_SL g672 ( .A(n_592), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_616), .B(n_579), .Y(n_673) );
INVx4_ASAP7_75t_L g674 ( .A(n_616), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_590), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_625), .A2(n_583), .B1(n_419), .B2(n_468), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_623), .B(n_568), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_625), .A2(n_468), .B1(n_482), .B2(n_386), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_612), .B(n_509), .Y(n_679) );
INVx8_ASAP7_75t_L g680 ( .A(n_626), .Y(n_680) );
AOI22xp5_ASAP7_75t_SL g681 ( .A1(n_592), .A2(n_358), .B1(n_514), .B2(n_410), .Y(n_681) );
INVx3_ASAP7_75t_L g682 ( .A(n_598), .Y(n_682) );
CKINVDCx8_ASAP7_75t_R g683 ( .A(n_592), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_598), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_601), .B(n_382), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_601), .A2(n_569), .B1(n_482), .B2(n_516), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_621), .A2(n_508), .B1(n_516), .B2(n_383), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_602), .A2(n_585), .B1(n_549), .B2(n_571), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_602), .B(n_509), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_608), .B(n_551), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_610), .B(n_611), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_610), .B(n_551), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_611), .B(n_552), .Y(n_693) );
NOR2xp33_ASAP7_75t_SL g694 ( .A(n_623), .B(n_508), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_619), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_628), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_613), .B(n_553), .Y(n_697) );
AND2x2_ASAP7_75t_SL g698 ( .A(n_613), .B(n_570), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_588), .B(n_564), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_588), .B(n_564), .Y(n_700) );
INVx3_ASAP7_75t_L g701 ( .A(n_588), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_593), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_593), .A2(n_585), .B1(n_549), .B2(n_571), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_640), .A2(n_562), .B(n_568), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_652), .A2(n_526), .B1(n_542), .B2(n_514), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_655), .B(n_383), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_652), .A2(n_542), .B1(n_526), .B2(n_427), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_682), .Y(n_708) );
OAI21x1_ASAP7_75t_L g709 ( .A1(n_650), .A2(n_578), .B(n_354), .Y(n_709) );
CKINVDCx8_ASAP7_75t_R g710 ( .A(n_654), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_659), .B(n_352), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_672), .A2(n_433), .B1(n_434), .B2(n_423), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_641), .B(n_371), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_637), .B(n_565), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_637), .B(n_396), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_644), .Y(n_716) );
O2A1O1Ixp33_ASAP7_75t_L g717 ( .A1(n_630), .A2(n_439), .B(n_444), .C(n_436), .Y(n_717) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_687), .Y(n_718) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_678), .Y(n_719) );
NOR2xp33_ASAP7_75t_SL g720 ( .A(n_647), .B(n_549), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_636), .B(n_499), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_649), .A2(n_360), .B(n_350), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_674), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_680), .A2(n_585), .B1(n_549), .B2(n_459), .Y(n_724) );
INVx3_ASAP7_75t_SL g725 ( .A(n_681), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_646), .B(n_379), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_657), .A2(n_387), .B(n_373), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_653), .B(n_381), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_636), .A2(n_407), .B1(n_424), .B2(n_388), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_651), .A2(n_462), .B1(n_473), .B2(n_446), .Y(n_730) );
INVx4_ASAP7_75t_L g731 ( .A(n_680), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_694), .B(n_355), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_632), .B(n_357), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_653), .B(n_648), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_657), .A2(n_397), .B(n_395), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_677), .A2(n_408), .B(n_404), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_680), .A2(n_585), .B1(n_476), .B2(n_477), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_632), .B(n_362), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_691), .Y(n_739) );
OAI22x1_ASAP7_75t_L g740 ( .A1(n_686), .A2(n_432), .B1(n_448), .B2(n_428), .Y(n_740) );
O2A1O1Ixp5_ASAP7_75t_L g741 ( .A1(n_668), .A2(n_662), .B(n_679), .C(n_663), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_679), .B(n_450), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_643), .A2(n_654), .B1(n_666), .B2(n_671), .Y(n_743) );
BUFx8_ASAP7_75t_L g744 ( .A(n_685), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_632), .B(n_369), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_683), .A2(n_475), .B1(n_494), .B2(n_480), .Y(n_746) );
NAND2xp33_ASAP7_75t_L g747 ( .A(n_632), .B(n_585), .Y(n_747) );
OAI22x1_ASAP7_75t_L g748 ( .A1(n_645), .A2(n_470), .B1(n_485), .B2(n_454), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_676), .B(n_512), .Y(n_749) );
INVx4_ASAP7_75t_L g750 ( .A(n_674), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_L g751 ( .A1(n_643), .A2(n_511), .B(n_513), .C(n_510), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_677), .A2(n_411), .B(n_409), .Y(n_752) );
INVxp67_ASAP7_75t_L g753 ( .A(n_689), .Y(n_753) );
O2A1O1Ixp33_ASAP7_75t_L g754 ( .A1(n_658), .A2(n_522), .B(n_531), .C(n_515), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_667), .A2(n_418), .B(n_415), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_634), .A2(n_495), .B1(n_519), .B2(n_486), .Y(n_756) );
INVx4_ASAP7_75t_L g757 ( .A(n_639), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_654), .B(n_536), .Y(n_758) );
INVx1_ASAP7_75t_SL g759 ( .A(n_642), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_642), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_634), .B(n_543), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_629), .B(n_533), .Y(n_762) );
INVx1_ASAP7_75t_SL g763 ( .A(n_684), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_697), .A2(n_421), .B(n_420), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_629), .B(n_584), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_662), .B(n_540), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_688), .B(n_479), .C(n_502), .Y(n_767) );
INVxp67_ASAP7_75t_L g768 ( .A(n_690), .Y(n_768) );
O2A1O1Ixp33_ASAP7_75t_SL g769 ( .A1(n_673), .A2(n_426), .B(n_430), .C(n_422), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_669), .A2(n_585), .B1(n_479), .B2(n_507), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_670), .A2(n_437), .B(n_431), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_669), .A2(n_585), .B1(n_479), .B2(n_447), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_698), .A2(n_452), .B(n_451), .Y(n_773) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_635), .Y(n_774) );
INVx6_ASAP7_75t_L g775 ( .A(n_635), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_692), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_695), .A2(n_479), .B1(n_457), .B2(n_465), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_690), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_664), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_660), .B(n_374), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_696), .B(n_375), .Y(n_781) );
AOI21x1_ASAP7_75t_L g782 ( .A1(n_699), .A2(n_600), .B(n_595), .Y(n_782) );
NAND2x1p5_ASAP7_75t_L g783 ( .A(n_635), .B(n_456), .Y(n_783) );
OAI21xp33_ASAP7_75t_L g784 ( .A1(n_693), .A2(n_402), .B(n_393), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_698), .B(n_414), .Y(n_785) );
AND2x4_ASAP7_75t_L g786 ( .A(n_656), .B(n_484), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_700), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g788 ( .A(n_635), .B(n_425), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_665), .A2(n_467), .B(n_460), .Y(n_789) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_675), .Y(n_790) );
AO21x1_ASAP7_75t_L g791 ( .A1(n_702), .A2(n_472), .B(n_469), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_688), .A2(n_489), .B1(n_497), .B2(n_487), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_701), .Y(n_793) );
AOI21x1_ASAP7_75t_L g794 ( .A1(n_703), .A2(n_617), .B(n_600), .Y(n_794) );
A2O1A1Ixp33_ASAP7_75t_L g795 ( .A1(n_662), .A2(n_505), .B(n_518), .C(n_504), .Y(n_795) );
A2O1A1Ixp33_ASAP7_75t_L g796 ( .A1(n_662), .A2(n_523), .B(n_524), .C(n_520), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_682), .Y(n_797) );
AOI21xp33_ASAP7_75t_L g798 ( .A1(n_631), .A2(n_438), .B(n_400), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_637), .B(n_443), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_633), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g801 ( .A1(n_640), .A2(n_528), .B(n_525), .Y(n_801) );
NOR2x1_ASAP7_75t_L g802 ( .A(n_661), .B(n_529), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_640), .A2(n_534), .B(n_530), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_633), .B(n_535), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_640), .A2(n_541), .B(n_537), .Y(n_805) );
INVx3_ASAP7_75t_L g806 ( .A(n_682), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_637), .B(n_442), .Y(n_807) );
BUFx12f_ASAP7_75t_L g808 ( .A(n_638), .Y(n_808) );
OAI221xp5_ASAP7_75t_L g809 ( .A1(n_636), .A2(n_498), .B1(n_521), .B2(n_492), .C(n_464), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g810 ( .A1(n_640), .A2(n_492), .B(n_464), .Y(n_810) );
AND2x4_ASAP7_75t_L g811 ( .A(n_633), .B(n_359), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_637), .B(n_445), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_633), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_776), .B(n_463), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_739), .B(n_466), .Y(n_815) );
BUFx3_ASAP7_75t_L g816 ( .A(n_808), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_704), .A2(n_627), .B(n_624), .Y(n_817) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_705), .Y(n_818) );
OAI21x1_ASAP7_75t_L g819 ( .A1(n_794), .A2(n_521), .B(n_498), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_779), .B(n_471), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_705), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_773), .A2(n_627), .B(n_390), .Y(n_822) );
AO31x2_ASAP7_75t_L g823 ( .A1(n_791), .A2(n_582), .A3(n_390), .B(n_627), .Y(n_823) );
AOI31xp67_ASAP7_75t_L g824 ( .A1(n_809), .A2(n_582), .A3(n_413), .B(n_416), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_759), .A2(n_412), .B(n_474), .Y(n_825) );
O2A1O1Ixp33_ASAP7_75t_L g826 ( .A1(n_717), .A2(n_389), .B(n_16), .C(n_14), .Y(n_826) );
A2O1A1Ixp33_ASAP7_75t_L g827 ( .A1(n_741), .A2(n_398), .B(n_458), .C(n_377), .Y(n_827) );
AOI21xp33_ASAP7_75t_L g828 ( .A1(n_807), .A2(n_483), .B(n_481), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_768), .B(n_490), .Y(n_829) );
OR2x2_ASAP7_75t_L g830 ( .A(n_707), .B(n_14), .Y(n_830) );
NAND2xp5_ASAP7_75t_SL g831 ( .A(n_759), .B(n_491), .Y(n_831) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_707), .Y(n_832) );
OAI21xp5_ASAP7_75t_L g833 ( .A1(n_709), .A2(n_496), .B(n_493), .Y(n_833) );
OAI21x1_ASAP7_75t_L g834 ( .A1(n_782), .A2(n_398), .B(n_377), .Y(n_834) );
AOI21xp33_ASAP7_75t_L g835 ( .A1(n_812), .A2(n_527), .B(n_506), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_763), .A2(n_539), .B(n_532), .Y(n_836) );
AO22x2_ASAP7_75t_L g837 ( .A1(n_712), .A2(n_17), .B1(n_15), .B2(n_16), .Y(n_837) );
CKINVDCx5p33_ASAP7_75t_R g838 ( .A(n_744), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_716), .Y(n_839) );
BUFx3_ASAP7_75t_L g840 ( .A(n_744), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_757), .Y(n_841) );
NAND2x1p5_ASAP7_75t_L g842 ( .A(n_750), .B(n_458), .Y(n_842) );
AND2x4_ASAP7_75t_L g843 ( .A(n_800), .B(n_18), .Y(n_843) );
OAI21xp5_ASAP7_75t_L g844 ( .A1(n_767), .A2(n_557), .B(n_554), .Y(n_844) );
OR2x2_ASAP7_75t_L g845 ( .A(n_715), .B(n_18), .Y(n_845) );
BUFx10_ASAP7_75t_L g846 ( .A(n_811), .Y(n_846) );
OAI21x1_ASAP7_75t_L g847 ( .A1(n_783), .A2(n_557), .B(n_554), .Y(n_847) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_725), .Y(n_848) );
AOI21xp5_ASAP7_75t_L g849 ( .A1(n_747), .A2(n_557), .B(n_153), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_720), .A2(n_159), .B(n_155), .Y(n_850) );
AOI221x1_ASAP7_75t_L g851 ( .A1(n_712), .A2(n_19), .B1(n_20), .B2(n_21), .C(n_22), .Y(n_851) );
INVx3_ASAP7_75t_L g852 ( .A(n_750), .Y(n_852) );
AOI21x1_ASAP7_75t_SL g853 ( .A1(n_766), .A2(n_166), .B(n_165), .Y(n_853) );
AO31x2_ASAP7_75t_L g854 ( .A1(n_792), .A2(n_23), .A3(n_20), .B(n_22), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_714), .A2(n_26), .B1(n_24), .B2(n_25), .Y(n_855) );
AO21x1_ASAP7_75t_L g856 ( .A1(n_720), .A2(n_170), .B(n_168), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_746), .A2(n_28), .B1(n_24), .B2(n_27), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_718), .B(n_721), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_813), .Y(n_859) );
OAI21x1_ASAP7_75t_L g860 ( .A1(n_810), .A2(n_179), .B(n_177), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_760), .Y(n_861) );
O2A1O1Ixp33_ASAP7_75t_L g862 ( .A1(n_795), .A2(n_30), .B(n_27), .C(n_29), .Y(n_862) );
A2O1A1Ixp33_ASAP7_75t_L g863 ( .A1(n_754), .A2(n_31), .B(n_29), .C(n_30), .Y(n_863) );
AND2x4_ASAP7_75t_L g864 ( .A(n_731), .B(n_31), .Y(n_864) );
CKINVDCx11_ASAP7_75t_R g865 ( .A(n_710), .Y(n_865) );
NAND2x1p5_ASAP7_75t_L g866 ( .A(n_723), .B(n_32), .Y(n_866) );
OAI21xp5_ASAP7_75t_L g867 ( .A1(n_755), .A2(n_185), .B(n_184), .Y(n_867) );
BUFx6f_ASAP7_75t_L g868 ( .A(n_774), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_753), .B(n_32), .Y(n_869) );
A2O1A1Ixp33_ASAP7_75t_L g870 ( .A1(n_762), .A2(n_35), .B(n_33), .C(n_34), .Y(n_870) );
NOR2x1_ASAP7_75t_SL g871 ( .A(n_731), .B(n_36), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_719), .B(n_36), .Y(n_872) );
AO31x2_ASAP7_75t_L g873 ( .A1(n_792), .A2(n_40), .A3(n_38), .B(n_39), .Y(n_873) );
AO31x2_ASAP7_75t_L g874 ( .A1(n_796), .A2(n_41), .A3(n_38), .B(n_40), .Y(n_874) );
NOR2xp33_ASAP7_75t_SL g875 ( .A(n_746), .B(n_42), .Y(n_875) );
OAI21x1_ASAP7_75t_L g876 ( .A1(n_724), .A2(n_188), .B(n_186), .Y(n_876) );
OAI21xp5_ASAP7_75t_L g877 ( .A1(n_722), .A2(n_195), .B(n_192), .Y(n_877) );
AOI21xp5_ASAP7_75t_L g878 ( .A1(n_713), .A2(n_199), .B(n_196), .Y(n_878) );
OAI21xp5_ASAP7_75t_L g879 ( .A1(n_727), .A2(n_201), .B(n_200), .Y(n_879) );
O2A1O1Ixp33_ASAP7_75t_L g880 ( .A1(n_751), .A2(n_44), .B(n_42), .C(n_43), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_743), .A2(n_48), .B1(n_45), .B2(n_47), .Y(n_881) );
INVx2_ASAP7_75t_SL g882 ( .A(n_804), .Y(n_882) );
OAI21xp5_ASAP7_75t_L g883 ( .A1(n_735), .A2(n_203), .B(n_202), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_711), .B(n_49), .Y(n_884) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_774), .Y(n_885) );
OA21x2_ASAP7_75t_L g886 ( .A1(n_737), .A2(n_752), .B(n_736), .Y(n_886) );
INVx8_ASAP7_75t_L g887 ( .A(n_804), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_758), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_734), .B(n_50), .Y(n_889) );
NOR2xp67_ASAP7_75t_L g890 ( .A(n_748), .B(n_51), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_765), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_787), .Y(n_892) );
NAND2x1p5_ASAP7_75t_L g893 ( .A(n_806), .B(n_53), .Y(n_893) );
O2A1O1Ixp33_ASAP7_75t_L g894 ( .A1(n_730), .A2(n_53), .B(n_54), .C(n_56), .Y(n_894) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_729), .B(n_56), .Y(n_895) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_799), .B(n_57), .Y(n_896) );
INVx4_ASAP7_75t_L g897 ( .A(n_806), .Y(n_897) );
AO21x1_ASAP7_75t_L g898 ( .A1(n_786), .A2(n_214), .B(n_213), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_749), .B(n_57), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_811), .Y(n_900) );
AO31x2_ASAP7_75t_L g901 ( .A1(n_730), .A2(n_58), .A3(n_59), .B(n_60), .Y(n_901) );
A2O1A1Ixp33_ASAP7_75t_L g902 ( .A1(n_778), .A2(n_58), .B(n_59), .C(n_60), .Y(n_902) );
OAI21xp5_ASAP7_75t_L g903 ( .A1(n_801), .A2(n_216), .B(n_215), .Y(n_903) );
AOI21xp5_ASAP7_75t_L g904 ( .A1(n_793), .A2(n_218), .B(n_217), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_740), .A2(n_62), .B1(n_65), .B2(n_66), .Y(n_905) );
A2O1A1Ixp33_ASAP7_75t_L g906 ( .A1(n_771), .A2(n_65), .B(n_66), .C(n_68), .Y(n_906) );
AOI31xp67_ASAP7_75t_L g907 ( .A1(n_708), .A2(n_237), .A3(n_346), .B(n_345), .Y(n_907) );
HB1xp67_ASAP7_75t_L g908 ( .A(n_706), .Y(n_908) );
AO31x2_ASAP7_75t_L g909 ( .A1(n_803), .A2(n_68), .A3(n_69), .B(n_70), .Y(n_909) );
OAI21x1_ASAP7_75t_L g910 ( .A1(n_797), .A2(n_223), .B(n_222), .Y(n_910) );
OAI21xp5_ASAP7_75t_L g911 ( .A1(n_805), .A2(n_764), .B(n_789), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_756), .B(n_69), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_726), .B(n_70), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_742), .A2(n_71), .B1(n_72), .B2(n_74), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_785), .A2(n_232), .B(n_231), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_728), .B(n_71), .Y(n_916) );
O2A1O1Ixp5_ASAP7_75t_L g917 ( .A1(n_732), .A2(n_248), .B(n_343), .C(n_340), .Y(n_917) );
A2O1A1Ixp33_ASAP7_75t_L g918 ( .A1(n_781), .A2(n_74), .B(n_75), .C(n_76), .Y(n_918) );
OAI21x1_ASAP7_75t_L g919 ( .A1(n_733), .A2(n_236), .B(n_235), .Y(n_919) );
BUFx6f_ASAP7_75t_L g920 ( .A(n_775), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_775), .Y(n_921) );
OAI21x1_ASAP7_75t_L g922 ( .A1(n_738), .A2(n_239), .B(n_238), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_769), .Y(n_923) );
INVxp67_ASAP7_75t_L g924 ( .A(n_802), .Y(n_924) );
BUFx6f_ASAP7_75t_L g925 ( .A(n_790), .Y(n_925) );
AOI221x1_ASAP7_75t_L g926 ( .A1(n_798), .A2(n_75), .B1(n_77), .B2(n_78), .C(n_79), .Y(n_926) );
AO31x2_ASAP7_75t_L g927 ( .A1(n_780), .A2(n_77), .A3(n_79), .B(n_80), .Y(n_927) );
OA21x2_ASAP7_75t_L g928 ( .A1(n_770), .A2(n_262), .B(n_334), .Y(n_928) );
AO32x2_ASAP7_75t_L g929 ( .A1(n_772), .A2(n_81), .A3(n_82), .B1(n_83), .B2(n_84), .Y(n_929) );
BUFx6f_ASAP7_75t_L g930 ( .A(n_790), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_761), .Y(n_931) );
OAI21x1_ASAP7_75t_L g932 ( .A1(n_745), .A2(n_266), .B(n_333), .Y(n_932) );
NAND2x1p5_ASAP7_75t_L g933 ( .A(n_790), .B(n_83), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_777), .A2(n_84), .B1(n_85), .B2(n_86), .Y(n_934) );
OAI21xp5_ASAP7_75t_L g935 ( .A1(n_788), .A2(n_269), .B(n_328), .Y(n_935) );
NAND2x1p5_ASAP7_75t_L g936 ( .A(n_784), .B(n_88), .Y(n_936) );
AND2x4_ASAP7_75t_L g937 ( .A(n_739), .B(n_90), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_757), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_779), .B(n_91), .Y(n_939) );
AO31x2_ASAP7_75t_L g940 ( .A1(n_791), .A2(n_92), .A3(n_93), .B(n_94), .Y(n_940) );
AO32x2_ASAP7_75t_L g941 ( .A1(n_712), .A2(n_94), .A3(n_95), .B1(n_96), .B2(n_97), .Y(n_941) );
AO31x2_ASAP7_75t_L g942 ( .A1(n_791), .A2(n_95), .A3(n_96), .B(n_99), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_776), .Y(n_943) );
OR2x2_ASAP7_75t_L g944 ( .A(n_705), .B(n_100), .Y(n_944) );
AO31x2_ASAP7_75t_L g945 ( .A1(n_791), .A2(n_101), .A3(n_102), .B(n_103), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_707), .A2(n_101), .B1(n_103), .B2(n_104), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_776), .B(n_106), .Y(n_947) );
NOR2xp33_ASAP7_75t_L g948 ( .A(n_779), .B(n_107), .Y(n_948) );
AO21x2_ASAP7_75t_L g949 ( .A1(n_709), .A2(n_283), .B(n_325), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_818), .A2(n_107), .B1(n_108), .B2(n_110), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_892), .Y(n_951) );
OAI22x1_ASAP7_75t_L g952 ( .A1(n_937), .A2(n_110), .B1(n_111), .B2(n_112), .Y(n_952) );
CKINVDCx11_ASAP7_75t_R g953 ( .A(n_816), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_861), .Y(n_954) );
BUFx2_ASAP7_75t_L g955 ( .A(n_887), .Y(n_955) );
INVx3_ASAP7_75t_L g956 ( .A(n_897), .Y(n_956) );
AO21x2_ASAP7_75t_L g957 ( .A1(n_827), .A2(n_281), .B(n_324), .Y(n_957) );
OAI21xp5_ASAP7_75t_L g958 ( .A1(n_858), .A2(n_111), .B(n_112), .Y(n_958) );
A2O1A1Ixp33_ASAP7_75t_L g959 ( .A1(n_826), .A2(n_113), .B(n_114), .C(n_115), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_839), .Y(n_960) );
BUFx3_ASAP7_75t_L g961 ( .A(n_840), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_891), .B(n_113), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_908), .B(n_116), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_832), .B(n_117), .Y(n_964) );
A2O1A1Ixp33_ASAP7_75t_L g965 ( .A1(n_931), .A2(n_118), .B(n_119), .C(n_120), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_859), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_843), .Y(n_967) );
OAI21x1_ASAP7_75t_SL g968 ( .A1(n_871), .A2(n_121), .B(n_122), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_837), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_916), .B(n_122), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_837), .Y(n_971) );
AO21x2_ASAP7_75t_L g972 ( .A1(n_833), .A2(n_287), .B(n_321), .Y(n_972) );
OAI21x1_ASAP7_75t_L g973 ( .A1(n_853), .A2(n_286), .B(n_318), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_944), .Y(n_974) );
AOI21xp5_ASAP7_75t_L g975 ( .A1(n_911), .A2(n_276), .B(n_317), .Y(n_975) );
A2O1A1Ixp33_ASAP7_75t_L g976 ( .A1(n_896), .A2(n_123), .B(n_124), .C(n_127), .Y(n_976) );
OA21x2_ASAP7_75t_L g977 ( .A1(n_844), .A2(n_275), .B(n_316), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_872), .B(n_123), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_884), .B(n_127), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_913), .B(n_889), .Y(n_980) );
AND2x4_ASAP7_75t_L g981 ( .A(n_852), .B(n_128), .Y(n_981) );
INVx2_ASAP7_75t_SL g982 ( .A(n_838), .Y(n_982) );
OAI21x1_ASAP7_75t_SL g983 ( .A1(n_898), .A2(n_128), .B(n_129), .Y(n_983) );
AO21x2_ASAP7_75t_L g984 ( .A1(n_949), .A2(n_291), .B(n_315), .Y(n_984) );
NAND2x1p5_ASAP7_75t_L g985 ( .A(n_864), .B(n_131), .Y(n_985) );
OR2x2_ASAP7_75t_L g986 ( .A(n_845), .B(n_133), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_830), .Y(n_987) );
AOI21xp33_ASAP7_75t_SL g988 ( .A1(n_848), .A2(n_133), .B(n_134), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_866), .Y(n_989) );
NOR3xp33_ASAP7_75t_L g990 ( .A(n_880), .B(n_134), .C(n_135), .Y(n_990) );
AOI22xp5_ASAP7_75t_L g991 ( .A1(n_875), .A2(n_135), .B1(n_136), .B2(n_137), .Y(n_991) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_882), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_899), .B(n_136), .Y(n_993) );
CKINVDCx11_ASAP7_75t_R g994 ( .A(n_846), .Y(n_994) );
OAI21x1_ASAP7_75t_L g995 ( .A1(n_847), .A2(n_274), .B(n_310), .Y(n_995) );
BUFx8_ASAP7_75t_SL g996 ( .A(n_900), .Y(n_996) );
OR2x2_ASAP7_75t_L g997 ( .A(n_814), .B(n_139), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_895), .B(n_139), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_947), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_869), .A2(n_245), .B1(n_247), .B2(n_250), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_923), .B(n_251), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_912), .B(n_348), .Y(n_1002) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_893), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_946), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_841), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_901), .Y(n_1006) );
AOI21xp5_ASAP7_75t_L g1007 ( .A1(n_822), .A2(n_254), .B(n_260), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_901), .Y(n_1008) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_938), .B(n_267), .Y(n_1009) );
CKINVDCx11_ASAP7_75t_R g1010 ( .A(n_865), .Y(n_1010) );
OA21x2_ASAP7_75t_L g1011 ( .A1(n_910), .A2(n_270), .B(n_295), .Y(n_1011) );
A2O1A1Ixp33_ASAP7_75t_L g1012 ( .A1(n_862), .A2(n_297), .B(n_300), .C(n_302), .Y(n_1012) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_890), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_874), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_857), .A2(n_303), .B1(n_304), .B2(n_305), .Y(n_1015) );
AO21x2_ASAP7_75t_L g1016 ( .A1(n_867), .A2(n_306), .B(n_307), .Y(n_1016) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_820), .B(n_924), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_933), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_815), .B(n_823), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_874), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_874), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_909), .Y(n_1022) );
BUFx3_ASAP7_75t_L g1023 ( .A(n_920), .Y(n_1023) );
OR2x6_ASAP7_75t_L g1024 ( .A(n_842), .B(n_894), .Y(n_1024) );
A2O1A1Ixp33_ASAP7_75t_L g1025 ( .A1(n_863), .A2(n_918), .B(n_870), .C(n_906), .Y(n_1025) );
AOI22xp33_ASAP7_75t_SL g1026 ( .A1(n_939), .A2(n_948), .B1(n_881), .B2(n_936), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_823), .B(n_886), .Y(n_1027) );
A2O1A1Ixp33_ASAP7_75t_L g1028 ( .A1(n_905), .A2(n_902), .B(n_825), .C(n_915), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_823), .B(n_829), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_940), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_940), .Y(n_1031) );
BUFx3_ASAP7_75t_L g1032 ( .A(n_920), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_855), .B(n_941), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_940), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_942), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_941), .B(n_888), .Y(n_1036) );
NAND2x1p5_ASAP7_75t_L g1037 ( .A(n_868), .B(n_885), .Y(n_1037) );
BUFx2_ASAP7_75t_L g1038 ( .A(n_925), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_942), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_921), .B(n_914), .Y(n_1040) );
INVx8_ASAP7_75t_L g1041 ( .A(n_868), .Y(n_1041) );
OAI21xp5_ASAP7_75t_L g1042 ( .A1(n_824), .A2(n_876), .B(n_878), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_925), .B(n_930), .Y(n_1043) );
AO31x2_ASAP7_75t_L g1044 ( .A1(n_856), .A2(n_926), .A3(n_851), .B(n_849), .Y(n_1044) );
INVx2_ASAP7_75t_SL g1045 ( .A(n_930), .Y(n_1045) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_828), .B(n_835), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_942), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_928), .A2(n_934), .B1(n_930), .B2(n_850), .Y(n_1048) );
INVxp33_ASAP7_75t_L g1049 ( .A(n_831), .Y(n_1049) );
OAI21x1_ASAP7_75t_SL g1050 ( .A1(n_935), .A2(n_928), .B(n_879), .Y(n_1050) );
AND2x4_ASAP7_75t_L g1051 ( .A(n_836), .B(n_919), .Y(n_1051) );
OAI21x1_ASAP7_75t_SL g1052 ( .A1(n_877), .A2(n_903), .B(n_883), .Y(n_1052) );
OAI21xp5_ASAP7_75t_L g1053 ( .A1(n_917), .A2(n_932), .B(n_922), .Y(n_1053) );
AND2x4_ASAP7_75t_L g1054 ( .A(n_945), .B(n_860), .Y(n_1054) );
OA21x2_ASAP7_75t_L g1055 ( .A1(n_904), .A2(n_907), .B(n_945), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_854), .Y(n_1056) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_927), .Y(n_1057) );
AOI21x1_ASAP7_75t_L g1058 ( .A1(n_927), .A2(n_873), .B(n_929), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_873), .B(n_927), .Y(n_1059) );
AO31x2_ASAP7_75t_L g1060 ( .A1(n_873), .A2(n_827), .A3(n_856), .B(n_898), .Y(n_1060) );
NAND3xp33_ASAP7_75t_L g1061 ( .A(n_929), .B(n_926), .C(n_827), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_929), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_943), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1064 ( .A1(n_817), .A2(n_720), .B(n_704), .Y(n_1064) );
AO21x2_ASAP7_75t_L g1065 ( .A1(n_827), .A2(n_819), .B(n_833), .Y(n_1065) );
OR2x6_ASAP7_75t_L g1066 ( .A(n_887), .B(n_678), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_892), .Y(n_1067) );
AO21x2_ASAP7_75t_L g1068 ( .A1(n_827), .A2(n_819), .B(n_833), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_821), .B(n_637), .Y(n_1069) );
OAI21x1_ASAP7_75t_SL g1070 ( .A1(n_871), .A2(n_712), .B(n_898), .Y(n_1070) );
OAI21xp5_ASAP7_75t_L g1071 ( .A1(n_827), .A2(n_741), .B(n_704), .Y(n_1071) );
NOR2x1_ASAP7_75t_SL g1072 ( .A(n_892), .B(n_739), .Y(n_1072) );
AO21x2_ASAP7_75t_L g1073 ( .A1(n_827), .A2(n_819), .B(n_833), .Y(n_1073) );
OA21x2_ASAP7_75t_L g1074 ( .A1(n_819), .A2(n_834), .B(n_827), .Y(n_1074) );
AOI21xp5_ASAP7_75t_L g1075 ( .A1(n_817), .A2(n_720), .B(n_704), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1063), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_960), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_951), .B(n_1067), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1069), .B(n_963), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1066), .B(n_985), .Y(n_1080) );
AO21x2_ASAP7_75t_L g1081 ( .A1(n_1042), .A2(n_1027), .B(n_1052), .Y(n_1081) );
INVx5_ASAP7_75t_SL g1082 ( .A(n_1066), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_969), .A2(n_971), .B1(n_990), .B2(n_1004), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_985), .B(n_955), .Y(n_1084) );
AO21x2_ASAP7_75t_L g1085 ( .A1(n_1027), .A2(n_1059), .B(n_1050), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_966), .Y(n_1086) );
AND2x4_ASAP7_75t_L g1087 ( .A(n_1072), .B(n_1009), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_987), .B(n_974), .Y(n_1088) );
OR2x6_ASAP7_75t_L g1089 ( .A(n_1009), .B(n_981), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_962), .Y(n_1090) );
AO21x2_ASAP7_75t_L g1091 ( .A1(n_1059), .A2(n_1061), .B(n_1031), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_958), .B(n_999), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_998), .B(n_967), .Y(n_1093) );
OAI21xp5_ASAP7_75t_L g1094 ( .A1(n_1025), .A2(n_959), .B(n_1028), .Y(n_1094) );
INVx5_ASAP7_75t_L g1095 ( .A(n_1041), .Y(n_1095) );
AO21x2_ASAP7_75t_L g1096 ( .A1(n_1061), .A2(n_1034), .B(n_1030), .Y(n_1096) );
OAI21xp5_ASAP7_75t_L g1097 ( .A1(n_980), .A2(n_1026), .B(n_964), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1014), .B(n_1020), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1021), .B(n_1033), .Y(n_1099) );
AO21x2_ASAP7_75t_L g1100 ( .A1(n_1035), .A2(n_1047), .B(n_1039), .Y(n_1100) );
OR2x6_ASAP7_75t_L g1101 ( .A(n_1003), .B(n_1041), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1005), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1006), .B(n_1008), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_1043), .Y(n_1104) );
AO21x2_ASAP7_75t_L g1105 ( .A1(n_1071), .A2(n_1022), .B(n_1058), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_952), .Y(n_1106) );
AO21x2_ASAP7_75t_L g1107 ( .A1(n_1071), .A2(n_1075), .B(n_1064), .Y(n_1107) );
NOR2xp33_ASAP7_75t_L g1108 ( .A(n_1046), .B(n_997), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1017), .B(n_993), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_991), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_991), .Y(n_1111) );
OAI21xp5_ASAP7_75t_L g1112 ( .A1(n_980), .A2(n_978), .B(n_979), .Y(n_1112) );
INVxp67_ASAP7_75t_L g1113 ( .A(n_992), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1013), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_970), .B(n_989), .Y(n_1115) );
OR2x6_ASAP7_75t_L g1116 ( .A(n_1024), .B(n_956), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1036), .B(n_1049), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_968), .Y(n_1118) );
HB1xp67_ASAP7_75t_L g1119 ( .A(n_1057), .Y(n_1119) );
BUFx6f_ASAP7_75t_L g1120 ( .A(n_1037), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1002), .B(n_976), .Y(n_1121) );
BUFx3_ASAP7_75t_L g1122 ( .A(n_961), .Y(n_1122) );
OA21x2_ASAP7_75t_L g1123 ( .A1(n_1056), .A2(n_1029), .B(n_1019), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1023), .B(n_1032), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_965), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1019), .B(n_1062), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1054), .Y(n_1127) );
OA21x2_ASAP7_75t_L g1128 ( .A1(n_1054), .A2(n_973), .B(n_1053), .Y(n_1128) );
AO21x2_ASAP7_75t_L g1129 ( .A1(n_1048), .A2(n_1053), .B(n_1070), .Y(n_1129) );
NOR2xp33_ASAP7_75t_L g1130 ( .A(n_996), .B(n_1040), .Y(n_1130) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1011), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_950), .B(n_1038), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1001), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1001), .Y(n_1134) );
OR2x2_ASAP7_75t_L g1135 ( .A(n_982), .B(n_1024), .Y(n_1135) );
INVx2_ASAP7_75t_L g1136 ( .A(n_995), .Y(n_1136) );
AO21x2_ASAP7_75t_L g1137 ( .A1(n_1048), .A2(n_983), .B(n_1065), .Y(n_1137) );
NAND2xp5_ASAP7_75t_SL g1138 ( .A(n_1051), .B(n_1015), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_988), .B(n_1024), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_1045), .B(n_1051), .Y(n_1140) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_1018), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_972), .B(n_1044), .Y(n_1142) );
OAI22xp33_ASAP7_75t_L g1143 ( .A1(n_1015), .A2(n_977), .B1(n_975), .B2(n_1055), .Y(n_1143) );
INVx6_ASAP7_75t_L g1144 ( .A(n_953), .Y(n_1144) );
BUFx3_ASAP7_75t_L g1145 ( .A(n_994), .Y(n_1145) );
INVx4_ASAP7_75t_L g1146 ( .A(n_1010), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1044), .B(n_1000), .Y(n_1147) );
AO21x2_ASAP7_75t_L g1148 ( .A1(n_1065), .A2(n_1068), .B(n_1073), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1060), .B(n_1012), .Y(n_1149) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1074), .Y(n_1150) );
INVx2_ASAP7_75t_SL g1151 ( .A(n_1060), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1073), .B(n_984), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_984), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_1016), .A2(n_1007), .B1(n_957), .B2(n_977), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1016), .B(n_957), .Y(n_1155) );
CKINVDCx5p33_ASAP7_75t_R g1156 ( .A(n_953), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1069), .B(n_986), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_954), .B(n_837), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1099), .B(n_1126), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1076), .Y(n_1160) );
BUFx2_ASAP7_75t_L g1161 ( .A(n_1089), .Y(n_1161) );
AND2x4_ASAP7_75t_L g1162 ( .A(n_1140), .B(n_1103), .Y(n_1162) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_1104), .Y(n_1163) );
HB1xp67_ASAP7_75t_L g1164 ( .A(n_1104), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_1117), .B(n_1119), .Y(n_1165) );
BUFx2_ASAP7_75t_L g1166 ( .A(n_1089), .Y(n_1166) );
NOR2xp67_ASAP7_75t_SL g1167 ( .A(n_1095), .B(n_1145), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1098), .B(n_1088), .Y(n_1168) );
INVx1_ASAP7_75t_SL g1169 ( .A(n_1122), .Y(n_1169) );
BUFx3_ASAP7_75t_L g1170 ( .A(n_1095), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1078), .B(n_1158), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_1097), .A2(n_1106), .B1(n_1111), .B2(n_1110), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_1119), .B(n_1157), .Y(n_1173) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_1108), .A2(n_1130), .B1(n_1109), .B2(n_1092), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1158), .B(n_1092), .Y(n_1175) );
OR2x6_ASAP7_75t_SL g1176 ( .A(n_1156), .B(n_1135), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1102), .B(n_1079), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1077), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1086), .Y(n_1179) );
OAI211xp5_ASAP7_75t_SL g1180 ( .A1(n_1113), .A2(n_1114), .B(n_1108), .C(n_1115), .Y(n_1180) );
INVx3_ASAP7_75t_L g1181 ( .A(n_1087), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1127), .B(n_1091), .Y(n_1182) );
HB1xp67_ASAP7_75t_L g1183 ( .A(n_1141), .Y(n_1183) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1100), .Y(n_1184) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1100), .Y(n_1185) );
AND2x4_ASAP7_75t_L g1186 ( .A(n_1087), .B(n_1116), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1123), .B(n_1096), .Y(n_1187) );
BUFx3_ASAP7_75t_L g1188 ( .A(n_1095), .Y(n_1188) );
INVx1_ASAP7_75t_SL g1189 ( .A(n_1122), .Y(n_1189) );
AND2x4_ASAP7_75t_L g1190 ( .A(n_1118), .B(n_1138), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1090), .B(n_1112), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1085), .B(n_1105), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1105), .B(n_1151), .Y(n_1193) );
NOR2xp33_ASAP7_75t_L g1194 ( .A(n_1139), .B(n_1130), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1150), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1093), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1081), .B(n_1094), .Y(n_1197) );
INVx4_ASAP7_75t_L g1198 ( .A(n_1101), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1084), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_1083), .A2(n_1082), .B1(n_1125), .B2(n_1080), .Y(n_1200) );
AND2x4_ASAP7_75t_L g1201 ( .A(n_1138), .B(n_1129), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1083), .B(n_1132), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1132), .B(n_1124), .Y(n_1203) );
OR2x2_ASAP7_75t_L g1204 ( .A(n_1133), .B(n_1134), .Y(n_1204) );
BUFx2_ASAP7_75t_L g1205 ( .A(n_1101), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1160), .Y(n_1206) );
NAND5xp2_ASAP7_75t_L g1207 ( .A(n_1200), .B(n_1121), .C(n_1154), .D(n_1147), .E(n_1155), .Y(n_1207) );
HB1xp67_ASAP7_75t_L g1208 ( .A(n_1183), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1159), .B(n_1137), .Y(n_1209) );
AND2x4_ASAP7_75t_L g1210 ( .A(n_1190), .B(n_1137), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1165), .B(n_1153), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1178), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1175), .B(n_1142), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1168), .B(n_1152), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1197), .B(n_1148), .Y(n_1215) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1195), .Y(n_1216) );
NOR2xp33_ASAP7_75t_L g1217 ( .A(n_1169), .B(n_1189), .Y(n_1217) );
AND2x4_ASAP7_75t_SL g1218 ( .A(n_1198), .B(n_1101), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1179), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1171), .B(n_1107), .Y(n_1220) );
NOR2xp33_ASAP7_75t_L g1221 ( .A(n_1194), .B(n_1146), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1162), .B(n_1128), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1162), .B(n_1155), .Y(n_1223) );
BUFx3_ASAP7_75t_L g1224 ( .A(n_1170), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1196), .B(n_1120), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1173), .B(n_1149), .Y(n_1226) );
INVx4_ASAP7_75t_L g1227 ( .A(n_1188), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1182), .B(n_1131), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1177), .Y(n_1229) );
NOR2xp33_ASAP7_75t_L g1230 ( .A(n_1194), .B(n_1146), .Y(n_1230) );
HB1xp67_ASAP7_75t_L g1231 ( .A(n_1163), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1192), .B(n_1136), .Y(n_1232) );
HB1xp67_ASAP7_75t_L g1233 ( .A(n_1164), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1216), .Y(n_1234) );
AND2x4_ASAP7_75t_L g1235 ( .A(n_1210), .B(n_1193), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1220), .B(n_1201), .Y(n_1236) );
OAI21xp33_ASAP7_75t_L g1237 ( .A1(n_1207), .A2(n_1172), .B(n_1174), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1206), .Y(n_1238) );
INVxp67_ASAP7_75t_SL g1239 ( .A(n_1208), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1240 ( .A(n_1231), .Y(n_1240) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_1210), .B(n_1187), .Y(n_1241) );
AND2x4_ASAP7_75t_L g1242 ( .A(n_1210), .B(n_1187), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1214), .B(n_1184), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1212), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1214), .B(n_1185), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1213), .B(n_1185), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1219), .Y(n_1247) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1228), .Y(n_1248) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1232), .Y(n_1249) );
INVx2_ASAP7_75t_L g1250 ( .A(n_1232), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1215), .B(n_1191), .Y(n_1251) );
AOI32xp33_ASAP7_75t_SL g1252 ( .A1(n_1239), .A2(n_1221), .A3(n_1230), .B1(n_1217), .B2(n_1229), .Y(n_1252) );
AOI211xp5_ASAP7_75t_L g1253 ( .A1(n_1237), .A2(n_1167), .B(n_1180), .C(n_1209), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1251), .B(n_1233), .Y(n_1254) );
NOR2xp33_ASAP7_75t_L g1255 ( .A(n_1240), .B(n_1176), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1238), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1238), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_1237), .A2(n_1223), .B1(n_1202), .B2(n_1226), .Y(n_1258) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1234), .Y(n_1259) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1259), .Y(n_1260) );
AOI22xp5_ASAP7_75t_L g1261 ( .A1(n_1258), .A2(n_1241), .B1(n_1242), .B2(n_1235), .Y(n_1261) );
AOI22xp5_ASAP7_75t_L g1262 ( .A1(n_1253), .A2(n_1241), .B1(n_1242), .B2(n_1235), .Y(n_1262) );
NAND2xp5_ASAP7_75t_SL g1263 ( .A(n_1255), .B(n_1227), .Y(n_1263) );
INVx1_ASAP7_75t_SL g1264 ( .A(n_1254), .Y(n_1264) );
A2O1A1Ixp33_ASAP7_75t_L g1265 ( .A1(n_1252), .A2(n_1218), .B(n_1205), .C(n_1186), .Y(n_1265) );
NAND3x2_ASAP7_75t_L g1266 ( .A(n_1252), .B(n_1166), .C(n_1161), .Y(n_1266) );
AOI22xp5_ASAP7_75t_L g1267 ( .A1(n_1261), .A2(n_1262), .B1(n_1264), .B2(n_1263), .Y(n_1267) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_1266), .A2(n_1223), .B1(n_1222), .B2(n_1236), .Y(n_1268) );
NAND3xp33_ASAP7_75t_L g1269 ( .A(n_1265), .B(n_1256), .C(n_1257), .Y(n_1269) );
NAND4xp75_ASAP7_75t_L g1270 ( .A(n_1260), .B(n_1243), .C(n_1245), .D(n_1246), .Y(n_1270) );
NAND3xp33_ASAP7_75t_L g1271 ( .A(n_1268), .B(n_1269), .C(n_1267), .Y(n_1271) );
NOR3xp33_ASAP7_75t_SL g1272 ( .A(n_1271), .B(n_1144), .C(n_1270), .Y(n_1272) );
AND2x4_ASAP7_75t_L g1273 ( .A(n_1272), .B(n_1199), .Y(n_1273) );
XNOR2x1_ASAP7_75t_L g1274 ( .A(n_1273), .B(n_1224), .Y(n_1274) );
INVx2_ASAP7_75t_L g1275 ( .A(n_1274), .Y(n_1275) );
AOI21xp5_ASAP7_75t_L g1276 ( .A1(n_1275), .A2(n_1244), .B(n_1247), .Y(n_1276) );
OAI21x1_ASAP7_75t_SL g1277 ( .A1(n_1276), .A2(n_1203), .B(n_1225), .Y(n_1277) );
AOI21xp33_ASAP7_75t_L g1278 ( .A1(n_1277), .A2(n_1204), .B(n_1211), .Y(n_1278) );
NOR3xp33_ASAP7_75t_L g1279 ( .A(n_1278), .B(n_1181), .C(n_1143), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_1279), .A2(n_1248), .B1(n_1250), .B2(n_1249), .Y(n_1280) );
endmodule