module real_aes_10713_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1346;
wire n_1383;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_269;
wire n_430;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1352;
wire n_729;
wire n_394;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_1369;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_0), .A2(n_23), .B1(n_531), .B2(n_541), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_0), .A2(n_231), .B1(n_367), .B2(n_544), .Y(n_611) );
INVx1_ASAP7_75t_L g813 ( .A(n_1), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_1), .A2(n_135), .B1(n_721), .B2(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g1259 ( .A(n_2), .Y(n_1259) );
OAI221xp5_ASAP7_75t_L g1311 ( .A1(n_2), .A2(n_76), .B1(n_1312), .B2(n_1317), .C(n_1321), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g1271 ( .A1(n_3), .A2(n_243), .B1(n_796), .B2(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1334 ( .A(n_3), .Y(n_1334) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_4), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_4), .A2(n_29), .B1(n_392), .B2(n_393), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_5), .A2(n_111), .B1(n_392), .B2(n_733), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_5), .A2(n_111), .B1(n_526), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_6), .A2(n_13), .B1(n_516), .B2(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g843 ( .A(n_6), .Y(n_843) );
INVx1_ASAP7_75t_L g866 ( .A(n_7), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_8), .A2(n_10), .B1(n_1047), .B2(n_1064), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_9), .Y(n_262) );
INVx1_ASAP7_75t_L g399 ( .A(n_9), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_9), .B(n_186), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_9), .B(n_346), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_11), .A2(n_95), .B1(n_606), .B2(n_656), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_11), .A2(n_95), .B1(n_691), .B2(n_693), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g454 ( .A1(n_12), .A2(n_201), .B1(n_378), .B2(n_379), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_12), .A2(n_201), .B1(n_408), .B2(n_419), .Y(n_465) );
INVx1_ASAP7_75t_L g844 ( .A(n_13), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_14), .A2(n_43), .B1(n_740), .B2(n_742), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_14), .A2(n_43), .B1(n_745), .B2(n_747), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g1067 ( .A1(n_15), .A2(n_214), .B1(n_1053), .B2(n_1056), .Y(n_1067) );
INVx1_ASAP7_75t_L g708 ( .A(n_16), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_17), .A2(n_171), .B1(n_378), .B2(n_379), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_17), .A2(n_171), .B1(n_406), .B2(n_408), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_18), .A2(n_240), .B1(n_408), .B2(n_419), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_18), .A2(n_240), .B1(n_544), .B2(n_554), .Y(n_1014) );
AO22x2_ASAP7_75t_L g852 ( .A1(n_19), .A2(n_853), .B1(n_913), .B2(n_914), .Y(n_852) );
INVx1_ASAP7_75t_L g913 ( .A(n_19), .Y(n_913) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_20), .Y(n_537) );
CKINVDCx14_ASAP7_75t_R g1072 ( .A(n_21), .Y(n_1072) );
INVx1_ASAP7_75t_L g295 ( .A(n_22), .Y(n_295) );
INVx1_ASAP7_75t_L g596 ( .A(n_23), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_24), .Y(n_807) );
AOI221xp5_ASAP7_75t_L g1268 ( .A1(n_25), .A2(n_41), .B1(n_526), .B2(n_747), .C(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1336 ( .A(n_25), .Y(n_1336) );
AOI22xp33_ASAP7_75t_L g1374 ( .A1(n_26), .A2(n_127), .B1(n_442), .B2(n_691), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_26), .A2(n_127), .B1(n_606), .B2(n_656), .Y(n_1385) );
AOI22xp33_ASAP7_75t_SL g885 ( .A1(n_27), .A2(n_239), .B1(n_886), .B2(n_887), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_27), .A2(n_239), .B1(n_747), .B2(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g811 ( .A(n_28), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_28), .A2(n_246), .B1(n_392), .B2(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g317 ( .A(n_29), .Y(n_317) );
INVx1_ASAP7_75t_L g429 ( .A(n_30), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_30), .A2(n_123), .B1(n_338), .B2(n_456), .Y(n_460) );
XNOR2xp5_ASAP7_75t_L g559 ( .A(n_31), .B(n_560), .Y(n_559) );
INVxp67_ASAP7_75t_SL g1368 ( .A(n_32), .Y(n_1368) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_32), .A2(n_196), .B1(n_830), .B2(n_1393), .Y(n_1392) );
INVxp33_ASAP7_75t_L g928 ( .A(n_33), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_33), .A2(n_212), .B1(n_960), .B2(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g279 ( .A(n_34), .Y(n_279) );
INVx2_ASAP7_75t_L g287 ( .A(n_35), .Y(n_287) );
OR2x2_ASAP7_75t_L g1266 ( .A(n_35), .B(n_1256), .Y(n_1266) );
INVx1_ASAP7_75t_L g638 ( .A(n_36), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_36), .A2(n_114), .B1(n_660), .B2(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g629 ( .A(n_37), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_37), .A2(n_101), .B1(n_674), .B2(n_675), .Y(n_673) );
BUFx2_ASAP7_75t_L g333 ( .A(n_38), .Y(n_333) );
BUFx2_ASAP7_75t_L g374 ( .A(n_38), .Y(n_374) );
INVx1_ASAP7_75t_L g672 ( .A(n_38), .Y(n_672) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_38), .B(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g650 ( .A(n_39), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_39), .A2(n_51), .B1(n_656), .B2(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g711 ( .A(n_40), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_40), .A2(n_99), .B1(n_381), .B2(n_721), .Y(n_735) );
INVx1_ASAP7_75t_L g1327 ( .A(n_41), .Y(n_1327) );
CKINVDCx5p33_ASAP7_75t_R g1276 ( .A(n_42), .Y(n_1276) );
INVx1_ASAP7_75t_L g717 ( .A(n_44), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_44), .A2(n_141), .B1(n_348), .B2(n_351), .Y(n_723) );
INVxp33_ASAP7_75t_L g774 ( .A(n_45), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_45), .A2(n_147), .B1(n_677), .B2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_46), .A2(n_56), .B1(n_392), .B2(n_738), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_46), .A2(n_56), .B1(n_749), .B2(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g609 ( .A(n_47), .Y(n_609) );
AO22x2_ASAP7_75t_L g618 ( .A1(n_48), .A2(n_619), .B1(n_620), .B2(n_696), .Y(n_618) );
INVx1_ASAP7_75t_L g696 ( .A(n_48), .Y(n_696) );
INVxp67_ASAP7_75t_SL g1353 ( .A(n_49), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_49), .A2(n_120), .B1(n_351), .B2(n_646), .Y(n_1366) );
INVx1_ASAP7_75t_L g937 ( .A(n_50), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_50), .A2(n_136), .B1(n_949), .B2(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g640 ( .A(n_51), .Y(n_640) );
INVx1_ASAP7_75t_L g433 ( .A(n_52), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_52), .A2(n_225), .B1(n_379), .B2(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g283 ( .A(n_53), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_53), .A2(n_185), .B1(n_338), .B2(n_381), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_54), .A2(n_237), .B1(n_408), .B2(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_54), .A2(n_172), .B1(n_367), .B2(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g859 ( .A(n_55), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_57), .A2(n_137), .B1(n_721), .B2(n_949), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_57), .A2(n_137), .B1(n_865), .B2(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g628 ( .A(n_58), .Y(n_628) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_58), .A2(n_72), .B1(n_680), .B2(n_683), .Y(n_679) );
INVxp33_ASAP7_75t_L g768 ( .A(n_59), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_59), .A2(n_92), .B1(n_747), .B2(n_796), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_60), .A2(n_86), .B1(n_529), .B2(n_531), .Y(n_978) );
INVx1_ASAP7_75t_L g994 ( .A(n_60), .Y(n_994) );
INVx1_ASAP7_75t_L g499 ( .A(n_61), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_61), .A2(n_172), .B1(n_529), .B2(n_531), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g1068 ( .A1(n_62), .A2(n_90), .B1(n_1047), .B2(n_1064), .Y(n_1068) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_63), .A2(n_227), .B1(n_540), .B2(n_541), .Y(n_984) );
AOI221xp5_ASAP7_75t_L g992 ( .A1(n_63), .A2(n_227), .B1(n_944), .B2(n_953), .C(n_993), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_64), .A2(n_234), .B1(n_303), .B2(n_463), .Y(n_832) );
INVx1_ASAP7_75t_L g838 ( .A(n_64), .Y(n_838) );
AOI22xp5_ASAP7_75t_SL g1058 ( .A1(n_65), .A2(n_82), .B1(n_1041), .B2(n_1047), .Y(n_1058) );
INVx1_ASAP7_75t_L g608 ( .A(n_66), .Y(n_608) );
INVx1_ASAP7_75t_L g575 ( .A(n_67), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_68), .A2(n_220), .B1(n_944), .B2(n_946), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_68), .A2(n_220), .B1(n_963), .B2(n_964), .Y(n_962) );
CKINVDCx16_ASAP7_75t_R g1045 ( .A(n_69), .Y(n_1045) );
INVx1_ASAP7_75t_L g764 ( .A(n_70), .Y(n_764) );
INVxp67_ASAP7_75t_SL g727 ( .A(n_71), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_71), .A2(n_140), .B1(n_660), .B2(n_754), .Y(n_753) );
OAI222xp33_ASAP7_75t_L g623 ( .A1(n_72), .A2(n_151), .B1(n_233), .B2(n_308), .C1(n_313), .C2(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g926 ( .A(n_73), .Y(n_926) );
INVx1_ASAP7_75t_L g451 ( .A(n_74), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_74), .A2(n_85), .B1(n_419), .B2(n_420), .Y(n_468) );
INVx1_ASAP7_75t_L g493 ( .A(n_75), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_75), .A2(n_164), .B1(n_540), .B2(n_541), .Y(n_539) );
INVx1_ASAP7_75t_L g1262 ( .A(n_76), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_77), .A2(n_145), .B1(n_338), .B2(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_77), .A2(n_145), .B1(n_303), .B2(n_463), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_78), .A2(n_105), .B1(n_313), .B2(n_438), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_78), .A2(n_105), .B1(n_351), .B2(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g364 ( .A(n_79), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_79), .A2(n_98), .B1(n_419), .B2(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g580 ( .A(n_80), .Y(n_580) );
OAI211xp5_ASAP7_75t_SL g612 ( .A1(n_80), .A2(n_546), .B(n_548), .C(n_613), .Y(n_612) );
AO22x2_ASAP7_75t_L g756 ( .A1(n_81), .A2(n_757), .B1(n_798), .B2(n_799), .Y(n_756) );
INVx1_ASAP7_75t_L g798 ( .A(n_81), .Y(n_798) );
INVxp33_ASAP7_75t_SL g706 ( .A(n_83), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_83), .A2(n_161), .B1(n_392), .B2(n_733), .Y(n_732) );
INVxp67_ASAP7_75t_SL g860 ( .A(n_84), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_84), .A2(n_191), .B1(n_674), .B2(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g449 ( .A(n_85), .Y(n_449) );
INVx1_ASAP7_75t_L g1013 ( .A(n_86), .Y(n_1013) );
INVx1_ASAP7_75t_L g331 ( .A(n_87), .Y(n_331) );
INVx1_ASAP7_75t_L g1256 ( .A(n_87), .Y(n_1256) );
INVxp33_ASAP7_75t_SL g873 ( .A(n_88), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_88), .A2(n_183), .B1(n_667), .B2(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g862 ( .A(n_89), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_89), .A2(n_176), .B1(n_887), .B2(n_895), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_91), .A2(n_190), .B1(n_674), .B2(n_883), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_91), .A2(n_190), .B1(n_901), .B2(n_903), .Y(n_900) );
INVx1_ASAP7_75t_L g763 ( .A(n_92), .Y(n_763) );
INVx1_ASAP7_75t_L g524 ( .A(n_93), .Y(n_524) );
OAI211xp5_ASAP7_75t_SL g545 ( .A1(n_93), .A2(n_546), .B(n_548), .C(n_549), .Y(n_545) );
NAND2xp33_ASAP7_75t_SL g1250 ( .A(n_94), .B(n_865), .Y(n_1250) );
INVx1_ASAP7_75t_L g1304 ( .A(n_94), .Y(n_1304) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_96), .A2(n_180), .B1(n_308), .B2(n_313), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_96), .A2(n_180), .B1(n_348), .B2(n_351), .Y(n_347) );
INVx1_ASAP7_75t_L g569 ( .A(n_97), .Y(n_569) );
INVxp67_ASAP7_75t_L g372 ( .A(n_98), .Y(n_372) );
INVxp33_ASAP7_75t_SL g705 ( .A(n_99), .Y(n_705) );
INVx1_ASAP7_75t_L g989 ( .A(n_100), .Y(n_989) );
INVx1_ASAP7_75t_L g632 ( .A(n_101), .Y(n_632) );
INVxp67_ASAP7_75t_SL g1357 ( .A(n_102), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_102), .A2(n_232), .B1(n_1380), .B2(n_1381), .Y(n_1379) );
INVx1_ASAP7_75t_L g600 ( .A(n_103), .Y(n_600) );
INVx1_ASAP7_75t_L g816 ( .A(n_104), .Y(n_816) );
OAI22xp33_ASAP7_75t_L g840 ( .A1(n_104), .A2(n_175), .B1(n_646), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_106), .A2(n_130), .B1(n_661), .B2(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_106), .A2(n_130), .B1(n_685), .B2(n_687), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_107), .A2(n_221), .B1(n_1053), .B2(n_1104), .Y(n_1103) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_108), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_108), .A2(n_179), .B1(n_408), .B2(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g1135 ( .A(n_109), .Y(n_1135) );
AOI222xp33_ASAP7_75t_L g1239 ( .A1(n_109), .A2(n_1240), .B1(n_1344), .B2(n_1346), .C1(n_1397), .C2(n_1401), .Y(n_1239) );
CKINVDCx5p33_ASAP7_75t_R g1283 ( .A(n_110), .Y(n_1283) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_112), .A2(n_217), .B1(n_378), .B2(n_379), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_112), .A2(n_217), .B1(n_750), .B2(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g579 ( .A(n_113), .Y(n_579) );
OAI22xp33_ASAP7_75t_SL g614 ( .A1(n_113), .A2(n_142), .B1(n_263), .B2(n_554), .Y(n_614) );
INVx1_ASAP7_75t_L g637 ( .A(n_114), .Y(n_637) );
INVx1_ASAP7_75t_L g254 ( .A(n_115), .Y(n_254) );
INVx1_ASAP7_75t_L g448 ( .A(n_116), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_116), .A2(n_195), .B1(n_416), .B2(n_463), .Y(n_467) );
INVx1_ASAP7_75t_L g1287 ( .A(n_117), .Y(n_1287) );
AOI221xp5_ASAP7_75t_L g986 ( .A1(n_118), .A2(n_197), .B1(n_674), .B2(n_987), .C(n_988), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_118), .A2(n_197), .B1(n_419), .B2(n_420), .Y(n_1004) );
INVx1_ASAP7_75t_L g983 ( .A(n_119), .Y(n_983) );
INVxp67_ASAP7_75t_SL g1354 ( .A(n_120), .Y(n_1354) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_121), .A2(n_206), .B1(n_1053), .B2(n_1056), .Y(n_1052) );
AOI22xp33_ASAP7_75t_SL g1247 ( .A1(n_122), .A2(n_205), .B1(n_419), .B2(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1309 ( .A(n_122), .Y(n_1309) );
INVx1_ASAP7_75t_L g436 ( .A(n_123), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g1375 ( .A1(n_124), .A2(n_156), .B1(n_685), .B2(n_1376), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_124), .A2(n_156), .B1(n_660), .B2(n_792), .Y(n_1384) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_125), .A2(n_126), .B1(n_1041), .B2(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g917 ( .A(n_128), .Y(n_917) );
CKINVDCx14_ASAP7_75t_R g975 ( .A(n_129), .Y(n_975) );
XOR2xp5_ASAP7_75t_L g470 ( .A(n_131), .B(n_471), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g1062 ( .A1(n_131), .A2(n_153), .B1(n_1053), .B2(n_1056), .Y(n_1062) );
INVx1_ASAP7_75t_L g982 ( .A(n_132), .Y(n_982) );
CKINVDCx5p33_ASAP7_75t_R g1267 ( .A(n_133), .Y(n_1267) );
INVx1_ASAP7_75t_L g769 ( .A(n_134), .Y(n_769) );
INVx1_ASAP7_75t_L g810 ( .A(n_135), .Y(n_810) );
INVxp33_ASAP7_75t_L g932 ( .A(n_136), .Y(n_932) );
INVxp33_ASAP7_75t_L g761 ( .A(n_138), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_138), .A2(n_146), .B1(n_526), .B2(n_750), .Y(n_797) );
INVx1_ASAP7_75t_L g572 ( .A(n_139), .Y(n_572) );
INVxp33_ASAP7_75t_L g725 ( .A(n_140), .Y(n_725) );
INVx1_ASAP7_75t_L g714 ( .A(n_141), .Y(n_714) );
INVx1_ASAP7_75t_L g584 ( .A(n_142), .Y(n_584) );
INVx1_ASAP7_75t_L g766 ( .A(n_143), .Y(n_766) );
INVxp67_ASAP7_75t_SL g933 ( .A(n_144), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_144), .A2(n_192), .B1(n_952), .B2(n_953), .Y(n_951) );
INVxp33_ASAP7_75t_L g760 ( .A(n_146), .Y(n_760) );
INVxp33_ASAP7_75t_L g776 ( .A(n_147), .Y(n_776) );
INVx1_ASAP7_75t_L g595 ( .A(n_148), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_148), .A2(n_169), .B1(n_529), .B2(n_540), .Y(n_602) );
INVx1_ASAP7_75t_L g482 ( .A(n_149), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_150), .A2(n_210), .B1(n_381), .B2(n_721), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_150), .A2(n_210), .B1(n_303), .B2(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g644 ( .A(n_151), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_152), .A2(n_223), .B1(n_787), .B2(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_152), .A2(n_223), .B1(n_303), .B2(n_463), .Y(n_828) );
CKINVDCx16_ASAP7_75t_R g1048 ( .A(n_154), .Y(n_1048) );
AO221x2_ASAP7_75t_L g1070 ( .A1(n_155), .A2(n_229), .B1(n_1047), .B2(n_1064), .C(n_1071), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_157), .A2(n_1347), .B1(n_1395), .B2(n_1396), .Y(n_1346) );
CKINVDCx5p33_ASAP7_75t_R g1396 ( .A(n_157), .Y(n_1396) );
INVx1_ASAP7_75t_L g921 ( .A(n_158), .Y(n_921) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_159), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_159), .B(n_254), .Y(n_1021) );
AND3x2_ASAP7_75t_L g1044 ( .A(n_159), .B(n_254), .C(n_1024), .Y(n_1044) );
AOI22xp5_ASAP7_75t_SL g1079 ( .A1(n_160), .A2(n_170), .B1(n_1041), .B2(n_1047), .Y(n_1079) );
INVxp33_ASAP7_75t_SL g709 ( .A(n_161), .Y(n_709) );
INVxp33_ASAP7_75t_SL g729 ( .A(n_162), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_162), .A2(n_211), .B1(n_745), .B2(n_747), .Y(n_752) );
INVxp33_ASAP7_75t_L g777 ( .A(n_163), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_163), .A2(n_168), .B1(n_721), .B2(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g496 ( .A(n_164), .Y(n_496) );
INVxp33_ASAP7_75t_SL g1359 ( .A(n_165), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_165), .A2(n_222), .B1(n_691), .B2(n_839), .Y(n_1378) );
INVx2_ASAP7_75t_L g267 ( .A(n_166), .Y(n_267) );
AOI22xp5_ASAP7_75t_SL g1078 ( .A1(n_167), .A2(n_226), .B1(n_1053), .B2(n_1056), .Y(n_1078) );
INVx1_ASAP7_75t_L g772 ( .A(n_168), .Y(n_772) );
INVx1_ASAP7_75t_L g598 ( .A(n_169), .Y(n_598) );
INVx1_ASAP7_75t_L g1024 ( .A(n_173), .Y(n_1024) );
INVxp67_ASAP7_75t_SL g922 ( .A(n_174), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_174), .A2(n_207), .B1(n_420), .B2(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g815 ( .A(n_175), .Y(n_815) );
INVxp33_ASAP7_75t_SL g856 ( .A(n_176), .Y(n_856) );
AO221x2_ASAP7_75t_L g1132 ( .A1(n_177), .A2(n_248), .B1(n_1106), .B2(n_1133), .C(n_1134), .Y(n_1132) );
INVxp67_ASAP7_75t_SL g1365 ( .A(n_178), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_178), .A2(n_219), .B1(n_1387), .B2(n_1390), .Y(n_1386) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_179), .Y(n_484) );
INVx1_ASAP7_75t_L g478 ( .A(n_181), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_182), .Y(n_431) );
INVxp33_ASAP7_75t_SL g874 ( .A(n_183), .Y(n_874) );
INVx1_ASAP7_75t_L g1006 ( .A(n_184), .Y(n_1006) );
INVx1_ASAP7_75t_L g306 ( .A(n_185), .Y(n_306) );
INVx1_ASAP7_75t_L g269 ( .A(n_186), .Y(n_269) );
INVx2_ASAP7_75t_L g346 ( .A(n_186), .Y(n_346) );
INVx1_ASAP7_75t_L g336 ( .A(n_187), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_187), .A2(n_236), .B1(n_415), .B2(n_416), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_188), .A2(n_216), .B1(n_381), .B2(n_385), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_188), .A2(n_216), .B1(n_402), .B2(n_403), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g425 ( .A(n_189), .B(n_426), .Y(n_425) );
INVxp33_ASAP7_75t_SL g857 ( .A(n_191), .Y(n_857) );
INVxp67_ASAP7_75t_SL g935 ( .A(n_192), .Y(n_935) );
OAI211xp5_ASAP7_75t_L g979 ( .A1(n_193), .A2(n_538), .B(n_980), .C(n_981), .Y(n_979) );
INVx1_ASAP7_75t_L g997 ( .A(n_193), .Y(n_997) );
CKINVDCx14_ASAP7_75t_R g1136 ( .A(n_194), .Y(n_1136) );
INVx1_ASAP7_75t_L g441 ( .A(n_195), .Y(n_441) );
INVxp33_ASAP7_75t_SL g1369 ( .A(n_196), .Y(n_1369) );
XNOR2xp5_ASAP7_75t_L g803 ( .A(n_198), .B(n_804), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_199), .Y(n_924) );
INVx1_ASAP7_75t_L g990 ( .A(n_200), .Y(n_990) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_202), .Y(n_631) );
CKINVDCx16_ASAP7_75t_R g1038 ( .A(n_203), .Y(n_1038) );
INVx1_ASAP7_75t_L g521 ( .A(n_204), .Y(n_521) );
OAI22xp33_ASAP7_75t_SL g553 ( .A1(n_204), .A2(n_237), .B1(n_263), .B2(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g1299 ( .A(n_205), .Y(n_1299) );
INVxp67_ASAP7_75t_SL g929 ( .A(n_207), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g1279 ( .A(n_208), .Y(n_1279) );
INVx1_ASAP7_75t_L g1356 ( .A(n_209), .Y(n_1356) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_211), .Y(n_722) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_212), .Y(n_925) );
INVx1_ASAP7_75t_L g1025 ( .A(n_213), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_213), .B(n_1023), .Y(n_1037) );
XOR2x2_ASAP7_75t_L g701 ( .A(n_214), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g566 ( .A(n_215), .Y(n_566) );
INVx1_ASAP7_75t_L g869 ( .A(n_218), .Y(n_869) );
INVxp33_ASAP7_75t_SL g1363 ( .A(n_219), .Y(n_1363) );
INVx1_ASAP7_75t_L g1352 ( .A(n_222), .Y(n_1352) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_224), .Y(n_536) );
INVx1_ASAP7_75t_L g434 ( .A(n_225), .Y(n_434) );
INVx2_ASAP7_75t_L g266 ( .A(n_228), .Y(n_266) );
AOI21xp33_ASAP7_75t_L g1251 ( .A1(n_230), .A2(n_796), .B(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g1307 ( .A(n_230), .Y(n_1307) );
INVx1_ASAP7_75t_L g586 ( .A(n_231), .Y(n_586) );
INVxp67_ASAP7_75t_SL g1360 ( .A(n_232), .Y(n_1360) );
INVx1_ASAP7_75t_L g647 ( .A(n_233), .Y(n_647) );
INVx1_ASAP7_75t_L g846 ( .A(n_234), .Y(n_846) );
INVxp33_ASAP7_75t_SL g879 ( .A(n_235), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_235), .A2(n_247), .B1(n_814), .B2(n_908), .Y(n_907) );
INVxp33_ASAP7_75t_L g356 ( .A(n_236), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g1033 ( .A(n_238), .Y(n_1033) );
BUFx3_ASAP7_75t_L g292 ( .A(n_241), .Y(n_292) );
INVx1_ASAP7_75t_L g325 ( .A(n_241), .Y(n_325) );
BUFx3_ASAP7_75t_L g294 ( .A(n_242), .Y(n_294) );
INVx1_ASAP7_75t_L g320 ( .A(n_242), .Y(n_320) );
INVx1_ASAP7_75t_L g1329 ( .A(n_243), .Y(n_1329) );
INVx1_ASAP7_75t_L g1007 ( .A(n_244), .Y(n_1007) );
INVx1_ASAP7_75t_L g502 ( .A(n_245), .Y(n_502) );
INVx1_ASAP7_75t_L g808 ( .A(n_246), .Y(n_808) );
INVx1_ASAP7_75t_L g876 ( .A(n_247), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_1015), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_257), .Y(n_251) );
AND2x4_ASAP7_75t_L g1345 ( .A(n_252), .B(n_258), .Y(n_1345) );
NOR2xp33_ASAP7_75t_SL g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx1_ASAP7_75t_SL g1400 ( .A(n_253), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_253), .B(n_255), .Y(n_1402) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_255), .B(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_263), .Y(n_258) );
INVxp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g373 ( .A(n_260), .B(n_374), .Y(n_373) );
OR2x6_ASAP7_75t_L g558 ( .A(n_260), .B(n_374), .Y(n_558) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g389 ( .A(n_261), .B(n_269), .Y(n_389) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g475 ( .A(n_262), .B(n_359), .Y(n_475) );
INVx8_ASAP7_75t_L g355 ( .A(n_263), .Y(n_355) );
OR2x6_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
OR2x6_ASAP7_75t_L g367 ( .A(n_264), .B(n_358), .Y(n_367) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_264), .Y(n_477) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_264), .Y(n_498) );
INVx2_ASAP7_75t_SL g591 ( .A(n_264), .Y(n_591) );
INVx2_ASAP7_75t_SL g996 ( .A(n_264), .Y(n_996) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_264), .B(n_1291), .Y(n_1290) );
BUFx2_ASAP7_75t_L g1333 ( .A(n_264), .Y(n_1333) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g340 ( .A(n_266), .Y(n_340) );
INVx1_ASAP7_75t_L g353 ( .A(n_266), .Y(n_353) );
INVx2_ASAP7_75t_L g361 ( .A(n_266), .Y(n_361) );
AND2x4_ASAP7_75t_L g371 ( .A(n_266), .B(n_341), .Y(n_371) );
AND2x2_ASAP7_75t_L g384 ( .A(n_266), .B(n_267), .Y(n_384) );
INVx2_ASAP7_75t_L g341 ( .A(n_267), .Y(n_341) );
INVx1_ASAP7_75t_L g350 ( .A(n_267), .Y(n_350) );
INVx1_ASAP7_75t_L g363 ( .A(n_267), .Y(n_363) );
INVx1_ASAP7_75t_L g481 ( .A(n_267), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_267), .B(n_361), .Y(n_487) );
AND2x4_ASAP7_75t_L g349 ( .A(n_268), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g351 ( .A(n_269), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g841 ( .A(n_269), .B(n_352), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B1(n_697), .B2(n_698), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_617), .B2(n_618), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
XOR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_469), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B1(n_424), .B2(n_425), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
XNOR2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AOI211xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_329), .B(n_334), .C(n_375), .Y(n_280) );
NAND4xp25_ASAP7_75t_L g281 ( .A(n_282), .B(n_299), .C(n_316), .D(n_326), .Y(n_281) );
AOI22xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_284), .B1(n_295), .B2(n_296), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_284), .A2(n_318), .B1(n_705), .B2(n_706), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_284), .A2(n_318), .B1(n_810), .B2(n_811), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_284), .A2(n_318), .B1(n_856), .B2(n_857), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_284), .A2(n_318), .B1(n_932), .B2(n_933), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_284), .A2(n_318), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
AND2x6_ASAP7_75t_L g322 ( .A(n_285), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g430 ( .A(n_285), .B(n_288), .Y(n_430) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g309 ( .A(n_286), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_287), .Y(n_298) );
INVx1_ASAP7_75t_L g302 ( .A(n_287), .Y(n_302) );
AND2x2_ASAP7_75t_L g412 ( .A(n_287), .B(n_331), .Y(n_412) );
INVx2_ASAP7_75t_L g423 ( .A(n_287), .Y(n_423) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g402 ( .A(n_289), .Y(n_402) );
INVx2_ASAP7_75t_L g657 ( .A(n_289), .Y(n_657) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_289), .Y(n_746) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_289), .Y(n_909) );
INVx2_ASAP7_75t_L g961 ( .A(n_289), .Y(n_961) );
INVx2_ASAP7_75t_SL g1389 ( .A(n_289), .Y(n_1389) );
INVx6_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g296 ( .A(n_290), .B(n_297), .Y(n_296) );
BUFx2_ASAP7_75t_L g415 ( .A(n_290), .Y(n_415) );
INVx2_ASAP7_75t_L g464 ( .A(n_290), .Y(n_464) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_290), .B(n_1254), .Y(n_1295) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g315 ( .A(n_291), .Y(n_315) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g305 ( .A(n_292), .B(n_294), .Y(n_305) );
AND2x4_ASAP7_75t_L g319 ( .A(n_292), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g312 ( .A(n_293), .Y(n_312) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g324 ( .A(n_294), .B(n_325), .Y(n_324) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_295), .A2(n_366), .B1(n_368), .B2(n_372), .Y(n_365) );
AOI22xp5_ASAP7_75t_SL g428 ( .A1(n_296), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_428) );
INVx4_ASAP7_75t_L g531 ( .A(n_296), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_296), .A2(n_322), .B1(n_631), .B2(n_632), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_296), .A2(n_322), .B1(n_708), .B2(n_709), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_296), .A2(n_322), .B1(n_327), .B2(n_769), .C(n_774), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_296), .A2(n_322), .B1(n_807), .B2(n_808), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_296), .A2(n_322), .B1(n_859), .B2(n_860), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_296), .A2(n_322), .B1(n_921), .B2(n_935), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_296), .A2(n_322), .B1(n_1356), .B2(n_1357), .Y(n_1355) );
AND2x2_ASAP7_75t_SL g715 ( .A(n_297), .B(n_716), .Y(n_715) );
AND2x4_ASAP7_75t_L g868 ( .A(n_297), .B(n_716), .Y(n_868) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_306), .B(n_307), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_300), .A2(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g980 ( .A(n_300), .Y(n_980) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
AND2x6_ASAP7_75t_L g318 ( .A(n_301), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g328 ( .A(n_301), .Y(n_328) );
INVx1_ASAP7_75t_L g530 ( .A(n_301), .Y(n_530) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x6_ASAP7_75t_L g314 ( .A(n_302), .B(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g327 ( .A(n_304), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g404 ( .A(n_304), .Y(n_404) );
INVx2_ASAP7_75t_L g607 ( .A(n_304), .Y(n_607) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_304), .Y(n_713) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_305), .Y(n_417) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g438 ( .A(n_309), .Y(n_438) );
AOI222xp33_ASAP7_75t_L g533 ( .A1(n_309), .A2(n_314), .B1(n_502), .B2(n_534), .C1(n_536), .C2(n_537), .Y(n_533) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_309), .A2(n_314), .B1(n_600), .B2(n_606), .C1(n_608), .C2(n_609), .Y(n_605) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g716 ( .A(n_311), .Y(n_716) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g1258 ( .A(n_312), .Y(n_1258) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_314), .A2(n_711), .B1(n_712), .B2(n_714), .C1(n_715), .C2(n_717), .Y(n_710) );
AOI222xp33_ASAP7_75t_L g771 ( .A1(n_314), .A2(n_712), .B1(n_715), .B2(n_764), .C1(n_766), .C2(n_772), .Y(n_771) );
AOI222xp33_ASAP7_75t_L g812 ( .A1(n_314), .A2(n_715), .B1(n_813), .B2(n_814), .C1(n_815), .C2(n_816), .Y(n_812) );
AOI222xp33_ASAP7_75t_L g861 ( .A1(n_314), .A2(n_862), .B1(n_863), .B2(n_866), .C1(n_867), .C2(n_869), .Y(n_861) );
AOI222xp33_ASAP7_75t_L g936 ( .A1(n_314), .A2(n_867), .B1(n_924), .B2(n_926), .C1(n_937), .C2(n_938), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_314), .A2(n_868), .B1(n_982), .B2(n_983), .Y(n_981) );
AOI222xp33_ASAP7_75t_L g1351 ( .A1(n_314), .A2(n_403), .B1(n_868), .B2(n_1352), .C1(n_1353), .C2(n_1354), .Y(n_1351) );
BUFx3_ASAP7_75t_L g1261 ( .A(n_315), .Y(n_1261) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_321), .B2(n_322), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_318), .A2(n_322), .B1(n_433), .B2(n_434), .Y(n_432) );
CKINVDCx6p67_ASAP7_75t_R g540 ( .A(n_318), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_318), .A2(n_430), .B1(n_628), .B2(n_629), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_318), .A2(n_430), .B1(n_776), .B2(n_777), .Y(n_775) );
INVx2_ASAP7_75t_SL g407 ( .A(n_319), .Y(n_407) );
BUFx3_ASAP7_75t_L g419 ( .A(n_319), .Y(n_419) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_319), .Y(n_516) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_319), .Y(n_526) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_319), .Y(n_568) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_319), .Y(n_583) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_319), .Y(n_667) );
BUFx2_ASAP7_75t_L g749 ( .A(n_319), .Y(n_749) );
INVx1_ASAP7_75t_L g510 ( .A(n_320), .Y(n_510) );
INVx4_ASAP7_75t_L g541 ( .A(n_322), .Y(n_541) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_323), .Y(n_420) );
INVx2_ASAP7_75t_L g585 ( .A(n_323), .Y(n_585) );
BUFx6f_ASAP7_75t_L g750 ( .A(n_323), .Y(n_750) );
INVx1_ASAP7_75t_L g793 ( .A(n_323), .Y(n_793) );
INVx1_ASAP7_75t_L g835 ( .A(n_323), .Y(n_835) );
INVx1_ASAP7_75t_L g1394 ( .A(n_323), .Y(n_1394) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_324), .Y(n_408) );
INVx2_ASAP7_75t_L g664 ( .A(n_324), .Y(n_664) );
INVx1_ASAP7_75t_L g965 ( .A(n_324), .Y(n_965) );
INVx1_ASAP7_75t_L g1249 ( .A(n_324), .Y(n_1249) );
INVx1_ASAP7_75t_L g509 ( .A(n_325), .Y(n_509) );
NAND4xp25_ASAP7_75t_L g427 ( .A(n_326), .B(n_428), .C(n_432), .D(n_435), .Y(n_427) );
NAND4xp25_ASAP7_75t_L g805 ( .A(n_326), .B(n_806), .C(n_809), .D(n_812), .Y(n_805) );
BUFx2_ASAP7_75t_L g870 ( .A(n_326), .Y(n_870) );
NAND4xp25_ASAP7_75t_L g930 ( .A(n_326), .B(n_931), .C(n_934), .D(n_936), .Y(n_930) );
INVx5_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
CKINVDCx8_ASAP7_75t_R g538 ( .A(n_327), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_327), .B(n_623), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_329), .A2(n_427), .B(n_439), .C(n_452), .Y(n_426) );
OAI31xp33_ASAP7_75t_SL g527 ( .A1(n_329), .A2(n_528), .A3(n_532), .B(n_539), .Y(n_527) );
OAI31xp33_ASAP7_75t_L g601 ( .A1(n_329), .A2(n_602), .A3(n_603), .B(n_604), .Y(n_601) );
AOI211xp5_ASAP7_75t_L g804 ( .A1(n_329), .A2(n_805), .B(n_817), .C(n_836), .Y(n_804) );
OAI31xp33_ASAP7_75t_L g977 ( .A1(n_329), .A2(n_978), .A3(n_979), .B(n_984), .Y(n_977) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
AND2x4_ASAP7_75t_L g634 ( .A(n_330), .B(n_332), .Y(n_634) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g422 ( .A(n_331), .B(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g388 ( .A(n_333), .Y(n_388) );
OR2x6_ASAP7_75t_L g474 ( .A(n_333), .B(n_475), .Y(n_474) );
AOI31xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_354), .A3(n_365), .B(n_373), .Y(n_334) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B(n_342), .C(n_347), .Y(n_335) );
AOI222xp33_ASAP7_75t_L g1011 ( .A1(n_337), .A2(n_349), .B1(n_550), .B2(n_982), .C1(n_983), .C2(n_1007), .Y(n_1011) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x6_ASAP7_75t_L g1305 ( .A(n_338), .B(n_1302), .Y(n_1305) );
NAND2x1p5_ASAP7_75t_L g1322 ( .A(n_338), .B(n_1316), .Y(n_1322) );
BUFx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g342 ( .A(n_339), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_339), .Y(n_444) );
BUFx2_ASAP7_75t_L g643 ( .A(n_339), .Y(n_643) );
BUFx3_ASAP7_75t_L g695 ( .A(n_339), .Y(n_695) );
BUFx6f_ASAP7_75t_L g821 ( .A(n_339), .Y(n_821) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g440 ( .A1(n_342), .A2(n_441), .B(n_442), .C(n_445), .Y(n_440) );
CKINVDCx11_ASAP7_75t_R g548 ( .A(n_342), .Y(n_548) );
AOI211xp5_ASAP7_75t_L g719 ( .A1(n_342), .A2(n_720), .B(n_722), .C(n_723), .Y(n_719) );
AOI211xp5_ASAP7_75t_L g837 ( .A1(n_342), .A2(n_838), .B(n_839), .C(n_840), .Y(n_837) );
AOI211xp5_ASAP7_75t_L g1364 ( .A1(n_342), .A2(n_385), .B(n_1365), .C(n_1366), .Y(n_1364) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVxp67_ASAP7_75t_L g552 ( .A(n_344), .Y(n_552) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_345), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g359 ( .A(n_346), .Y(n_359) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g446 ( .A(n_349), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_349), .A2(n_536), .B1(n_537), .B2(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_349), .A2(n_550), .B1(n_608), .B2(n_609), .Y(n_613) );
INVx2_ASAP7_75t_L g646 ( .A(n_349), .Y(n_646) );
INVx1_ASAP7_75t_L g1315 ( .A(n_350), .Y(n_1315) );
INVx1_ASAP7_75t_L g551 ( .A(n_352), .Y(n_551) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_353), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g501 ( .A(n_353), .B(n_481), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_356), .B1(n_357), .B2(n_364), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_355), .A2(n_357), .B1(n_448), .B2(n_449), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_355), .A2(n_631), .B1(n_650), .B2(n_651), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_355), .A2(n_366), .B1(n_708), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_355), .A2(n_366), .B1(n_768), .B2(n_769), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g845 ( .A1(n_355), .A2(n_651), .B1(n_807), .B2(n_846), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_355), .A2(n_366), .B1(n_859), .B2(n_879), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g927 ( .A1(n_355), .A2(n_726), .B1(n_928), .B2(n_929), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_355), .A2(n_651), .B1(n_1006), .B2(n_1013), .Y(n_1012) );
AOI22xp5_ASAP7_75t_L g1362 ( .A1(n_355), .A2(n_366), .B1(n_1356), .B2(n_1363), .Y(n_1362) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_357), .A2(n_368), .B1(n_637), .B2(n_638), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_357), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_357), .A2(n_726), .B1(n_760), .B2(n_761), .Y(n_759) );
AOI22xp33_ASAP7_75t_SL g842 ( .A1(n_357), .A2(n_726), .B1(n_843), .B2(n_844), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_357), .A2(n_726), .B1(n_873), .B2(n_874), .Y(n_872) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_357), .A2(n_651), .B1(n_921), .B2(n_922), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g1367 ( .A1(n_357), .A2(n_368), .B1(n_1368), .B2(n_1369), .Y(n_1367) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
AND2x4_ASAP7_75t_L g368 ( .A(n_358), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g555 ( .A(n_358), .Y(n_555) );
AND2x4_ASAP7_75t_L g726 ( .A(n_358), .B(n_369), .Y(n_726) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_360), .Y(n_378) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_360), .Y(n_392) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_360), .Y(n_459) );
BUFx2_ASAP7_75t_L g674 ( .A(n_360), .Y(n_674) );
INVx1_ASAP7_75t_L g686 ( .A(n_360), .Y(n_686) );
INVx1_ASAP7_75t_L g785 ( .A(n_360), .Y(n_785) );
BUFx2_ASAP7_75t_L g952 ( .A(n_360), .Y(n_952) );
AND2x4_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g1320 ( .A(n_361), .Y(n_1320) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_366), .A2(n_368), .B1(n_431), .B2(n_451), .Y(n_450) );
INVx5_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx4_ASAP7_75t_L g651 ( .A(n_367), .Y(n_651) );
INVx5_ASAP7_75t_SL g544 ( .A(n_368), .Y(n_544) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_370), .Y(n_394) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_371), .Y(n_379) );
INVx3_ASAP7_75t_L g491 ( .A(n_371), .Y(n_491) );
INVx1_ASAP7_75t_L g678 ( .A(n_371), .Y(n_678) );
AOI31xp33_ASAP7_75t_L g439 ( .A1(n_373), .A2(n_440), .A3(n_447), .B(n_450), .Y(n_439) );
AOI31xp33_ASAP7_75t_L g1361 ( .A1(n_373), .A2(n_1362), .A3(n_1364), .B(n_1367), .Y(n_1361) );
AND2x4_ASAP7_75t_L g421 ( .A(n_374), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g518 ( .A(n_374), .B(n_422), .Y(n_518) );
AND2x4_ASAP7_75t_L g1294 ( .A(n_374), .B(n_1295), .Y(n_1294) );
NAND4xp25_ASAP7_75t_L g375 ( .A(n_376), .B(n_390), .C(n_400), .D(n_413), .Y(n_375) );
NAND3xp33_ASAP7_75t_L g376 ( .A(n_377), .B(n_380), .C(n_387), .Y(n_376) );
INVx2_ASAP7_75t_SL g884 ( .A(n_379), .Y(n_884) );
INVx4_ASAP7_75t_L g893 ( .A(n_379), .Y(n_893) );
INVx2_ASAP7_75t_SL g954 ( .A(n_379), .Y(n_954) );
BUFx3_ASAP7_75t_L g987 ( .A(n_379), .Y(n_987) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g456 ( .A(n_382), .Y(n_456) );
INVx2_ASAP7_75t_SL g787 ( .A(n_382), .Y(n_787) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx2_ASAP7_75t_L g826 ( .A(n_383), .Y(n_826) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx3_ASAP7_75t_L g682 ( .A(n_384), .Y(n_682) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_387), .B(n_454), .C(n_455), .Y(n_453) );
AOI33xp33_ASAP7_75t_L g668 ( .A1(n_387), .A2(n_669), .A3(n_673), .B1(n_679), .B2(n_684), .B3(n_690), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g736 ( .A(n_387), .B(n_737), .C(n_739), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g779 ( .A(n_387), .B(n_780), .C(n_781), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g818 ( .A(n_387), .B(n_819), .C(n_820), .Y(n_818) );
INVx2_ASAP7_75t_L g889 ( .A(n_387), .Y(n_889) );
BUFx3_ASAP7_75t_L g991 ( .A(n_387), .Y(n_991) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
AND2x2_ASAP7_75t_L g396 ( .A(n_388), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g410 ( .A(n_388), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g563 ( .A(n_388), .B(n_564), .Y(n_563) );
OR2x6_ASAP7_75t_L g905 ( .A(n_388), .B(n_564), .Y(n_905) );
BUFx2_ASAP7_75t_L g1286 ( .A(n_388), .Y(n_1286) );
AND2x4_ASAP7_75t_L g1373 ( .A(n_388), .B(n_389), .Y(n_1373) );
NAND3xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .C(n_396), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_396), .B(n_458), .C(n_460), .Y(n_457) );
INVx1_ASAP7_75t_L g503 ( .A(n_396), .Y(n_503) );
NAND3xp33_ASAP7_75t_L g782 ( .A(n_396), .B(n_783), .C(n_786), .Y(n_782) );
NAND3xp33_ASAP7_75t_L g822 ( .A(n_396), .B(n_823), .C(n_825), .Y(n_822) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x6_ASAP7_75t_L g670 ( .A(n_398), .B(n_671), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_405), .C(n_409), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g830 ( .A(n_407), .Y(n_830) );
INVx1_ASAP7_75t_L g570 ( .A(n_408), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_409), .B(n_462), .C(n_465), .Y(n_461) );
AOI33xp33_ASAP7_75t_L g653 ( .A1(n_409), .A2(n_654), .A3(n_655), .B1(n_659), .B2(n_665), .B3(n_666), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_409), .B(n_744), .C(n_748), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g788 ( .A(n_409), .B(n_789), .C(n_791), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g827 ( .A(n_409), .B(n_828), .C(n_829), .Y(n_827) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI22xp5_ASAP7_75t_SL g504 ( .A1(n_410), .A2(n_505), .B1(n_517), .B2(n_519), .Y(n_504) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g564 ( .A(n_412), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_418), .C(n_421), .Y(n_413) );
INVx1_ASAP7_75t_L g973 ( .A(n_416), .Y(n_973) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_SL g535 ( .A(n_417), .Y(n_535) );
BUFx4f_ASAP7_75t_L g747 ( .A(n_417), .Y(n_747) );
BUFx3_ASAP7_75t_L g814 ( .A(n_417), .Y(n_814) );
AND2x4_ASAP7_75t_L g1264 ( .A(n_417), .B(n_1265), .Y(n_1264) );
AND2x4_ASAP7_75t_L g1273 ( .A(n_417), .B(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1391 ( .A(n_417), .Y(n_1391) );
INVx2_ASAP7_75t_SL g970 ( .A(n_419), .Y(n_970) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_421), .B(n_467), .C(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g587 ( .A(n_421), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_421), .B(n_752), .C(n_753), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g794 ( .A(n_421), .B(n_795), .C(n_797), .Y(n_794) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_421), .B(n_832), .C(n_833), .Y(n_831) );
AOI33xp33_ASAP7_75t_L g1382 ( .A1(n_421), .A2(n_1383), .A3(n_1384), .B1(n_1385), .B2(n_1386), .B3(n_1392), .Y(n_1382) );
CKINVDCx5p33_ASAP7_75t_R g1252 ( .A(n_422), .Y(n_1252) );
AND2x4_ASAP7_75t_L g1254 ( .A(n_423), .B(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g742 ( .A(n_443), .Y(n_742) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_444), .Y(n_683) );
INVx1_ASAP7_75t_L g765 ( .A(n_446), .Y(n_765) );
NAND4xp25_ASAP7_75t_L g452 ( .A(n_453), .B(n_457), .C(n_461), .D(n_466), .Y(n_452) );
INVx2_ASAP7_75t_SL g945 ( .A(n_459), .Y(n_945) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_459), .B(n_1302), .Y(n_1310) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_SL g796 ( .A(n_464), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_559), .B1(n_615), .B2(n_616), .Y(n_469) );
INVx1_ASAP7_75t_L g615 ( .A(n_470), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_527), .C(n_542), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_504), .Y(n_472) );
OAI33xp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_476), .A3(n_483), .B1(n_492), .B2(n_497), .B3(n_503), .Y(n_473) );
OAI33xp33_ASAP7_75t_L g588 ( .A1(n_474), .A2(n_503), .A3(n_589), .B1(n_592), .B2(n_593), .B3(n_597), .Y(n_588) );
OAI33xp33_ASAP7_75t_L g1323 ( .A1(n_474), .A2(n_1324), .A3(n_1330), .B1(n_1337), .B2(n_1338), .B3(n_1341), .Y(n_1323) );
OAI22xp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B1(n_479), .B2(n_482), .Y(n_476) );
OAI221xp5_ASAP7_75t_L g505 ( .A1(n_478), .A2(n_482), .B1(n_506), .B2(n_511), .C(n_515), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_479), .A2(n_572), .B1(n_575), .B2(n_590), .Y(n_589) );
BUFx3_ASAP7_75t_L g1335 ( .A(n_479), .Y(n_1335) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI22xp33_ASAP7_75t_SL g483 ( .A1(n_484), .A2(n_485), .B1(n_488), .B2(n_489), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_485), .A2(n_493), .B1(n_494), .B2(n_496), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_485), .A2(n_494), .B1(n_566), .B2(n_569), .Y(n_592) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g594 ( .A(n_486), .Y(n_594) );
INVx1_ASAP7_75t_L g1326 ( .A(n_486), .Y(n_1326) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g556 ( .A(n_487), .Y(n_556) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g1377 ( .A(n_490), .Y(n_1377) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g495 ( .A(n_491), .Y(n_495) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_491), .Y(n_734) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_494), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_593) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g947 ( .A(n_495), .Y(n_947) );
AND2x4_ASAP7_75t_L g1301 ( .A(n_495), .B(n_1302), .Y(n_1301) );
BUFx3_ASAP7_75t_L g1343 ( .A(n_495), .Y(n_1343) );
OAI22xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B1(n_500), .B2(n_502), .Y(n_497) );
OAI22xp33_ASAP7_75t_L g988 ( .A1(n_498), .A2(n_599), .B1(n_989), .B2(n_990), .Y(n_988) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g547 ( .A(n_501), .Y(n_547) );
INVx3_ASAP7_75t_L g599 ( .A(n_501), .Y(n_599) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g520 ( .A(n_507), .Y(n_520) );
INVx2_ASAP7_75t_L g1001 ( .A(n_507), .Y(n_1001) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g529 ( .A(n_508), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g574 ( .A(n_508), .Y(n_574) );
OR2x2_ASAP7_75t_L g1278 ( .A(n_508), .B(n_1266), .Y(n_1278) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
AND2x2_ASAP7_75t_L g514 ( .A(n_509), .B(n_510), .Y(n_514) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g523 ( .A(n_514), .Y(n_523) );
BUFx4f_ASAP7_75t_L g577 ( .A(n_514), .Y(n_577) );
INVx1_ASAP7_75t_L g626 ( .A(n_514), .Y(n_626) );
INVx2_ASAP7_75t_L g1003 ( .A(n_514), .Y(n_1003) );
INVx1_ASAP7_75t_L g967 ( .A(n_517), .Y(n_967) );
OAI22xp5_ASAP7_75t_SL g999 ( .A1(n_517), .A2(n_563), .B1(n_1000), .B2(n_1005), .Y(n_999) );
INVx4_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx4f_ASAP7_75t_L g654 ( .A(n_518), .Y(n_654) );
BUFx4f_ASAP7_75t_L g912 ( .A(n_518), .Y(n_912) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B1(n_522), .B2(n_524), .C(n_525), .Y(n_519) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g902 ( .A(n_526), .Y(n_902) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_533), .B(n_538), .Y(n_532) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g658 ( .A(n_535), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_538), .B(n_605), .Y(n_604) );
NAND4xp25_ASAP7_75t_L g703 ( .A(n_538), .B(n_704), .C(n_707), .D(n_710), .Y(n_703) );
NAND4xp25_ASAP7_75t_SL g1350 ( .A(n_538), .B(n_1351), .C(n_1355), .D(n_1358), .Y(n_1350) );
OAI31xp33_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_545), .A3(n_553), .B(n_557), .Y(n_542) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g1340 ( .A(n_547), .Y(n_1340) );
NAND4xp25_ASAP7_75t_SL g635 ( .A(n_548), .B(n_636), .C(n_639), .D(n_649), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g758 ( .A(n_548), .B(n_759), .C(n_762), .D(n_767), .Y(n_758) );
NAND4xp25_ASAP7_75t_SL g871 ( .A(n_548), .B(n_872), .C(n_875), .D(n_878), .Y(n_871) );
NAND4xp25_ASAP7_75t_L g919 ( .A(n_548), .B(n_920), .C(n_923), .D(n_927), .Y(n_919) );
NAND3xp33_ASAP7_75t_L g1010 ( .A(n_548), .B(n_1011), .C(n_1012), .Y(n_1010) );
AOI222xp33_ASAP7_75t_L g875 ( .A1(n_550), .A2(n_645), .B1(n_866), .B2(n_869), .C1(n_876), .C2(n_877), .Y(n_875) );
AOI222xp33_ASAP7_75t_L g923 ( .A1(n_550), .A2(n_645), .B1(n_839), .B2(n_924), .C1(n_925), .C2(n_926), .Y(n_923) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AND2x4_ASAP7_75t_L g648 ( .A(n_551), .B(n_552), .Y(n_648) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
OAI31xp33_ASAP7_75t_SL g610 ( .A1(n_557), .A2(n_611), .A3(n_612), .B(n_614), .Y(n_610) );
AOI221x1_ASAP7_75t_L g620 ( .A1(n_557), .A2(n_621), .B1(n_633), .B2(n_635), .C(n_652), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_557), .A2(n_634), .B1(n_703), .B2(n_718), .C(n_730), .Y(n_702) );
AOI221x1_ASAP7_75t_L g757 ( .A1(n_557), .A2(n_634), .B1(n_758), .B2(n_770), .C(n_778), .Y(n_757) );
AOI221x1_ASAP7_75t_L g853 ( .A1(n_557), .A2(n_633), .B1(n_854), .B2(n_871), .C(n_880), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g918 ( .A1(n_557), .A2(n_919), .B1(n_930), .B2(n_939), .C(n_941), .Y(n_918) );
OAI21xp5_ASAP7_75t_L g1009 ( .A1(n_557), .A2(n_1010), .B(n_1014), .Y(n_1009) );
CKINVDCx16_ASAP7_75t_R g557 ( .A(n_558), .Y(n_557) );
AOI31xp33_ASAP7_75t_L g836 ( .A1(n_558), .A2(n_837), .A3(n_842), .B(n_845), .Y(n_836) );
INVx1_ASAP7_75t_L g616 ( .A(n_559), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_601), .C(n_610), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_588), .Y(n_561) );
OAI33xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .A3(n_571), .B1(n_578), .B2(n_581), .B3(n_587), .Y(n_562) );
INVx1_ASAP7_75t_L g1270 ( .A(n_564), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B1(n_569), .B2(n_570), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx4f_ASAP7_75t_L g660 ( .A(n_568), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_575), .B2(n_576), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_573), .A2(n_576), .B1(n_579), .B2(n_580), .Y(n_578) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_584), .B1(n_585), .B2(n_586), .Y(n_581) );
INVx1_ASAP7_75t_L g963 ( .A(n_582), .Y(n_963) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g1284 ( .A(n_583), .B(n_1265), .Y(n_1284) );
INVx1_ASAP7_75t_L g903 ( .A(n_585), .Y(n_903) );
INVx1_ASAP7_75t_L g911 ( .A(n_585), .Y(n_911) );
OAI22xp33_ASAP7_75t_L g597 ( .A1(n_590), .A2(n_598), .B1(n_599), .B2(n_600), .Y(n_597) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI22xp33_ASAP7_75t_SL g993 ( .A1(n_599), .A2(n_994), .B1(n_995), .B2(n_997), .Y(n_993) );
INVx3_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g865 ( .A(n_607), .Y(n_865) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_627), .C(n_630), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g940 ( .A(n_634), .Y(n_940) );
AOI211x1_ASAP7_75t_SL g1349 ( .A1(n_634), .A2(n_1350), .B(n_1361), .C(n_1370), .Y(n_1349) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_641), .B1(n_644), .B2(n_645), .C1(n_647), .C2(n_648), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g877 ( .A(n_642), .Y(n_877) );
INVx1_ASAP7_75t_L g887 ( .A(n_642), .Y(n_887) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI222xp33_ASAP7_75t_L g762 ( .A1(n_643), .A2(n_648), .B1(n_763), .B2(n_764), .C1(n_765), .C2(n_766), .Y(n_762) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_668), .Y(n_652) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_SL g754 ( .A(n_662), .Y(n_754) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g1272 ( .A(n_664), .Y(n_1272) );
OR2x2_ASAP7_75t_L g1281 ( .A(n_664), .B(n_1266), .Y(n_1281) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_669), .B(n_732), .C(n_735), .Y(n_731) );
NAND3xp33_ASAP7_75t_L g890 ( .A(n_669), .B(n_891), .C(n_894), .Y(n_890) );
NAND3xp33_ASAP7_75t_L g950 ( .A(n_669), .B(n_951), .C(n_955), .Y(n_950) );
CKINVDCx8_ASAP7_75t_R g1337 ( .A(n_669), .Y(n_1337) );
AOI33xp33_ASAP7_75t_L g1371 ( .A1(n_669), .A2(n_1372), .A3(n_1374), .B1(n_1375), .B2(n_1378), .B3(n_1379), .Y(n_1371) );
INVx5_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx6_ASAP7_75t_L g998 ( .A(n_670), .Y(n_998) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x4_ASAP7_75t_L g1302 ( .A(n_672), .B(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g738 ( .A(n_676), .Y(n_738) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g689 ( .A(n_678), .Y(n_689) );
BUFx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_SL g692 ( .A(n_682), .Y(n_692) );
INVx2_ASAP7_75t_L g886 ( .A(n_682), .Y(n_886) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g1328 ( .A(n_689), .Y(n_1328) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g741 ( .A(n_692), .Y(n_741) );
INVx1_ASAP7_75t_L g896 ( .A(n_692), .Y(n_896) );
AND2x4_ASAP7_75t_L g1308 ( .A(n_692), .B(n_1302), .Y(n_1308) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_695), .Y(n_721) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
XNOR2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_849), .Y(n_698) );
AO22x2_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_801), .B1(n_847), .B2(n_848), .Y(n_699) );
INVx1_ASAP7_75t_L g847 ( .A(n_700), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_755), .B1(n_756), .B2(n_800), .Y(n_700) );
INVx1_ASAP7_75t_L g800 ( .A(n_701), .Y(n_800) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_724), .C(n_728), .Y(n_718) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND4xp25_ASAP7_75t_L g730 ( .A(n_731), .B(n_736), .C(n_743), .D(n_751), .Y(n_730) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_SL g824 ( .A(n_734), .Y(n_824) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g790 ( .A(n_746), .Y(n_790) );
INVx4_ASAP7_75t_L g899 ( .A(n_746), .Y(n_899) );
BUFx2_ASAP7_75t_L g938 ( .A(n_747), .Y(n_938) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g799 ( .A(n_757), .Y(n_799) );
NAND3xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .C(n_775), .Y(n_770) );
NAND4xp25_ASAP7_75t_L g778 ( .A(n_779), .B(n_782), .C(n_788), .D(n_794), .Y(n_778) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g1380 ( .A(n_785), .Y(n_1380) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g848 ( .A(n_801), .Y(n_848) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND4xp25_ASAP7_75t_L g817 ( .A(n_818), .B(n_822), .C(n_827), .D(n_831), .Y(n_817) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_821), .Y(n_839) );
INVx2_ASAP7_75t_SL g957 ( .A(n_821), .Y(n_957) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
XNOR2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_915), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g914 ( .A(n_853), .Y(n_914) );
NAND4xp25_ASAP7_75t_L g854 ( .A(n_855), .B(n_858), .C(n_861), .D(n_870), .Y(n_854) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
BUFx4f_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
NAND4xp25_ASAP7_75t_L g880 ( .A(n_881), .B(n_890), .C(n_897), .D(n_906), .Y(n_880) );
NAND3xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_885), .C(n_888), .Y(n_881) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
BUFx3_ASAP7_75t_L g949 ( .A(n_886), .Y(n_949) );
NAND3xp33_ASAP7_75t_L g942 ( .A(n_888), .B(n_943), .C(n_948), .Y(n_942) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
NAND3xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_900), .C(n_904), .Y(n_897) );
INVx2_ASAP7_75t_SL g901 ( .A(n_902), .Y(n_901) );
NAND3xp33_ASAP7_75t_L g958 ( .A(n_904), .B(n_959), .C(n_962), .Y(n_958) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_905), .Y(n_904) );
INVx2_ASAP7_75t_L g1383 ( .A(n_905), .Y(n_1383) );
NAND3xp33_ASAP7_75t_L g906 ( .A(n_907), .B(n_910), .C(n_912), .Y(n_906) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
XNOR2x2_ASAP7_75t_L g915 ( .A(n_916), .B(n_974), .Y(n_915) );
XNOR2xp5_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
NAND4xp25_ASAP7_75t_L g941 ( .A(n_942), .B(n_950), .C(n_958), .D(n_966), .Y(n_941) );
INVx3_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVxp67_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx2_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
BUFx3_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
NAND3xp33_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .C(n_971), .Y(n_966) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
XNOR2xp5_ASAP7_75t_L g974 ( .A(n_975), .B(n_976), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g1071 ( .A1(n_975), .A2(n_1020), .B1(n_1036), .B2(n_1072), .Y(n_1071) );
NAND3x1_ASAP7_75t_SL g976 ( .A(n_977), .B(n_985), .C(n_1009), .Y(n_976) );
AOI221xp5_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_991), .B1(n_992), .B2(n_998), .C(n_999), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g1000 ( .A1(n_989), .A2(n_990), .B1(n_1001), .B2(n_1002), .C(n_1004), .Y(n_1000) );
INVx3_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
OAI221xp5_ASAP7_75t_L g1005 ( .A1(n_1001), .A2(n_1002), .B1(n_1006), .B2(n_1007), .C(n_1008), .Y(n_1005) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
OAI21xp5_ASAP7_75t_L g1015 ( .A1(n_1016), .A2(n_1026), .B(n_1239), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
OAI22xp33_ASAP7_75t_L g1134 ( .A1(n_1018), .A2(n_1135), .B1(n_1136), .B2(n_1137), .Y(n_1134) );
BUFx3_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_1019), .A2(n_1033), .B1(n_1034), .B2(n_1038), .Y(n_1032) );
BUFx6f_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1022), .Y(n_1020) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_1021), .B(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1021), .Y(n_1055) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1022), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1025), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1025), .Y(n_1043) );
AOI221xp5_ASAP7_75t_L g1026 ( .A1(n_1027), .A2(n_1130), .B1(n_1131), .B2(n_1138), .C(n_1178), .Y(n_1026) );
A2O1A1Ixp33_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1073), .B(n_1099), .C(n_1107), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1049), .Y(n_1028) );
INVxp67_ASAP7_75t_L g1084 ( .A(n_1029), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1030), .B(n_1077), .Y(n_1076) );
INVx2_ASAP7_75t_SL g1096 ( .A(n_1030), .Y(n_1096) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1030), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1030), .B(n_1051), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1030), .B(n_1050), .Y(n_1155) );
NOR2xp33_ASAP7_75t_L g1186 ( .A(n_1030), .B(n_1050), .Y(n_1186) );
AND2x4_ASAP7_75t_L g1198 ( .A(n_1030), .B(n_1093), .Y(n_1198) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_1031), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1031), .B(n_1093), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1031), .B(n_1077), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1039), .Y(n_1031) );
HB1xp67_ASAP7_75t_L g1137 ( .A(n_1034), .Y(n_1137) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1037), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_1040), .A2(n_1045), .B1(n_1046), .B2(n_1048), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
BUFx3_ASAP7_75t_L g1133 ( .A(n_1041), .Y(n_1133) );
AND2x4_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1044), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1042), .B(n_1044), .Y(n_1064) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
AND2x4_ASAP7_75t_L g1047 ( .A(n_1043), .B(n_1044), .Y(n_1047) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1046), .Y(n_1106) );
INVx2_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1049), .B(n_1172), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1059), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1050), .B(n_1087), .Y(n_1086) );
NAND3xp33_ASAP7_75t_L g1184 ( .A(n_1050), .B(n_1070), .C(n_1132), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1050), .B(n_1080), .Y(n_1217) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
BUFx2_ASAP7_75t_L g1075 ( .A(n_1051), .Y(n_1075) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1051), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1051), .B(n_1080), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1051), .B(n_1092), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1051), .B(n_1088), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1051), .B(n_1124), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1051), .B(n_1060), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1058), .Y(n_1051) );
AND2x4_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1055), .Y(n_1053) );
OAI21xp33_ASAP7_75t_SL g1401 ( .A1(n_1054), .A2(n_1400), .B(n_1402), .Y(n_1401) );
AND2x4_ASAP7_75t_L g1056 ( .A(n_1055), .B(n_1057), .Y(n_1056) );
BUFx2_ASAP7_75t_L g1104 ( .A(n_1056), .Y(n_1104) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1059), .Y(n_1174) );
NOR2xp33_ASAP7_75t_L g1182 ( .A(n_1059), .B(n_1080), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1065), .Y(n_1059) );
OR2x2_ASAP7_75t_L g1128 ( .A(n_1060), .B(n_1089), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1060), .B(n_1157), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1060), .B(n_1069), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1060), .B(n_1070), .Y(n_1226) );
BUFx3_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVxp67_ASAP7_75t_L g1081 ( .A(n_1061), .Y(n_1081) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_1061), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1061), .B(n_1120), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_1061), .B(n_1070), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1063), .Y(n_1061) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1065), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1065), .B(n_1081), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1069), .Y(n_1065) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1066), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1066), .B(n_1070), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_1066), .B(n_1070), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1068), .Y(n_1066) );
AOI221xp5_ASAP7_75t_L g1073 ( .A1(n_1069), .A2(n_1074), .B1(n_1080), .B2(n_1084), .C(n_1085), .Y(n_1073) );
NOR2x1_ASAP7_75t_L g1140 ( .A(n_1069), .B(n_1088), .Y(n_1140) );
INVx2_ASAP7_75t_SL g1069 ( .A(n_1070), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1070), .B(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1074), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1076), .Y(n_1074) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1075), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1075), .B(n_1161), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1075), .B(n_1087), .Y(n_1176) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1076), .Y(n_1117) );
OAI221xp5_ASAP7_75t_L g1085 ( .A1(n_1077), .A2(n_1086), .B1(n_1089), .B2(n_1091), .C(n_1094), .Y(n_1085) );
INVx3_ASAP7_75t_L g1093 ( .A(n_1077), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1077), .B(n_1101), .Y(n_1111) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1077), .B(n_1102), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1079), .Y(n_1077) );
O2A1O1Ixp33_ASAP7_75t_L g1214 ( .A1(n_1080), .A2(n_1141), .B(n_1199), .C(n_1215), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1082), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1081), .B(n_1120), .Y(n_1119) );
AOI322xp5_ASAP7_75t_L g1145 ( .A1(n_1081), .A2(n_1093), .A3(n_1146), .B1(n_1150), .B2(n_1152), .C1(n_1153), .C2(n_1156), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1081), .B(n_1211), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1082), .B(n_1097), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1082), .B(n_1088), .Y(n_1115) );
OAI21xp33_ASAP7_75t_L g1129 ( .A1(n_1082), .A2(n_1087), .B(n_1095), .Y(n_1129) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1082), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1082), .B(n_1195), .Y(n_1194) );
NOR2xp33_ASAP7_75t_L g1087 ( .A(n_1083), .B(n_1088), .Y(n_1087) );
AOI21xp5_ASAP7_75t_L g1094 ( .A1(n_1083), .A2(n_1095), .B(n_1098), .Y(n_1094) );
NAND4xp25_ASAP7_75t_L g1185 ( .A(n_1083), .B(n_1132), .C(n_1172), .D(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1087), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1088), .B(n_1090), .Y(n_1236) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1090), .B(n_1097), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1090), .B(n_1238), .Y(n_1237) );
OAI222xp33_ASAP7_75t_SL g1230 ( .A1(n_1091), .A2(n_1170), .B1(n_1231), .B2(n_1233), .C1(n_1235), .C2(n_1237), .Y(n_1230) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1093), .Y(n_1152) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1093), .B(n_1193), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1093), .B(n_1102), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1095), .B(n_1164), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1097), .Y(n_1095) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1096), .Y(n_1114) );
NOR2xp33_ASAP7_75t_L g1150 ( .A(n_1096), .B(n_1151), .Y(n_1150) );
NOR2xp33_ASAP7_75t_L g1191 ( .A(n_1096), .B(n_1192), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1096), .B(n_1228), .Y(n_1227) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1097), .B(n_1121), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1097), .B(n_1198), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1097), .B(n_1226), .Y(n_1225) );
O2A1O1Ixp33_ASAP7_75t_L g1223 ( .A1(n_1099), .A2(n_1152), .B(n_1224), .C(n_1227), .Y(n_1223) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1100), .B(n_1110), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1100), .B(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1101), .Y(n_1165) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1102), .Y(n_1124) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1102), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1105), .Y(n_1102) );
NOR3xp33_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1116), .C(n_1125), .Y(n_1107) );
OAI21xp33_ASAP7_75t_L g1108 ( .A1(n_1109), .A2(n_1112), .B(n_1113), .Y(n_1108) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1109), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1110), .B(n_1234), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1111), .B(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1111), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1115), .Y(n_1113) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1115), .Y(n_1122) );
AOI22xp5_ASAP7_75t_L g1171 ( .A1(n_1115), .A2(n_1172), .B1(n_1173), .B2(n_1177), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1115), .B(n_1155), .Y(n_1215) );
O2A1O1Ixp33_ASAP7_75t_L g1116 ( .A1(n_1117), .A2(n_1118), .B(n_1122), .C(n_1123), .Y(n_1116) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
A2O1A1Ixp33_ASAP7_75t_L g1205 ( .A1(n_1122), .A2(n_1206), .B(n_1207), .C(n_1209), .Y(n_1205) );
NOR3xp33_ASAP7_75t_L g1153 ( .A(n_1123), .B(n_1148), .C(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
A2O1A1Ixp33_ASAP7_75t_L g1139 ( .A1(n_1124), .A2(n_1140), .B(n_1141), .C(n_1143), .Y(n_1139) );
OAI21xp33_ASAP7_75t_L g1125 ( .A1(n_1126), .A2(n_1128), .B(n_1129), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1127), .B(n_1203), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1127), .B(n_1140), .Y(n_1229) );
NOR2xp33_ASAP7_75t_L g1167 ( .A(n_1128), .B(n_1168), .Y(n_1167) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
INVx3_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1132), .B(n_1166), .Y(n_1188) );
XNOR2xp5_ASAP7_75t_L g1242 ( .A(n_1135), .B(n_1243), .Y(n_1242) );
NAND4xp25_ASAP7_75t_SL g1138 ( .A(n_1139), .B(n_1145), .C(n_1158), .D(n_1171), .Y(n_1138) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1149), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1148), .B(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1151), .Y(n_1172) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
O2A1O1Ixp33_ASAP7_75t_L g1158 ( .A1(n_1159), .A2(n_1162), .B(n_1166), .C(n_1167), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
CKINVDCx5p33_ASAP7_75t_R g1170 ( .A(n_1161), .Y(n_1170) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1165), .Y(n_1169) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1166), .Y(n_1221) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1170), .Y(n_1168) );
OAI221xp5_ASAP7_75t_SL g1181 ( .A1(n_1170), .A2(n_1182), .B1(n_1183), .B2(n_1184), .C(n_1185), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1175), .Y(n_1173) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
NAND3xp33_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1200), .C(n_1219), .Y(n_1178) );
NOR4xp25_ASAP7_75t_SL g1179 ( .A(n_1180), .B(n_1181), .C(n_1187), .D(n_1196), .Y(n_1179) );
OAI21xp33_ASAP7_75t_L g1187 ( .A1(n_1188), .A2(n_1189), .B(n_1190), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1194), .Y(n_1190) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1192), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1199), .Y(n_1196) );
AOI221xp5_ASAP7_75t_L g1200 ( .A1(n_1198), .A2(n_1201), .B1(n_1204), .B2(n_1205), .C(n_1212), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
OAI21xp5_ASAP7_75t_L g1216 ( .A1(n_1210), .A2(n_1217), .B(n_1218), .Y(n_1216) );
OAI21xp5_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1214), .B(n_1216), .Y(n_1212) );
NOR3xp33_ASAP7_75t_SL g1219 ( .A(n_1220), .B(n_1223), .C(n_1230), .Y(n_1219) );
NOR2xp33_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1222), .Y(n_1220) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1232), .Y(n_1238) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1296), .Y(n_1243) );
AOI22xp5_ASAP7_75t_L g1244 ( .A1(n_1245), .A2(n_1285), .B1(n_1287), .B2(n_1288), .Y(n_1244) );
NAND4xp25_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1263), .C(n_1275), .D(n_1282), .Y(n_1245) );
AOI322xp5_ASAP7_75t_L g1246 ( .A1(n_1247), .A2(n_1250), .A3(n_1251), .B1(n_1253), .B2(n_1259), .C1(n_1260), .C2(n_1262), .Y(n_1246) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
AND2x4_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1257), .Y(n_1253) );
AND2x4_ASAP7_75t_L g1260 ( .A(n_1254), .B(n_1261), .Y(n_1260) );
BUFx2_ASAP7_75t_L g1274 ( .A(n_1254), .Y(n_1274) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx2_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
AOI221xp5_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1267), .B1(n_1268), .B2(n_1271), .C(n_1273), .Y(n_1263) );
INVx2_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
OAI22xp33_ASAP7_75t_L g1338 ( .A1(n_1267), .A2(n_1276), .B1(n_1339), .B2(n_1340), .Y(n_1338) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_1276), .A2(n_1277), .B1(n_1279), .B2(n_1280), .Y(n_1275) );
INVx6_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
OAI22xp5_ASAP7_75t_L g1341 ( .A1(n_1279), .A2(n_1283), .B1(n_1325), .B2(n_1342), .Y(n_1341) );
INVx4_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1284), .Y(n_1282) );
CKINVDCx8_ASAP7_75t_R g1285 ( .A(n_1286), .Y(n_1285) );
INVx2_ASAP7_75t_SL g1288 ( .A(n_1289), .Y(n_1288) );
AND2x4_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1293), .Y(n_1289) );
INVx3_ASAP7_75t_L g1316 ( .A(n_1291), .Y(n_1316) );
INVx2_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
NOR3xp33_ASAP7_75t_SL g1296 ( .A(n_1297), .B(n_1311), .C(n_1323), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1306), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1300), .B1(n_1304), .B2(n_1305), .Y(n_1298) );
BUFx2_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_1307), .A2(n_1308), .B1(n_1309), .B2(n_1310), .Y(n_1306) );
HB1xp67_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
NAND2x1_ASAP7_75t_SL g1313 ( .A(n_1314), .B(n_1316), .Y(n_1313) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
NAND2x1p5_ASAP7_75t_L g1318 ( .A(n_1316), .B(n_1319), .Y(n_1318) );
BUFx4f_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
BUFx3_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_1325), .A2(n_1327), .B1(n_1328), .B2(n_1329), .Y(n_1324) );
BUFx2_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
OAI22xp33_ASAP7_75t_L g1330 ( .A1(n_1331), .A2(n_1334), .B1(n_1335), .B2(n_1336), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
INVx2_ASAP7_75t_SL g1339 ( .A(n_1332), .Y(n_1339) );
INVx2_ASAP7_75t_SL g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
BUFx2_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1347), .Y(n_1395) );
HB1xp67_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1382), .Y(n_1370) );
BUFx2_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
INVx2_ASAP7_75t_SL g1376 ( .A(n_1377), .Y(n_1376) );
INVx2_ASAP7_75t_L g1381 ( .A(n_1377), .Y(n_1381) );
INVx2_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
CKINVDCx5p33_ASAP7_75t_R g1398 ( .A(n_1399), .Y(n_1398) );
endmodule