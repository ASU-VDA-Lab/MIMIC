module fake_netlist_5_2549_n_1147 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_211, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_1147);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1147;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_523;
wire n_268;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_947;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_1145;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_1016;
wire n_546;
wire n_856;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1096;
wire n_1095;
wire n_234;
wire n_343;
wire n_379;
wire n_428;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_1020;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_681;
wire n_584;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_866;
wire n_573;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_1058;
wire n_874;
wire n_465;
wire n_846;
wire n_358;
wire n_838;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_832;
wire n_695;
wire n_795;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1072;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_996;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_491;
wire n_272;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_811;
wire n_952;
wire n_766;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_1032;
wire n_360;
wire n_594;
wire n_890;
wire n_872;
wire n_1056;
wire n_764;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_167),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_39),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_68),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_30),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_123),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_153),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_91),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_78),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_187),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_50),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_172),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_16),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_104),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_184),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_72),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_108),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_17),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_154),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_131),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_133),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_6),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_7),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_74),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_67),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

BUFx8_ASAP7_75t_SL g242 ( 
.A(n_19),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_95),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_22),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_47),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_31),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_111),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_191),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_141),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_45),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_17),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_25),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_9),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_57),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_92),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_59),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_158),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_157),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_97),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_103),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_166),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_42),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_150),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_71),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_203),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_26),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_136),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_145),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_15),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_7),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_143),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_121),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_194),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_1),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_117),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_94),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_23),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_181),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_149),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_22),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_101),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_242),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_242),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_255),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_238),
.Y(n_293)
);

INVxp33_ASAP7_75t_SL g294 ( 
.A(n_214),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_216),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_212),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_226),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_226),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_236),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_232),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_220),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_239),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_244),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_216),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_220),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_221),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_241),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_246),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_270),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_254),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_227),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_227),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_234),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_257),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_273),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_260),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_263),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_234),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_254),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_245),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_267),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_277),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_229),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_302),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_302),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_317),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_306),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_319),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_301),
.B(n_231),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

AOI22x1_ASAP7_75t_SL g355 ( 
.A1(n_330),
.A2(n_256),
.B1(n_245),
.B2(n_281),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_298),
.B(n_304),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_285),
.Y(n_359)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_306),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_327),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_329),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_294),
.B(n_247),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_297),
.B(n_213),
.Y(n_364)
);

BUFx8_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_306),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_294),
.B(n_265),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_286),
.B(n_222),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_305),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_307),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_320),
.B(n_215),
.Y(n_376)
);

NAND2x1_ASAP7_75t_L g377 ( 
.A(n_323),
.B(n_324),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_325),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

OA21x2_ASAP7_75t_L g380 ( 
.A1(n_332),
.A2(n_284),
.B(n_218),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_289),
.A2(n_256),
.B1(n_282),
.B2(n_280),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_290),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_308),
.B(n_222),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_299),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_326),
.A2(n_283),
.B1(n_279),
.B2(n_275),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_310),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_334),
.A2(n_248),
.B(n_219),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_382),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_372),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_378),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_308),
.Y(n_393)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_372),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_345),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_388),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_378),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_345),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_347),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_335),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_335),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_365),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_365),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_388),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_368),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_365),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_322),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_384),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

BUFx6f_ASAP7_75t_SL g415 ( 
.A(n_384),
.Y(n_415)
);

BUFx10_ASAP7_75t_L g416 ( 
.A(n_383),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_369),
.Y(n_417)
);

NAND2xp33_ASAP7_75t_SL g418 ( 
.A(n_384),
.B(n_321),
.Y(n_418)
);

NOR2x1p5_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_287),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_355),
.B(n_330),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_384),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_377),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_L g423 ( 
.A(n_381),
.B(n_353),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_385),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_345),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_355),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_370),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_364),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_373),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_R g431 ( 
.A(n_380),
.B(n_321),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_386),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_349),
.B(n_322),
.Y(n_433)
);

NAND2xp33_ASAP7_75t_R g434 ( 
.A(n_380),
.B(n_288),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_359),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_385),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_370),
.B(n_336),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_338),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_338),
.Y(n_439)
);

INVxp33_ASAP7_75t_L g440 ( 
.A(n_357),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_349),
.B(n_217),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_344),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_344),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_357),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_345),
.Y(n_445)
);

AO21x2_ASAP7_75t_L g446 ( 
.A1(n_389),
.A2(n_225),
.B(n_223),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_357),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_346),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_373),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_373),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_373),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_380),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_373),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_379),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_R g455 ( 
.A(n_374),
.B(n_288),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_379),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_379),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_379),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_374),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_374),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_375),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_375),
.B(n_293),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_349),
.B(n_228),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_437),
.B(n_380),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_413),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_392),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_398),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_422),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_336),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_406),
.Y(n_472)
);

INVxp33_ASAP7_75t_SL g473 ( 
.A(n_391),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_425),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_417),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_400),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_437),
.B(n_463),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_395),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_437),
.B(n_342),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_428),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_421),
.B(n_389),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_442),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_402),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_436),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_405),
.B(n_233),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_394),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_409),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_442),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_438),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_410),
.B(n_235),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_402),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_437),
.B(n_342),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_439),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_418),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_414),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_464),
.B(n_371),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_423),
.B(n_341),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_424),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_428),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_444),
.B(n_371),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_443),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_433),
.B(n_343),
.Y(n_507)
);

BUFx4f_ASAP7_75t_L g508 ( 
.A(n_430),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_457),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_457),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_464),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_460),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_461),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_435),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_414),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_452),
.A2(n_248),
.B1(n_350),
.B2(n_348),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g517 ( 
.A(n_393),
.B(n_343),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_393),
.B(n_243),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_462),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_440),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_414),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_447),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_429),
.B(n_339),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_396),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_451),
.B(n_348),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_450),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_399),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_419),
.B(n_337),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_453),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_426),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_456),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_397),
.B(n_337),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_445),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_448),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_415),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_412),
.B(n_295),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_412),
.B(n_295),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_454),
.B(n_340),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_415),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_458),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_432),
.B(n_340),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_459),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_441),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_416),
.B(n_249),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_431),
.A2(n_434),
.B1(n_446),
.B2(n_416),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_446),
.B(n_250),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_404),
.B(n_352),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_408),
.Y(n_551)
);

AO22x2_ASAP7_75t_L g552 ( 
.A1(n_537),
.A2(n_420),
.B1(n_316),
.B2(n_328),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_509),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_486),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_489),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_528),
.B(n_510),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_468),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_528),
.B(n_505),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_517),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_500),
.B(n_367),
.Y(n_560)
);

OR2x2_ASAP7_75t_SL g561 ( 
.A(n_542),
.B(n_309),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_489),
.Y(n_562)
);

NOR2x1p5_ASAP7_75t_L g563 ( 
.A(n_467),
.B(n_411),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_511),
.B(n_367),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_511),
.B(n_309),
.Y(n_565)
);

AO22x2_ASAP7_75t_L g566 ( 
.A1(n_538),
.A2(n_328),
.B1(n_316),
.B2(n_427),
.Y(n_566)
);

NAND3x1_ASAP7_75t_L g567 ( 
.A(n_518),
.B(n_403),
.C(n_401),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_485),
.B(n_480),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_518),
.B(n_258),
.C(n_252),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_470),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_545),
.B(n_523),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_469),
.Y(n_572)
);

AO22x2_ASAP7_75t_L g573 ( 
.A1(n_503),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_480),
.B(n_367),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_475),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_523),
.B(n_361),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_472),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_505),
.B(n_352),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

NAND2x1p5_ASAP7_75t_L g580 ( 
.A(n_467),
.B(n_358),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_533),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_470),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_482),
.Y(n_583)
);

BUFx6f_ASAP7_75t_SL g584 ( 
.A(n_497),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_488),
.B(n_493),
.Y(n_585)
);

NAND2x1p5_ASAP7_75t_L g586 ( 
.A(n_487),
.B(n_358),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_549),
.A2(n_517),
.B1(n_516),
.B2(n_474),
.Y(n_587)
);

OAI221xp5_ASAP7_75t_L g588 ( 
.A1(n_516),
.A2(n_520),
.B1(n_488),
.B2(n_493),
.C(n_491),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_525),
.B(n_346),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_474),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_524),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_526),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_476),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_525),
.B(n_346),
.Y(n_594)
);

OAI221xp5_ASAP7_75t_L g595 ( 
.A1(n_483),
.A2(n_266),
.B1(n_268),
.B2(n_259),
.C(n_269),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_502),
.B(n_350),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_524),
.Y(n_597)
);

OR2x2_ASAP7_75t_SL g598 ( 
.A(n_551),
.B(n_248),
.Y(n_598)
);

OAI221xp5_ASAP7_75t_L g599 ( 
.A1(n_548),
.A2(n_512),
.B1(n_519),
.B2(n_513),
.C(n_543),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_549),
.A2(n_346),
.B1(n_362),
.B2(n_356),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_476),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_530),
.Y(n_602)
);

INVx3_ASAP7_75t_R g603 ( 
.A(n_490),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_539),
.B(n_346),
.Y(n_604)
);

BUFx8_ASAP7_75t_L g605 ( 
.A(n_506),
.Y(n_605)
);

NAND3x1_ASAP7_75t_L g606 ( 
.A(n_536),
.B(n_0),
.C(n_2),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_517),
.A2(n_264),
.B1(n_271),
.B2(n_272),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_514),
.B(n_3),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_532),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_534),
.Y(n_610)
);

BUFx8_ASAP7_75t_L g611 ( 
.A(n_522),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_535),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_486),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_477),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_546),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_539),
.B(n_351),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_531),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_477),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_565),
.B(n_546),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_585),
.B(n_487),
.Y(n_621)
);

OAI321xp33_ASAP7_75t_L g622 ( 
.A1(n_588),
.A2(n_547),
.A3(n_498),
.B1(n_540),
.B2(n_481),
.C(n_501),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_571),
.B(n_529),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_616),
.B(n_473),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_554),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_576),
.B(n_564),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_589),
.A2(n_466),
.B(n_495),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_615),
.B(n_529),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_594),
.A2(n_466),
.B(n_495),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_560),
.A2(n_495),
.B(n_544),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_SL g631 ( 
.A1(n_619),
.A2(n_481),
.B(n_501),
.C(n_479),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_557),
.B(n_572),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_559),
.A2(n_544),
.B(n_479),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_559),
.A2(n_544),
.B(n_496),
.Y(n_634)
);

AOI21x1_ASAP7_75t_L g635 ( 
.A1(n_604),
.A2(n_496),
.B(n_471),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_558),
.B(n_541),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_575),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_554),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_553),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_570),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_599),
.A2(n_517),
.B1(n_507),
.B2(n_541),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_574),
.B(n_517),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_592),
.B(n_507),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_554),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_587),
.A2(n_471),
.B(n_508),
.C(n_550),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_570),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_558),
.B(n_556),
.Y(n_647)
);

BUFx12f_ASAP7_75t_L g648 ( 
.A(n_605),
.Y(n_648)
);

A2O1A1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_577),
.A2(n_508),
.B(n_550),
.C(n_484),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_559),
.A2(n_521),
.B1(n_478),
.B2(n_515),
.Y(n_650)
);

NAND2x1p5_ASAP7_75t_L g651 ( 
.A(n_601),
.B(n_521),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_609),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_556),
.A2(n_507),
.B1(n_527),
.B2(n_504),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_582),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_590),
.A2(n_499),
.B(n_494),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_568),
.B(n_527),
.Y(n_656)
);

NOR2x1_ASAP7_75t_L g657 ( 
.A(n_569),
.B(n_527),
.Y(n_657)
);

AOI21x1_ASAP7_75t_L g658 ( 
.A1(n_610),
.A2(n_354),
.B(n_351),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_555),
.B(n_507),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_600),
.A2(n_341),
.B(n_356),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_562),
.B(n_507),
.Y(n_661)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_583),
.A2(n_613),
.B(n_617),
.C(n_578),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_617),
.A2(n_614),
.B(n_579),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_581),
.B(n_3),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_578),
.B(n_354),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_602),
.A2(n_366),
.B(n_360),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_593),
.B(n_4),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_596),
.B(n_366),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_579),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_612),
.B(n_4),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_579),
.A2(n_341),
.B(n_356),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_614),
.A2(n_362),
.B(n_356),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_561),
.B(n_5),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_618),
.A2(n_360),
.B(n_356),
.Y(n_674)
);

BUFx4f_ASAP7_75t_L g675 ( 
.A(n_580),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_596),
.B(n_362),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_591),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_614),
.A2(n_362),
.B(n_360),
.Y(n_678)
);

OA22x2_ASAP7_75t_L g679 ( 
.A1(n_566),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_679)
);

O2A1O1Ixp5_ASAP7_75t_L g680 ( 
.A1(n_597),
.A2(n_109),
.B(n_210),
.C(n_207),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_595),
.B(n_8),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_586),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_607),
.B(n_362),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_608),
.A2(n_360),
.B(n_33),
.Y(n_684)
);

BUFx4f_ASAP7_75t_L g685 ( 
.A(n_603),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_567),
.B(n_360),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_626),
.A2(n_629),
.B(n_627),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_SL g688 ( 
.A1(n_681),
.A2(n_598),
.B(n_552),
.C(n_566),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_621),
.B(n_623),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_637),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_620),
.B(n_552),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_645),
.A2(n_563),
.B(n_606),
.C(n_573),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_632),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_652),
.Y(n_694)
);

AO32x1_ASAP7_75t_L g695 ( 
.A1(n_650),
.A2(n_573),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_695)
);

O2A1O1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_673),
.A2(n_662),
.B(n_628),
.C(n_664),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_647),
.B(n_9),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_631),
.A2(n_634),
.B(n_633),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_624),
.B(n_584),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_675),
.B(n_605),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_644),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_639),
.B(n_611),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_668),
.B(n_665),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_647),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_675),
.B(n_611),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_SL g706 ( 
.A1(n_659),
.A2(n_584),
.B(n_110),
.C(n_112),
.Y(n_706)
);

O2A1O1Ixp5_ASAP7_75t_L g707 ( 
.A1(n_661),
.A2(n_10),
.B(n_11),
.C(n_13),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_683),
.A2(n_34),
.B(n_32),
.Y(n_708)
);

O2A1O1Ixp5_ASAP7_75t_L g709 ( 
.A1(n_649),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_630),
.A2(n_36),
.B(n_35),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_682),
.B(n_14),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_668),
.B(n_16),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_651),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_656),
.B(n_18),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_644),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_640),
.Y(n_716)
);

NOR3xp33_ASAP7_75t_SL g717 ( 
.A(n_667),
.B(n_670),
.C(n_636),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_685),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_685),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_622),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_679),
.B(n_20),
.Y(n_721)
);

AO32x1_ASAP7_75t_L g722 ( 
.A1(n_646),
.A2(n_21),
.A3(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_677),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_654),
.B(n_682),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_676),
.B(n_642),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_641),
.A2(n_38),
.B(n_37),
.Y(n_726)
);

O2A1O1Ixp5_ASAP7_75t_L g727 ( 
.A1(n_684),
.A2(n_21),
.B(n_24),
.C(n_26),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_663),
.B(n_27),
.Y(n_728)
);

A2O1A1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_643),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_648),
.B(n_40),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_SL g731 ( 
.A1(n_682),
.A2(n_638),
.B1(n_653),
.B2(n_657),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_644),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_625),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_638),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_625),
.B(n_206),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_680),
.A2(n_686),
.B(n_674),
.C(n_666),
.Y(n_736)
);

O2A1O1Ixp5_ASAP7_75t_L g737 ( 
.A1(n_635),
.A2(n_28),
.B(n_29),
.C(n_41),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_658),
.A2(n_43),
.B(n_44),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_669),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_669),
.B(n_205),
.Y(n_740)
);

A2O1A1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_655),
.A2(n_48),
.B(n_49),
.C(n_51),
.Y(n_741)
);

OAI21xp33_ASAP7_75t_L g742 ( 
.A1(n_660),
.A2(n_52),
.B(n_53),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_678),
.B(n_54),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_672),
.Y(n_744)
);

AND2x2_ASAP7_75t_SL g745 ( 
.A(n_671),
.B(n_55),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_620),
.B(n_56),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_637),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_685),
.B(n_58),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_644),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_621),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_721),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_751)
);

INVx5_ASAP7_75t_L g752 ( 
.A(n_701),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_701),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_715),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_719),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_739),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_718),
.Y(n_757)
);

NAND2x1_ASAP7_75t_L g758 ( 
.A(n_743),
.B(n_66),
.Y(n_758)
);

INVx6_ASAP7_75t_L g759 ( 
.A(n_734),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_732),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_694),
.Y(n_761)
);

OR2x6_ASAP7_75t_L g762 ( 
.A(n_731),
.B(n_69),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_715),
.Y(n_763)
);

INVx8_ASAP7_75t_L g764 ( 
.A(n_749),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_735),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_734),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_749),
.Y(n_767)
);

OR2x6_ASAP7_75t_L g768 ( 
.A(n_743),
.B(n_70),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_690),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_735),
.Y(n_770)
);

BUFx2_ASAP7_75t_SL g771 ( 
.A(n_700),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_704),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_702),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_747),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_697),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_705),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_740),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_716),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_713),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_733),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_725),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_693),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_689),
.B(n_73),
.Y(n_783)
);

BUFx2_ASAP7_75t_R g784 ( 
.A(n_691),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_703),
.Y(n_785)
);

BUFx2_ASAP7_75t_R g786 ( 
.A(n_711),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_699),
.Y(n_787)
);

BUFx2_ASAP7_75t_SL g788 ( 
.A(n_746),
.Y(n_788)
);

BUFx8_ASAP7_75t_SL g789 ( 
.A(n_730),
.Y(n_789)
);

BUFx10_ASAP7_75t_L g790 ( 
.A(n_724),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_723),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_712),
.Y(n_792)
);

BUFx2_ASAP7_75t_SL g793 ( 
.A(n_744),
.Y(n_793)
);

NAND2x1p5_ASAP7_75t_L g794 ( 
.A(n_745),
.B(n_75),
.Y(n_794)
);

INVx6_ASAP7_75t_L g795 ( 
.A(n_730),
.Y(n_795)
);

INVx8_ASAP7_75t_L g796 ( 
.A(n_748),
.Y(n_796)
);

BUFx10_ASAP7_75t_L g797 ( 
.A(n_717),
.Y(n_797)
);

INVx3_ASAP7_75t_SL g798 ( 
.A(n_688),
.Y(n_798)
);

AO21x2_ASAP7_75t_L g799 ( 
.A1(n_698),
.A2(n_687),
.B(n_736),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_728),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_738),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_714),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_692),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_696),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_708),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_710),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_706),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_741),
.Y(n_808)
);

INVx6_ASAP7_75t_L g809 ( 
.A(n_729),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_737),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_709),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_722),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_722),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_707),
.B(n_76),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_695),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_750),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_695),
.Y(n_817)
);

INVx6_ASAP7_75t_SL g818 ( 
.A(n_727),
.Y(n_818)
);

CKINVDCx8_ASAP7_75t_R g819 ( 
.A(n_720),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_726),
.B(n_77),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_742),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_769),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_769),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_774),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_781),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_801),
.A2(n_79),
.B(n_80),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_781),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_801),
.A2(n_81),
.B(n_82),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_782),
.Y(n_829)
);

NAND3xp33_ASAP7_75t_L g830 ( 
.A(n_819),
.B(n_83),
.C(n_84),
.Y(n_830)
);

OAI21x1_ASAP7_75t_L g831 ( 
.A1(n_810),
.A2(n_85),
.B(n_86),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_755),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_777),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_804),
.A2(n_809),
.B1(n_803),
.B2(n_797),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_785),
.B(n_87),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_760),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_759),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_785),
.B(n_88),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_752),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_777),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_821),
.A2(n_89),
.B(n_90),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_792),
.B(n_93),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_816),
.A2(n_96),
.B(n_98),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_802),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_844)
);

NAND3xp33_ASAP7_75t_SL g845 ( 
.A(n_805),
.B(n_105),
.C(n_106),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_800),
.B(n_107),
.Y(n_846)
);

OAI21x1_ASAP7_75t_L g847 ( 
.A1(n_816),
.A2(n_113),
.B(n_114),
.Y(n_847)
);

OAI21x1_ASAP7_75t_L g848 ( 
.A1(n_821),
.A2(n_115),
.B(n_116),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_809),
.A2(n_204),
.B1(n_118),
.B2(n_120),
.Y(n_849)
);

OAI21x1_ASAP7_75t_L g850 ( 
.A1(n_814),
.A2(n_782),
.B(n_758),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_778),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_785),
.B(n_792),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_812),
.A2(n_122),
.B(n_124),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_761),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_SL g855 ( 
.A1(n_783),
.A2(n_806),
.B(n_817),
.C(n_815),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_800),
.B(n_125),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_759),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_780),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_777),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_770),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_791),
.B(n_126),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_793),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_797),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_863)
);

AO21x2_ASAP7_75t_L g864 ( 
.A1(n_799),
.A2(n_130),
.B(n_132),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_786),
.B(n_134),
.Y(n_865)
);

AOI211xp5_ASAP7_75t_L g866 ( 
.A1(n_798),
.A2(n_135),
.B(n_137),
.C(n_138),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_812),
.A2(n_139),
.B(n_140),
.Y(n_867)
);

NOR2x1_ASAP7_75t_SL g868 ( 
.A(n_762),
.B(n_142),
.Y(n_868)
);

AOI221xp5_ASAP7_75t_L g869 ( 
.A1(n_811),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.C(n_148),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_SL g870 ( 
.A1(n_783),
.A2(n_817),
.B(n_815),
.C(n_813),
.Y(n_870)
);

AO21x2_ASAP7_75t_L g871 ( 
.A1(n_813),
.A2(n_820),
.B(n_818),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_794),
.A2(n_151),
.B(n_152),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_794),
.A2(n_155),
.B(n_156),
.Y(n_873)
);

OA21x2_ASAP7_75t_L g874 ( 
.A1(n_818),
.A2(n_159),
.B(n_161),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_786),
.B(n_162),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_800),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_772),
.B(n_163),
.Y(n_877)
);

AO21x2_ASAP7_75t_L g878 ( 
.A1(n_807),
.A2(n_164),
.B(n_165),
.Y(n_878)
);

OA21x2_ASAP7_75t_L g879 ( 
.A1(n_807),
.A2(n_168),
.B(n_169),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_765),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_762),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_822),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_862),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_850),
.B(n_762),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_829),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_832),
.B(n_787),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_823),
.Y(n_887)
);

BUFx4f_ASAP7_75t_SL g888 ( 
.A(n_832),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_860),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_823),
.B(n_751),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_825),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_827),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_858),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_824),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_824),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_SL g896 ( 
.A1(n_868),
.A2(n_796),
.B1(n_808),
.B2(n_795),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_852),
.B(n_751),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_871),
.Y(n_898)
);

NAND2x1_ASAP7_75t_L g899 ( 
.A(n_874),
.B(n_795),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_851),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_829),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_854),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_870),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_880),
.Y(n_904)
);

AO21x1_ASAP7_75t_L g905 ( 
.A1(n_866),
.A2(n_808),
.B(n_770),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_880),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_881),
.A2(n_796),
.B1(n_768),
.B2(n_775),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_SL g908 ( 
.A(n_830),
.B(n_771),
.Y(n_908)
);

AOI21x1_ASAP7_75t_L g909 ( 
.A1(n_841),
.A2(n_768),
.B(n_776),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_876),
.B(n_768),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_871),
.Y(n_911)
);

CKINVDCx11_ASAP7_75t_R g912 ( 
.A(n_833),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_836),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_850),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_833),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_855),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_855),
.Y(n_917)
);

AO21x2_ASAP7_75t_L g918 ( 
.A1(n_864),
.A2(n_807),
.B(n_796),
.Y(n_918)
);

AOI31xp33_ASAP7_75t_L g919 ( 
.A1(n_881),
.A2(n_772),
.A3(n_789),
.B(n_784),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_853),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_831),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_834),
.A2(n_784),
.B1(n_788),
.B2(n_773),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_833),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_833),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_882),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_888),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_912),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_R g928 ( 
.A(n_910),
.B(n_874),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_SL g929 ( 
.A(n_905),
.B(n_834),
.C(n_865),
.Y(n_929)
);

NAND2xp33_ASAP7_75t_SL g930 ( 
.A(n_908),
.B(n_839),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_893),
.B(n_840),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_883),
.B(n_859),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_919),
.A2(n_875),
.B(n_865),
.C(n_844),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_907),
.A2(n_875),
.B1(n_905),
.B2(n_922),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_913),
.B(n_840),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_894),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_891),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_894),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_883),
.B(n_859),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_923),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_887),
.B(n_842),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_896),
.B(n_860),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_924),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_897),
.B(n_859),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_895),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_SL g946 ( 
.A1(n_890),
.A2(n_874),
.B1(n_879),
.B2(n_864),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_912),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_886),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_R g949 ( 
.A(n_910),
.B(n_879),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_892),
.Y(n_950)
);

BUFx5_ASAP7_75t_L g951 ( 
.A(n_920),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_904),
.B(n_859),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_SL g953 ( 
.A1(n_890),
.A2(n_863),
.B(n_849),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_SL g954 ( 
.A(n_908),
.B(n_861),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_897),
.B(n_773),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_904),
.B(n_867),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_903),
.Y(n_957)
);

CKINVDCx11_ASAP7_75t_R g958 ( 
.A(n_923),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_904),
.B(n_906),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_900),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_959),
.B(n_898),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_959),
.B(n_911),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_925),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_936),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_943),
.B(n_911),
.Y(n_965)
);

INVx8_ASAP7_75t_L g966 ( 
.A(n_927),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_938),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_945),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_944),
.B(n_884),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_937),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_950),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_931),
.B(n_902),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_960),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_957),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_939),
.B(n_884),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_935),
.B(n_884),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_941),
.Y(n_977)
);

NOR2x1p5_ASAP7_75t_L g978 ( 
.A(n_929),
.B(n_899),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_952),
.B(n_884),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_955),
.B(n_956),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_952),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_956),
.B(n_914),
.Y(n_982)
);

AOI222xp33_ASAP7_75t_L g983 ( 
.A1(n_953),
.A2(n_869),
.B1(n_863),
.B2(n_845),
.C1(n_916),
.C2(n_917),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_932),
.B(n_885),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_951),
.Y(n_985)
);

NAND2x1_ASAP7_75t_L g986 ( 
.A(n_979),
.B(n_932),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_969),
.B(n_947),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_983),
.A2(n_953),
.B(n_930),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_963),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_970),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_965),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_978),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_979),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_966),
.A2(n_933),
.B(n_934),
.C(n_954),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_971),
.Y(n_995)
);

OAI211xp5_ASAP7_75t_L g996 ( 
.A1(n_974),
.A2(n_934),
.B(n_946),
.C(n_942),
.Y(n_996)
);

NAND3xp33_ASAP7_75t_L g997 ( 
.A(n_965),
.B(n_949),
.C(n_928),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_973),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_964),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_966),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_966),
.B(n_926),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_964),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_993),
.B(n_961),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_992),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_999),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_993),
.B(n_992),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_991),
.B(n_961),
.Y(n_1007)
);

OAI221xp5_ASAP7_75t_L g1008 ( 
.A1(n_994),
.A2(n_948),
.B1(n_984),
.B2(n_972),
.C(n_977),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_989),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_991),
.B(n_986),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_990),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_995),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_997),
.B(n_981),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_987),
.B(n_962),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_998),
.B(n_962),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_998),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_1014),
.B(n_1000),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_1004),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_L g1019 ( 
.A(n_1010),
.B(n_996),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_1006),
.B(n_988),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_1010),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_1013),
.B(n_1002),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_1006),
.B(n_979),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1006),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1009),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1011),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_1019),
.A2(n_1008),
.B1(n_1016),
.B2(n_1007),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_1020),
.B(n_1018),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1023),
.B(n_1014),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1025),
.Y(n_1030)
);

INVxp67_ASAP7_75t_L g1031 ( 
.A(n_1020),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_1022),
.B(n_1012),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_1023),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1029),
.B(n_1017),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1032),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_1031),
.B(n_966),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_1033),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1028),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1030),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1027),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_1027),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1029),
.B(n_1023),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1031),
.B(n_1024),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_1038),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1043),
.B(n_1024),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_1037),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1042),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1034),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1038),
.B(n_1036),
.Y(n_1049)
);

CKINVDCx16_ASAP7_75t_R g1050 ( 
.A(n_1036),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1037),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_1035),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1046),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1047),
.A2(n_1041),
.B1(n_1040),
.B2(n_1021),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1051),
.Y(n_1055)
);

AOI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_1044),
.A2(n_1039),
.B1(n_1021),
.B2(n_1026),
.C(n_1005),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1050),
.A2(n_1015),
.B1(n_1003),
.B2(n_1007),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1051),
.Y(n_1058)
);

OAI21xp33_ASAP7_75t_L g1059 ( 
.A1(n_1049),
.A2(n_1015),
.B(n_1003),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1048),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1054),
.B(n_1052),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1053),
.B(n_1058),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1055),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1060),
.B(n_1045),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1059),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1062),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1061),
.B(n_1057),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1064),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1063),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1065),
.A2(n_1056),
.B1(n_1005),
.B2(n_1001),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1063),
.Y(n_1071)
);

OAI321xp33_ASAP7_75t_L g1072 ( 
.A1(n_1067),
.A2(n_837),
.A3(n_857),
.B1(n_849),
.B2(n_846),
.C(n_877),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1070),
.B(n_982),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_1068),
.B(n_756),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1071),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1069),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1066),
.B(n_982),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_1075),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_1076),
.A2(n_757),
.B(n_873),
.C(n_872),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_1074),
.A2(n_878),
.B(n_846),
.C(n_879),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1073),
.A2(n_856),
.B(n_773),
.Y(n_1081)
);

NAND4xp25_ASAP7_75t_SL g1082 ( 
.A(n_1077),
.B(n_1072),
.C(n_969),
.D(n_976),
.Y(n_1082)
);

AOI22x1_ASAP7_75t_L g1083 ( 
.A1(n_1078),
.A2(n_766),
.B1(n_763),
.B2(n_767),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_SL g1084 ( 
.A1(n_1081),
.A2(n_838),
.B(n_835),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_1080),
.A2(n_1079),
.B(n_1082),
.C(n_878),
.Y(n_1085)
);

AOI211xp5_ASAP7_75t_L g1086 ( 
.A1(n_1078),
.A2(n_753),
.B(n_754),
.C(n_767),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1078),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_1078),
.Y(n_1088)
);

AOI222xp33_ASAP7_75t_L g1089 ( 
.A1(n_1078),
.A2(n_779),
.B1(n_873),
.B2(n_872),
.C1(n_790),
.C2(n_985),
.Y(n_1089)
);

NAND2x1p5_ASAP7_75t_SL g1090 ( 
.A(n_1078),
.B(n_766),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1087),
.Y(n_1091)
);

AOI211x1_ASAP7_75t_L g1092 ( 
.A1(n_1090),
.A2(n_909),
.B(n_976),
.C(n_980),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_1088),
.B(n_1086),
.C(n_1083),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_1085),
.B(n_1089),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_1084),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1088),
.A2(n_764),
.B(n_752),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1088),
.B(n_980),
.Y(n_1097)
);

AOI322xp5_ASAP7_75t_L g1098 ( 
.A1(n_1088),
.A2(n_975),
.A3(n_910),
.B1(n_915),
.B2(n_752),
.C1(n_764),
.C2(n_940),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1088),
.A2(n_790),
.B1(n_764),
.B2(n_767),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1087),
.Y(n_1100)
);

OAI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_1091),
.A2(n_753),
.B(n_754),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_L g1102 ( 
.A(n_1100),
.B(n_843),
.C(n_847),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_SL g1103 ( 
.A1(n_1096),
.A2(n_174),
.B(n_175),
.C(n_176),
.Y(n_1103)
);

NAND2x1p5_ASAP7_75t_L g1104 ( 
.A(n_1097),
.B(n_753),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1095),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1099),
.B(n_975),
.Y(n_1106)
);

AND3x2_ASAP7_75t_L g1107 ( 
.A(n_1093),
.B(n_177),
.C(n_178),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_L g1108 ( 
.A(n_1094),
.B(n_179),
.Y(n_1108)
);

NOR2x1_ASAP7_75t_L g1109 ( 
.A(n_1092),
.B(n_754),
.Y(n_1109)
);

NAND5xp2_ASAP7_75t_L g1110 ( 
.A(n_1098),
.B(n_909),
.C(n_183),
.D(n_185),
.E(n_186),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_1097),
.B(n_940),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_1097),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_SL g1113 ( 
.A(n_1093),
.B(n_889),
.C(n_967),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1112),
.Y(n_1114)
);

CKINVDCx16_ASAP7_75t_R g1115 ( 
.A(n_1105),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1108),
.A2(n_843),
.B(n_826),
.Y(n_1116)
);

CKINVDCx16_ASAP7_75t_R g1117 ( 
.A(n_1113),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_1107),
.Y(n_1118)
);

CKINVDCx14_ASAP7_75t_R g1119 ( 
.A(n_1111),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_1104),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1103),
.A2(n_826),
.B(n_828),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1114),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1115),
.Y(n_1123)
);

XNOR2xp5_ASAP7_75t_L g1124 ( 
.A(n_1118),
.B(n_1109),
.Y(n_1124)
);

BUFx2_ASAP7_75t_SL g1125 ( 
.A(n_1120),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1119),
.B(n_1106),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1117),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1116),
.B(n_1101),
.Y(n_1128)
);

OR3x2_ASAP7_75t_L g1129 ( 
.A(n_1123),
.B(n_1110),
.C(n_1121),
.Y(n_1129)
);

OA21x2_ASAP7_75t_L g1130 ( 
.A1(n_1126),
.A2(n_1102),
.B(n_848),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1124),
.A2(n_828),
.B(n_831),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1129),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1132),
.A2(n_1127),
.B1(n_1122),
.B2(n_1125),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1133),
.A2(n_1128),
.B(n_1130),
.Y(n_1134)
);

XOR2xp5_ASAP7_75t_L g1135 ( 
.A(n_1134),
.B(n_182),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1134),
.A2(n_1131),
.B1(n_940),
.B2(n_923),
.Y(n_1136)
);

NAND5xp2_ASAP7_75t_L g1137 ( 
.A(n_1134),
.B(n_188),
.C(n_189),
.D(n_190),
.E(n_192),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1135),
.Y(n_1138)
);

AOI222xp33_ASAP7_75t_L g1139 ( 
.A1(n_1136),
.A2(n_958),
.B1(n_967),
.B2(n_968),
.C1(n_915),
.C2(n_923),
.Y(n_1139)
);

XNOR2xp5_ASAP7_75t_L g1140 ( 
.A(n_1137),
.B(n_195),
.Y(n_1140)
);

AOI322xp5_ASAP7_75t_L g1141 ( 
.A1(n_1138),
.A2(n_968),
.A3(n_923),
.B1(n_921),
.B2(n_914),
.C1(n_906),
.C2(n_901),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1140),
.A2(n_918),
.B1(n_951),
.B2(n_889),
.Y(n_1142)
);

OAI31xp33_ASAP7_75t_L g1143 ( 
.A1(n_1139),
.A2(n_196),
.A3(n_197),
.B(n_198),
.Y(n_1143)
);

AO21x2_ASAP7_75t_L g1144 ( 
.A1(n_1142),
.A2(n_199),
.B(n_200),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1143),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1145),
.A2(n_1141),
.B1(n_918),
.B2(n_951),
.Y(n_1146)
);

AOI211xp5_ASAP7_75t_L g1147 ( 
.A1(n_1146),
.A2(n_1144),
.B(n_201),
.C(n_202),
.Y(n_1147)
);


endmodule