module real_aes_16600_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_831, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_831;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g116 ( .A(n_0), .B(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_1), .A2(n_4), .B1(n_158), .B2(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_2), .A2(n_40), .B1(n_165), .B2(n_201), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_3), .A2(n_23), .B1(n_201), .B2(n_243), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_5), .A2(n_15), .B1(n_155), .B2(n_232), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_6), .A2(n_58), .B1(n_215), .B2(n_245), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_7), .A2(n_16), .B1(n_165), .B2(n_186), .Y(n_601) );
INVx1_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_9), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_10), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_11), .A2(n_17), .B1(n_214), .B2(n_217), .Y(n_213) );
BUFx2_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
OR2x2_ASAP7_75t_L g127 ( .A(n_12), .B(n_36), .Y(n_127) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_13), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_14), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_18), .A2(n_99), .B1(n_155), .B2(n_158), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_19), .A2(n_37), .B1(n_190), .B2(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_20), .B(n_156), .Y(n_187) );
OAI21x1_ASAP7_75t_L g173 ( .A1(n_21), .A2(n_54), .B(n_174), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_22), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_24), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_25), .B(n_162), .Y(n_521) );
INVx4_ASAP7_75t_R g569 ( .A(n_26), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_27), .A2(n_45), .B1(n_203), .B2(n_204), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_28), .A2(n_51), .B1(n_155), .B2(n_204), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_29), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_30), .B(n_190), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_31), .Y(n_266) );
INVx1_ASAP7_75t_L g500 ( .A(n_32), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_33), .B(n_201), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_SL g512 ( .A1(n_34), .A2(n_161), .B(n_165), .C(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_35), .A2(n_52), .B1(n_165), .B2(n_204), .Y(n_489) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_36), .Y(n_107) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_38), .A2(n_85), .B1(n_165), .B2(n_242), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_39), .A2(n_44), .B1(n_165), .B2(n_186), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_41), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_42), .A2(n_56), .B1(n_155), .B2(n_164), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_43), .A2(n_69), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_43), .Y(n_131) );
INVx1_ASAP7_75t_L g524 ( .A(n_46), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_47), .B(n_165), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_48), .Y(n_541) );
INVx2_ASAP7_75t_L g122 ( .A(n_49), .Y(n_122) );
INVx1_ASAP7_75t_L g111 ( .A(n_50), .Y(n_111) );
BUFx3_ASAP7_75t_L g125 ( .A(n_50), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_53), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_55), .A2(n_86), .B1(n_165), .B2(n_204), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_57), .A2(n_65), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_57), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_59), .A2(n_73), .B1(n_164), .B2(n_203), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_60), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_61), .A2(n_75), .B1(n_165), .B2(n_186), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_62), .A2(n_98), .B1(n_155), .B2(n_217), .Y(n_263) );
AND2x4_ASAP7_75t_L g151 ( .A(n_63), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g174 ( .A(n_64), .Y(n_174) );
INVx1_ASAP7_75t_L g806 ( .A(n_65), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_66), .A2(n_89), .B1(n_203), .B2(n_204), .Y(n_496) );
AO22x1_ASAP7_75t_L g558 ( .A1(n_67), .A2(n_74), .B1(n_229), .B2(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g152 ( .A(n_68), .Y(n_152) );
INVx1_ASAP7_75t_L g130 ( .A(n_69), .Y(n_130) );
AND2x2_ASAP7_75t_L g516 ( .A(n_70), .B(n_196), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_71), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_72), .B(n_245), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_76), .B(n_201), .Y(n_542) );
INVx2_ASAP7_75t_L g162 ( .A(n_77), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_78), .B(n_196), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_79), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_80), .A2(n_97), .B1(n_204), .B2(n_245), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_81), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_82), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_83), .B(n_172), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_84), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g827 ( .A(n_87), .Y(n_827) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_88), .B(n_196), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_90), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_91), .B(n_196), .Y(n_538) );
INVx1_ASAP7_75t_L g115 ( .A(n_92), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_92), .B(n_812), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g815 ( .A1(n_93), .A2(n_816), .B(n_823), .Y(n_815) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_94), .B(n_156), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_95), .A2(n_220), .B(n_245), .C(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g571 ( .A(n_96), .B(n_572), .Y(n_571) );
NAND2xp33_ASAP7_75t_L g546 ( .A(n_100), .B(n_191), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_118), .B(n_828), .Y(n_101) );
NOR2xp33_ASAP7_75t_SL g828 ( .A(n_102), .B(n_829), .Y(n_828) );
BUFx12f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x6_ASAP7_75t_SL g103 ( .A(n_104), .B(n_108), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
AND3x2_ASAP7_75t_L g826 ( .A(n_110), .B(n_114), .C(n_126), .Y(n_826) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g812 ( .A(n_111), .Y(n_812) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g137 ( .A(n_115), .Y(n_137) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_128), .B(n_802), .Y(n_118) );
BUFx12f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x6_ASAP7_75t_SL g120 ( .A(n_121), .B(n_123), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g814 ( .A(n_122), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_122), .B(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NOR2x1_ASAP7_75t_L g822 ( .A(n_125), .B(n_127), .Y(n_822) );
AND2x6_ASAP7_75t_SL g810 ( .A(n_126), .B(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
XNOR2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_132), .Y(n_128) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_138), .B1(n_478), .B2(n_479), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_136), .Y(n_478) );
BUFx8_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g821 ( .A(n_137), .B(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
XOR2xp5_ASAP7_75t_L g804 ( .A(n_139), .B(n_805), .Y(n_804) );
OR2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_381), .Y(n_139) );
NAND4xp25_ASAP7_75t_L g140 ( .A(n_141), .B(n_305), .C(n_336), .D(n_365), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_272), .Y(n_141) );
OAI322xp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_208), .A3(n_237), .B1(n_250), .B2(n_258), .C1(n_267), .C2(n_269), .Y(n_142) );
INVxp67_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_144), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_178), .Y(n_144) );
AND2x2_ASAP7_75t_L g302 ( .A(n_145), .B(n_303), .Y(n_302) );
INVx4_ASAP7_75t_L g338 ( .A(n_145), .Y(n_338) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g313 ( .A(n_146), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g316 ( .A(n_146), .B(n_210), .Y(n_316) );
AND2x2_ASAP7_75t_L g333 ( .A(n_146), .B(n_226), .Y(n_333) );
AND2x2_ASAP7_75t_L g431 ( .A(n_146), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g254 ( .A(n_147), .Y(n_254) );
AND2x4_ASAP7_75t_L g437 ( .A(n_147), .B(n_432), .Y(n_437) );
AO31x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_153), .A3(n_169), .B(n_175), .Y(n_147) );
AO31x2_ASAP7_75t_L g261 ( .A1(n_148), .A2(n_221), .A3(n_262), .B(n_265), .Y(n_261) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_149), .A2(n_564), .B(n_567), .Y(n_563) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AO31x2_ASAP7_75t_L g198 ( .A1(n_150), .A2(n_199), .A3(n_205), .B(n_206), .Y(n_198) );
AO31x2_ASAP7_75t_L g211 ( .A1(n_150), .A2(n_212), .A3(n_221), .B(n_223), .Y(n_211) );
AO31x2_ASAP7_75t_L g226 ( .A1(n_150), .A2(n_227), .A3(n_234), .B(n_235), .Y(n_226) );
AO31x2_ASAP7_75t_L g599 ( .A1(n_150), .A2(n_177), .A3(n_600), .B(n_603), .Y(n_599) );
BUFx10_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g194 ( .A(n_151), .Y(n_194) );
BUFx10_ASAP7_75t_L g491 ( .A(n_151), .Y(n_491) );
INVx1_ASAP7_75t_L g515 ( .A(n_151), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_160), .B1(n_163), .B2(n_166), .Y(n_153) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_156), .Y(n_559) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g159 ( .A(n_157), .Y(n_159) );
INVx3_ASAP7_75t_L g165 ( .A(n_157), .Y(n_165) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_157), .Y(n_191) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_157), .Y(n_201) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
INVx1_ASAP7_75t_L g216 ( .A(n_157), .Y(n_216) );
INVx1_ASAP7_75t_L g230 ( .A(n_157), .Y(n_230) );
INVx1_ASAP7_75t_L g233 ( .A(n_157), .Y(n_233) );
INVx2_ASAP7_75t_L g243 ( .A(n_157), .Y(n_243) );
INVx1_ASAP7_75t_L g245 ( .A(n_157), .Y(n_245) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_159), .B(n_509), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_160), .A2(n_189), .B(n_192), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_160), .A2(n_166), .B1(n_200), .B2(n_202), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_160), .A2(n_213), .B1(n_218), .B2(n_219), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_160), .A2(n_166), .B1(n_228), .B2(n_231), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_160), .A2(n_241), .B1(n_244), .B2(n_246), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_160), .A2(n_219), .B1(n_263), .B2(n_264), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_160), .A2(n_166), .B1(n_282), .B2(n_283), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_160), .A2(n_488), .B1(n_489), .B2(n_490), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_160), .A2(n_246), .B1(n_496), .B2(n_497), .Y(n_495) );
OAI22x1_ASAP7_75t_L g600 ( .A1(n_160), .A2(n_246), .B1(n_601), .B2(n_602), .Y(n_600) );
INVx6_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
O2A1O1Ixp5_ASAP7_75t_L g184 ( .A1(n_161), .A2(n_185), .B(n_186), .C(n_187), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_161), .A2(n_546), .B(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_161), .B(n_558), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g615 ( .A1(n_161), .A2(n_554), .B(n_558), .C(n_561), .Y(n_615) );
BUFx8_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g168 ( .A(n_162), .Y(n_168) );
INVx1_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
INVx1_ASAP7_75t_L g511 ( .A(n_162), .Y(n_511) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx4_ASAP7_75t_L g186 ( .A(n_165), .Y(n_186) );
INVx1_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g490 ( .A(n_167), .Y(n_490) );
BUFx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g544 ( .A(n_168), .Y(n_544) );
AO31x2_ASAP7_75t_L g280 ( .A1(n_169), .A2(n_247), .A3(n_281), .B(n_284), .Y(n_280) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_169), .A2(n_563), .B(n_571), .Y(n_562) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g223 ( .A(n_171), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_171), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g177 ( .A(n_172), .Y(n_177) );
INVx2_ASAP7_75t_L g222 ( .A(n_172), .Y(n_222) );
OAI21xp33_ASAP7_75t_L g561 ( .A1(n_172), .A2(n_515), .B(n_556), .Y(n_561) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_173), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_177), .B(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g442 ( .A(n_178), .B(n_343), .Y(n_442) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g271 ( .A(n_179), .Y(n_271) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_179), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_197), .Y(n_179) );
AND2x2_ASAP7_75t_L g259 ( .A(n_180), .B(n_198), .Y(n_259) );
INVx1_ASAP7_75t_L g300 ( .A(n_180), .Y(n_300) );
OAI21x1_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_183), .B(n_195), .Y(n_180) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_181), .A2(n_183), .B(n_195), .Y(n_295) );
INVx2_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
INVx4_ASAP7_75t_L g196 ( .A(n_182), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_182), .B(n_207), .Y(n_206) );
BUFx3_ASAP7_75t_L g234 ( .A(n_182), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_182), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_182), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g528 ( .A(n_182), .B(n_491), .Y(n_528) );
OAI21x1_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_188), .B(n_193), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_186), .A2(n_541), .B(n_542), .C(n_543), .Y(n_540) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g203 ( .A(n_191), .Y(n_203) );
OAI22xp33_ASAP7_75t_L g568 ( .A1(n_191), .A2(n_233), .B1(n_569), .B2(n_570), .Y(n_568) );
INVx2_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_SL g247 ( .A(n_194), .Y(n_247) );
INVx2_ASAP7_75t_L g205 ( .A(n_196), .Y(n_205) );
NOR2x1_ASAP7_75t_L g548 ( .A(n_196), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g291 ( .A(n_197), .Y(n_291) );
AND2x2_ASAP7_75t_L g355 ( .A(n_197), .B(n_294), .Y(n_355) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g309 ( .A(n_198), .Y(n_309) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_198), .Y(n_362) );
OR2x2_ASAP7_75t_L g433 ( .A(n_198), .B(n_239), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_201), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g498 ( .A(n_204), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_204), .B(n_523), .Y(n_522) );
AO31x2_ASAP7_75t_L g486 ( .A1(n_205), .A2(n_487), .A3(n_491), .B(n_492), .Y(n_486) );
NAND4xp25_ASAP7_75t_L g311 ( .A(n_208), .B(n_312), .C(n_315), .D(n_317), .Y(n_311) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g449 ( .A(n_209), .B(n_437), .Y(n_449) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_225), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_210), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g303 ( .A(n_210), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g323 ( .A(n_210), .Y(n_323) );
INVx1_ASAP7_75t_L g340 ( .A(n_210), .Y(n_340) );
INVx1_ASAP7_75t_L g348 ( .A(n_210), .Y(n_348) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_210), .Y(n_462) );
INVx4_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_211), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g380 ( .A(n_211), .B(n_280), .Y(n_380) );
AND2x2_ASAP7_75t_L g388 ( .A(n_211), .B(n_226), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_211), .B(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g453 ( .A(n_211), .Y(n_453) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_216), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g246 ( .A(n_220), .Y(n_246) );
AO31x2_ASAP7_75t_L g494 ( .A1(n_221), .A2(n_247), .A3(n_495), .B(n_499), .Y(n_494) );
AOI21x1_ASAP7_75t_L g503 ( .A1(n_221), .A2(n_504), .B(n_516), .Y(n_503) );
BUFx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_222), .B(n_493), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_222), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g572 ( .A(n_222), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_222), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g257 ( .A(n_226), .Y(n_257) );
OR2x2_ASAP7_75t_L g318 ( .A(n_226), .B(n_280), .Y(n_318) );
INVx2_ASAP7_75t_L g325 ( .A(n_226), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_226), .B(n_278), .Y(n_349) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_226), .Y(n_436) );
OAI21xp33_ASAP7_75t_SL g520 ( .A1(n_229), .A2(n_521), .B(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AO31x2_ASAP7_75t_L g239 ( .A1(n_234), .A2(n_240), .A3(n_247), .B(n_248), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_237), .B(n_408), .Y(n_407) );
BUFx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g260 ( .A(n_239), .B(n_261), .Y(n_260) );
BUFx2_ASAP7_75t_L g270 ( .A(n_239), .Y(n_270) );
INVx2_ASAP7_75t_L g288 ( .A(n_239), .Y(n_288) );
AND2x4_ASAP7_75t_L g320 ( .A(n_239), .B(n_292), .Y(n_320) );
OR2x2_ASAP7_75t_L g400 ( .A(n_239), .B(n_300), .Y(n_400) );
INVx2_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_243), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_246), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_255), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_252), .B(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g317 ( .A(n_252), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_252), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_253), .B(n_323), .Y(n_331) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g276 ( .A(n_254), .Y(n_276) );
OR2x2_ASAP7_75t_L g369 ( .A(n_254), .B(n_279), .Y(n_369) );
INVx1_ASAP7_75t_L g296 ( .A(n_255), .Y(n_296) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g268 ( .A(n_256), .Y(n_268) );
INVx1_ASAP7_75t_L g304 ( .A(n_257), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
OAI322xp33_ASAP7_75t_L g272 ( .A1(n_259), .A2(n_273), .A3(n_286), .B1(n_289), .B2(n_296), .C1(n_297), .C2(n_301), .Y(n_272) );
AND2x4_ASAP7_75t_L g319 ( .A(n_259), .B(n_320), .Y(n_319) );
AOI211xp5_ASAP7_75t_SL g350 ( .A1(n_259), .A2(n_351), .B(n_352), .C(n_356), .Y(n_350) );
AND2x2_ASAP7_75t_L g370 ( .A(n_259), .B(n_260), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_259), .B(n_287), .Y(n_376) );
AND2x4_ASAP7_75t_SL g298 ( .A(n_260), .B(n_299), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g389 ( .A(n_260), .B(n_316), .C(n_344), .Y(n_389) );
AND2x2_ASAP7_75t_L g420 ( .A(n_260), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g287 ( .A(n_261), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g292 ( .A(n_261), .Y(n_292) );
BUFx2_ASAP7_75t_L g360 ( .A(n_261), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_270), .B(n_294), .Y(n_293) );
NAND2x1_ASAP7_75t_L g334 ( .A(n_270), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g353 ( .A(n_270), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_271), .B(n_287), .Y(n_418) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g361 ( .A(n_276), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_280), .Y(n_314) );
AND2x4_ASAP7_75t_L g324 ( .A(n_280), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g411 ( .A(n_280), .Y(n_411) );
INVx2_ASAP7_75t_L g432 ( .A(n_280), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_286), .A2(n_445), .B1(n_447), .B2(n_448), .Y(n_444) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g356 ( .A(n_287), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g310 ( .A(n_288), .B(n_294), .Y(n_310) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g329 ( .A(n_290), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x4_ASAP7_75t_L g299 ( .A(n_291), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g421 ( .A(n_291), .Y(n_421) );
INVx2_ASAP7_75t_L g307 ( .A(n_292), .Y(n_307) );
AND2x2_ASAP7_75t_L g335 ( .A(n_292), .B(n_294), .Y(n_335) );
INVx3_ASAP7_75t_L g343 ( .A(n_292), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_292), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g328 ( .A(n_293), .Y(n_328) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_L g344 ( .A(n_295), .Y(n_344) );
OAI222xp33_ASAP7_75t_L g467 ( .A1(n_297), .A2(n_457), .B1(n_468), .B2(n_471), .C1(n_473), .C2(n_475), .Y(n_467) );
INVx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g408 ( .A(n_299), .Y(n_408) );
AND2x2_ASAP7_75t_L g472 ( .A(n_299), .B(n_342), .Y(n_472) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_302), .B(n_393), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_311), .B1(n_319), .B2(n_321), .C(n_326), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g394 ( .A(n_307), .Y(n_394) );
INVx2_ASAP7_75t_L g456 ( .A(n_308), .Y(n_456) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g357 ( .A(n_309), .Y(n_357) );
AND2x2_ASAP7_75t_L g393 ( .A(n_309), .B(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g359 ( .A(n_310), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g385 ( .A(n_310), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g474 ( .A(n_310), .Y(n_474) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g423 ( .A(n_314), .Y(n_423) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g446 ( .A(n_316), .B(n_324), .Y(n_446) );
AND2x2_ASAP7_75t_L g469 ( .A(n_316), .B(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g330 ( .A(n_318), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g465 ( .A(n_318), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_319), .A2(n_373), .B1(n_407), .B2(n_409), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_319), .A2(n_435), .B(n_438), .Y(n_434) );
INVxp67_ASAP7_75t_L g351 ( .A(n_320), .Y(n_351) );
INVx2_ASAP7_75t_SL g455 ( .A(n_320), .Y(n_455) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
OR2x2_ASAP7_75t_L g368 ( .A(n_322), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g466 ( .A(n_322), .B(n_465), .Y(n_466) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g339 ( .A(n_324), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_324), .B(n_348), .Y(n_364) );
INVx2_ASAP7_75t_L g391 ( .A(n_324), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .B1(n_332), .B2(n_334), .Y(n_326) );
NOR2xp33_ASAP7_75t_SL g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_328), .A2(n_402), .B1(n_415), .B2(n_417), .Y(n_414) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g424 ( .A(n_333), .B(n_425), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_341), .B(n_345), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g405 ( .A(n_338), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_338), .B(n_388), .Y(n_416) );
INVx1_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_342), .B(n_355), .Y(n_447) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI21xp33_ASAP7_75t_L g460 ( .A1(n_343), .A2(n_461), .B(n_463), .Y(n_460) );
OAI21xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_350), .B(n_358), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g404 ( .A(n_349), .Y(n_404) );
INVx1_ASAP7_75t_L g470 ( .A(n_349), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g443 ( .A(n_353), .Y(n_443) );
OR2x2_ASAP7_75t_L g454 ( .A(n_354), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND3xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .C(n_363), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_359), .A2(n_420), .B1(n_422), .B2(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g386 ( .A(n_360), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_361), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g399 ( .A(n_362), .Y(n_399) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_364), .B(n_368), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_364), .A2(n_427), .B1(n_430), .B2(n_433), .C(n_434), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_370), .B(n_371), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g375 ( .A(n_369), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_376), .B1(n_377), .B2(n_831), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g458 ( .A(n_380), .B(n_436), .Y(n_458) );
NAND4xp25_ASAP7_75t_L g381 ( .A(n_382), .B(n_412), .C(n_439), .D(n_459), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_395), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B1(n_389), .B2(n_390), .C(n_392), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_385), .A2(n_442), .B1(n_464), .B2(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g422 ( .A(n_388), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_388), .B(n_431), .Y(n_430) );
NAND2x1_ASAP7_75t_L g475 ( .A(n_388), .B(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_390), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g397 ( .A(n_394), .B(n_398), .Y(n_397) );
OAI21xp33_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_401), .B(n_406), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g425 ( .A(n_411), .Y(n_425) );
AOI211xp5_ASAP7_75t_L g439 ( .A1(n_411), .A2(n_440), .B(n_444), .C(n_450), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_426), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_414), .B(n_419), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g473 ( .A(n_421), .B(n_474), .Y(n_473) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx3_ASAP7_75t_L g477 ( .A(n_437), .Y(n_477) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI22xp33_ASAP7_75t_R g450 ( .A1(n_451), .A2(n_454), .B1(n_456), .B2(n_457), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g464 ( .A(n_453), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_467), .Y(n_459) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_694), .Y(n_479) );
NOR2xp67_ASAP7_75t_L g480 ( .A(n_481), .B(n_636), .Y(n_480) );
NAND3xp33_ASAP7_75t_SL g481 ( .A(n_482), .B(n_573), .C(n_618), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_529), .B(n_550), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_483), .A2(n_574), .B1(n_593), .B2(n_605), .Y(n_573) );
AOI22x1_ASAP7_75t_L g698 ( .A1(n_483), .A2(n_699), .B1(n_703), .B2(n_704), .Y(n_698) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_501), .Y(n_484) );
OR2x2_ASAP7_75t_L g659 ( .A(n_485), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .Y(n_485) );
OR2x2_ASAP7_75t_L g534 ( .A(n_486), .B(n_494), .Y(n_534) );
AND2x2_ASAP7_75t_L g577 ( .A(n_486), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g585 ( .A(n_486), .Y(n_585) );
BUFx2_ASAP7_75t_L g635 ( .A(n_486), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_490), .A2(n_526), .B(n_527), .Y(n_525) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_490), .A2(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g549 ( .A(n_491), .Y(n_549) );
AND2x2_ASAP7_75t_L g580 ( .A(n_494), .B(n_517), .Y(n_580) );
INVx1_ASAP7_75t_L g587 ( .A(n_494), .Y(n_587) );
INVx1_ASAP7_75t_L g592 ( .A(n_494), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_494), .B(n_585), .Y(n_654) );
INVx1_ASAP7_75t_L g675 ( .A(n_494), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_494), .B(n_578), .Y(n_745) );
INVx1_ASAP7_75t_L g638 ( .A(n_501), .Y(n_638) );
OR2x2_ASAP7_75t_L g690 ( .A(n_501), .B(n_654), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_517), .Y(n_501) );
AND2x2_ASAP7_75t_L g535 ( .A(n_502), .B(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g583 ( .A(n_502), .B(n_584), .Y(n_583) );
INVxp67_ASAP7_75t_L g589 ( .A(n_502), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_502), .B(n_532), .Y(n_666) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g578 ( .A(n_503), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_512), .B(n_515), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_508), .B(n_510), .Y(n_505) );
BUFx4f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_511), .B(n_524), .Y(n_523) );
INVx3_ASAP7_75t_L g532 ( .A(n_517), .Y(n_532) );
INVx1_ASAP7_75t_L g632 ( .A(n_517), .Y(n_632) );
AND2x2_ASAP7_75t_L g634 ( .A(n_517), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g652 ( .A(n_517), .B(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g674 ( .A(n_517), .B(n_675), .Y(n_674) );
NAND2x1p5_ASAP7_75t_SL g685 ( .A(n_517), .B(n_661), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_517), .B(n_592), .Y(n_775) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_525), .B(n_528), .Y(n_519) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_535), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_530), .A2(n_714), .B1(n_715), .B2(n_717), .Y(n_713) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_531), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_531), .B(n_770), .Y(n_769) );
OR2x2_ASAP7_75t_L g792 ( .A(n_531), .B(n_650), .Y(n_792) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g591 ( .A(n_532), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_532), .B(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g680 ( .A(n_532), .B(n_681), .Y(n_680) );
AND2x4_ASAP7_75t_L g631 ( .A(n_533), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g721 ( .A(n_534), .Y(n_721) );
OR2x2_ASAP7_75t_L g795 ( .A(n_534), .B(n_722), .Y(n_795) );
INVx1_ASAP7_75t_L g626 ( .A(n_535), .Y(n_626) );
INVx3_ASAP7_75t_L g630 ( .A(n_536), .Y(n_630) );
BUFx2_ASAP7_75t_L g641 ( .A(n_536), .Y(n_641) );
BUFx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g611 ( .A(n_537), .B(n_562), .Y(n_611) );
INVx2_ASAP7_75t_L g657 ( .A(n_537), .Y(n_657) );
INVx1_ASAP7_75t_L g689 ( .A(n_537), .Y(n_689) );
AND2x2_ASAP7_75t_L g702 ( .A(n_537), .B(n_599), .Y(n_702) );
AND2x2_ASAP7_75t_L g724 ( .A(n_537), .B(n_623), .Y(n_724) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_545), .B(n_548), .Y(n_539) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g715 ( .A(n_551), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_551), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g740 ( .A(n_551), .B(n_608), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_551), .B(n_742), .Y(n_741) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_562), .Y(n_551) );
INVx2_ASAP7_75t_L g597 ( .A(n_552), .Y(n_597) );
AND2x2_ASAP7_75t_L g624 ( .A(n_552), .B(n_625), .Y(n_624) );
AOI21x1_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_557), .B(n_560), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g598 ( .A(n_562), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g617 ( .A(n_562), .Y(n_617) );
INVx2_ASAP7_75t_L g625 ( .A(n_562), .Y(n_625) );
OR2x2_ASAP7_75t_L g645 ( .A(n_562), .B(n_599), .Y(n_645) );
AND2x2_ASAP7_75t_L g656 ( .A(n_562), .B(n_657), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_579), .B1(n_581), .B2(n_586), .C(n_588), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI32xp33_ASAP7_75t_L g686 ( .A1(n_576), .A2(n_590), .A3(n_687), .B1(n_690), .B2(n_691), .Y(n_686) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g676 ( .A(n_577), .Y(n_676) );
AND2x2_ASAP7_75t_L g712 ( .A(n_577), .B(n_591), .Y(n_712) );
INVx1_ASAP7_75t_L g776 ( .A(n_577), .Y(n_776) );
OR2x2_ASAP7_75t_L g650 ( .A(n_578), .B(n_585), .Y(n_650) );
INVx2_ASAP7_75t_L g661 ( .A(n_578), .Y(n_661) );
BUFx2_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g800 ( .A(n_580), .B(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVxp67_ASAP7_75t_L g787 ( .A(n_583), .Y(n_787) );
INVx1_ASAP7_75t_L g801 ( .A(n_583), .Y(n_801) );
OR2x2_ASAP7_75t_L g681 ( .A(n_584), .B(n_661), .Y(n_681) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_586), .B(n_681), .Y(n_703) );
INVx1_ASAP7_75t_L g734 ( .A(n_586), .Y(n_734) );
BUFx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g768 ( .A(n_587), .Y(n_768) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2x1_ASAP7_75t_L g737 ( .A(n_589), .B(n_738), .Y(n_737) );
OAI21xp5_ASAP7_75t_SL g759 ( .A1(n_590), .A2(n_760), .B(n_765), .Y(n_759) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
AND2x2_ASAP7_75t_L g669 ( .A(n_595), .B(n_611), .Y(n_669) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_595), .Y(n_799) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g701 ( .A(n_596), .Y(n_701) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g683 ( .A(n_597), .B(n_657), .Y(n_683) );
AND2x2_ASAP7_75t_L g754 ( .A(n_597), .B(n_625), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_598), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g682 ( .A(n_598), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g761 ( .A(n_598), .B(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g610 ( .A(n_599), .Y(n_610) );
INVx2_ASAP7_75t_L g623 ( .A(n_599), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_599), .B(n_614), .Y(n_671) );
AND2x2_ASAP7_75t_L g731 ( .A(n_599), .B(n_625), .Y(n_731) );
NAND2xp33_ASAP7_75t_SL g605 ( .A(n_606), .B(n_612), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g706 ( .A(n_609), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_609), .B(n_689), .Y(n_781) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g613 ( .A(n_610), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g742 ( .A(n_610), .B(n_657), .Y(n_742) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_616), .Y(n_612) );
OR2x2_ASAP7_75t_L g687 ( .A(n_613), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g644 ( .A(n_614), .Y(n_644) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g670 ( .A(n_617), .B(n_671), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_631), .B1(n_633), .B2(n_634), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_626), .B(n_627), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g633 ( .A(n_621), .B(n_630), .Y(n_633) );
BUFx2_ASAP7_75t_L g651 ( .A(n_621), .Y(n_651) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g662 ( .A(n_622), .Y(n_662) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g677 ( .A(n_624), .B(n_641), .Y(n_677) );
INVx2_ASAP7_75t_L g693 ( .A(n_624), .Y(n_693) );
AND2x2_ASAP7_75t_L g735 ( .A(n_624), .B(n_657), .Y(n_735) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g710 ( .A(n_630), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g757 ( .A(n_631), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g788 ( .A(n_632), .Y(n_788) );
INVx2_ASAP7_75t_L g727 ( .A(n_635), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_637), .B(n_646), .C(n_663), .D(n_678), .Y(n_636) );
NAND2xp33_ASAP7_75t_SL g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_639), .A2(n_717), .B1(n_733), .B2(n_735), .C(n_736), .Y(n_732) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2x1_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g714 ( .A(n_643), .Y(n_714) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx2_ASAP7_75t_L g707 ( .A(n_644), .Y(n_707) );
INVx2_ASAP7_75t_L g779 ( .A(n_645), .Y(n_779) );
AOI222xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_651), .B1(n_652), .B2(n_655), .C1(n_658), .C2(n_662), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g733 ( .A(n_649), .B(n_734), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_649), .A2(n_761), .B(n_763), .Y(n_760) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g772 ( .A(n_650), .B(n_716), .Y(n_772) );
OAI21xp33_ASAP7_75t_SL g746 ( .A1(n_651), .A2(n_672), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g665 ( .A(n_654), .B(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_SL g717 ( .A(n_654), .Y(n_717) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
BUFx2_ASAP7_75t_L g716 ( .A(n_657), .Y(n_716) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g722 ( .A(n_661), .Y(n_722) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_664), .A2(n_667), .B1(n_672), .B2(n_677), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_669), .A2(n_679), .B1(n_682), .B2(n_684), .C(n_686), .Y(n_678) );
INVx3_ASAP7_75t_R g793 ( .A(n_670), .Y(n_793) );
INVx1_ASAP7_75t_L g711 ( .A(n_671), .Y(n_711) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVxp67_ASAP7_75t_SL g728 ( .A(n_674), .Y(n_728) );
INVx1_ASAP7_75t_L g738 ( .A(n_674), .Y(n_738) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_683), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g756 ( .A(n_683), .Y(n_756) );
AND2x2_ASAP7_75t_L g784 ( .A(n_683), .B(n_731), .Y(n_784) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g778 ( .A(n_688), .B(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx3_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NOR2x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_750), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_732), .C(n_746), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_708), .C(n_718), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI21xp33_ASAP7_75t_L g709 ( .A1(n_699), .A2(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g749 ( .A(n_701), .Y(n_749) );
AND2x2_ASAP7_75t_L g790 ( .A(n_701), .B(n_779), .Y(n_790) );
NAND2x1_ASAP7_75t_L g748 ( .A(n_702), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g770 ( .A(n_707), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_713), .Y(n_708) );
INVx1_ASAP7_75t_L g762 ( .A(n_716), .Y(n_762) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_723), .B1(n_725), .B2(n_729), .Y(n_718) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g758 ( .A(n_722), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_724), .B(n_754), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g797 ( .A(n_730), .Y(n_797) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI22xp33_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_739), .B1(n_741), .B2(n_743), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_777), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_755), .B(n_757), .C(n_759), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OAI21xp33_ASAP7_75t_L g766 ( .A1(n_753), .A2(n_767), .B(n_769), .Y(n_766) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
O2A1O1Ixp5_ASAP7_75t_SL g777 ( .A1(n_757), .A2(n_778), .B(n_780), .C(n_782), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_761), .A2(n_766), .B1(n_771), .B2(n_773), .Y(n_765) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
OAI211xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_785), .B(n_789), .C(n_796), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B1(n_793), .B2(n_794), .Y(n_789) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI21xp5_ASAP7_75t_SL g796 ( .A1(n_797), .A2(n_798), .B(n_800), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI21xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_813), .B(n_815), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_808), .Y(n_803) );
BUFx2_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
INVx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
BUFx8_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
BUFx10_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_827), .Y(n_823) );
BUFx2_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
INVx4_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
endmodule