module real_aes_8118_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_0), .A2(n_72), .B1(n_193), .B2(n_194), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_0), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_1), .A2(n_262), .B(n_263), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_2), .A2(n_235), .B(n_237), .C(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_3), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g211 ( .A(n_4), .Y(n_211) );
AND2x6_ASAP7_75t_L g235 ( .A(n_4), .B(n_209), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_4), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g336 ( .A(n_5), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_6), .B(n_246), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_7), .A2(n_43), .B1(n_139), .B2(n_144), .Y(n_138) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_8), .A2(n_31), .B1(n_97), .B2(n_98), .Y(n_96) );
INVx1_ASAP7_75t_L g227 ( .A(n_9), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_10), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_11), .A2(n_281), .B(n_321), .C(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_12), .B(n_273), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_13), .Y(n_176) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_14), .A2(n_33), .B1(n_97), .B2(n_101), .Y(n_100) );
AOI22xp33_ASAP7_75t_L g113 ( .A1(n_15), .A2(n_47), .B1(n_114), .B2(n_119), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_16), .B(n_368), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g297 ( .A1(n_17), .A2(n_267), .B(n_298), .C(n_301), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_18), .A2(n_191), .B1(n_192), .B2(n_195), .Y(n_190) );
INVx1_ASAP7_75t_L g195 ( .A(n_18), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_19), .B(n_246), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_20), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_21), .B(n_246), .Y(n_282) );
INVx1_ASAP7_75t_L g548 ( .A(n_21), .Y(n_548) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_22), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_23), .Y(n_131) );
INVx1_ASAP7_75t_L g279 ( .A(n_24), .Y(n_279) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_25), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_26), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_27), .A2(n_59), .B1(n_159), .B2(n_164), .Y(n_158) );
INVx1_ASAP7_75t_L g365 ( .A(n_28), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_29), .Y(n_184) );
INVx2_ASAP7_75t_L g233 ( .A(n_30), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_32), .Y(n_316) );
OAI221xp5_ASAP7_75t_L g202 ( .A1(n_33), .A2(n_48), .B1(n_58), .B2(n_203), .C(n_204), .Y(n_202) );
INVxp67_ASAP7_75t_L g205 ( .A(n_33), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_34), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_35), .A2(n_267), .B(n_268), .C(n_270), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_36), .Y(n_112) );
XOR2xp5_ASAP7_75t_L g549 ( .A(n_37), .B(n_86), .Y(n_549) );
INVxp67_ASAP7_75t_L g366 ( .A(n_38), .Y(n_366) );
CKINVDCx14_ASAP7_75t_R g264 ( .A(n_39), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_40), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_41), .A2(n_237), .B(n_278), .C(n_285), .Y(n_277) );
AOI22xp5_ASAP7_75t_SL g538 ( .A1(n_41), .A2(n_86), .B1(n_186), .B2(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_41), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g333 ( .A1(n_42), .A2(n_248), .B(n_334), .C(n_335), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_44), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_45), .Y(n_362) );
INVx1_ASAP7_75t_L g296 ( .A(n_46), .Y(n_296) );
AO22x2_ASAP7_75t_L g104 ( .A1(n_48), .A2(n_69), .B1(n_97), .B2(n_101), .Y(n_104) );
INVxp67_ASAP7_75t_L g206 ( .A(n_48), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_49), .A2(n_190), .B1(n_196), .B2(n_197), .Y(n_189) );
INVx1_ASAP7_75t_L g196 ( .A(n_49), .Y(n_196) );
CKINVDCx14_ASAP7_75t_R g332 ( .A(n_50), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_51), .Y(n_137) );
INVx1_ASAP7_75t_L g209 ( .A(n_52), .Y(n_209) );
INVx1_ASAP7_75t_L g226 ( .A(n_53), .Y(n_226) );
INVx1_ASAP7_75t_SL g269 ( .A(n_54), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_55), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_56), .B(n_273), .Y(n_303) );
INVx1_ASAP7_75t_L g241 ( .A(n_57), .Y(n_241) );
AO22x2_ASAP7_75t_L g106 ( .A1(n_58), .A2(n_74), .B1(n_97), .B2(n_98), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_60), .A2(n_262), .B(n_331), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_61), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_62), .A2(n_262), .B(n_319), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_63), .A2(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g85 ( .A(n_64), .Y(n_85) );
CKINVDCx16_ASAP7_75t_R g276 ( .A(n_65), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_66), .A2(n_188), .B1(n_189), .B2(n_198), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g188 ( .A(n_66), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_67), .A2(n_262), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g322 ( .A(n_68), .Y(n_322) );
INVx2_ASAP7_75t_L g224 ( .A(n_70), .Y(n_224) );
INVx1_ASAP7_75t_L g313 ( .A(n_71), .Y(n_313) );
INVx1_ASAP7_75t_L g194 ( .A(n_72), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g81 ( .A1(n_73), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_73), .Y(n_82) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_73), .A2(n_237), .B(n_240), .C(n_250), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_75), .B(n_222), .Y(n_337) );
INVx1_ASAP7_75t_L g97 ( .A(n_76), .Y(n_97) );
INVx1_ASAP7_75t_L g99 ( .A(n_76), .Y(n_99) );
INVx2_ASAP7_75t_L g299 ( .A(n_77), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_199), .B1(n_212), .B2(n_532), .C(n_537), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_187), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_86), .B1(n_185), .B2(n_186), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_81), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
O2A1O1Ixp33_ASAP7_75t_SL g319 ( .A1(n_85), .A2(n_251), .B(n_265), .C(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g186 ( .A(n_86), .Y(n_186) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_147), .Y(n_86) );
NOR2xp33_ASAP7_75t_L g87 ( .A(n_88), .B(n_125), .Y(n_87) );
OAI221xp5_ASAP7_75t_SL g88 ( .A1(n_89), .A2(n_107), .B1(n_108), .B2(n_112), .C(n_113), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx11_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x6_ASAP7_75t_L g92 ( .A(n_93), .B(n_102), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
OR2x2_ASAP7_75t_L g151 ( .A(n_94), .B(n_152), .Y(n_151) );
OR2x2_ASAP7_75t_L g94 ( .A(n_95), .B(n_100), .Y(n_94) );
AND2x2_ASAP7_75t_L g111 ( .A(n_95), .B(n_100), .Y(n_111) );
AND2x2_ASAP7_75t_L g117 ( .A(n_95), .B(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g163 ( .A(n_96), .B(n_104), .Y(n_163) );
AND2x2_ASAP7_75t_L g169 ( .A(n_96), .B(n_100), .Y(n_169) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g101 ( .A(n_99), .Y(n_101) );
INVx2_ASAP7_75t_L g118 ( .A(n_100), .Y(n_118) );
INVx1_ASAP7_75t_L g146 ( .A(n_100), .Y(n_146) );
AND2x4_ASAP7_75t_L g110 ( .A(n_102), .B(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g116 ( .A(n_102), .B(n_117), .Y(n_116) );
AND2x6_ASAP7_75t_L g178 ( .A(n_102), .B(n_169), .Y(n_178) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
AND2x2_ASAP7_75t_L g130 ( .A(n_103), .B(n_106), .Y(n_130) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g123 ( .A(n_104), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_104), .B(n_106), .Y(n_136) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g124 ( .A(n_106), .Y(n_124) );
INVx1_ASAP7_75t_L g175 ( .A(n_106), .Y(n_175) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g143 ( .A(n_111), .B(n_123), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g156 ( .A(n_111), .B(n_130), .Y(n_156) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g122 ( .A(n_117), .B(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g129 ( .A(n_117), .B(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g134 ( .A(n_117), .B(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g174 ( .A(n_118), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
OAI221xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_131), .B1(n_132), .B2(n_137), .C(n_138), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g152 ( .A(n_130), .Y(n_152) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx2_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x6_ASAP7_75t_L g145 ( .A(n_136), .B(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx8_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g147 ( .A(n_148), .B(n_170), .Y(n_147) );
OAI221xp5_ASAP7_75t_SL g148 ( .A1(n_149), .A2(n_153), .B1(n_154), .B2(n_157), .C(n_158), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
AND2x4_ASAP7_75t_L g173 ( .A(n_163), .B(n_174), .Y(n_173) );
AND2x4_ASAP7_75t_L g182 ( .A(n_163), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
OAI222xp33_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_176), .B1(n_177), .B2(n_179), .C1(n_180), .C2(n_184), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx4f_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g183 ( .A(n_175), .Y(n_183) );
INVx2_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_189), .Y(n_198) );
INVx1_ASAP7_75t_L g197 ( .A(n_190), .Y(n_197) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_201), .Y(n_200) );
AND3x1_ASAP7_75t_SL g201 ( .A(n_202), .B(n_207), .C(n_210), .Y(n_201) );
INVxp67_ASAP7_75t_L g541 ( .A(n_202), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
INVx1_ASAP7_75t_SL g542 ( .A(n_207), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_207), .A2(n_545), .B(n_547), .Y(n_544) );
INVx1_ASAP7_75t_L g553 ( .A(n_207), .Y(n_553) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_208), .B(n_211), .Y(n_547) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_SL g552 ( .A(n_210), .B(n_553), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_211), .Y(n_210) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_214), .B(n_487), .Y(n_213) );
NOR4xp25_ASAP7_75t_L g214 ( .A(n_215), .B(n_424), .C(n_458), .D(n_474), .Y(n_214) );
NAND4xp25_ASAP7_75t_SL g215 ( .A(n_216), .B(n_350), .C(n_388), .D(n_404), .Y(n_215) );
AOI222xp33_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_288), .B1(n_325), .B2(n_338), .C1(n_343), .C2(n_349), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AOI31xp33_ASAP7_75t_L g520 ( .A1(n_218), .A2(n_521), .A3(n_522), .B(n_524), .Y(n_520) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_256), .Y(n_218) );
AND2x2_ASAP7_75t_L g495 ( .A(n_219), .B(n_258), .Y(n_495) );
BUFx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_SL g342 ( .A(n_220), .Y(n_342) );
AND2x2_ASAP7_75t_L g349 ( .A(n_220), .B(n_274), .Y(n_349) );
AND2x2_ASAP7_75t_L g409 ( .A(n_220), .B(n_259), .Y(n_409) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_228), .B(n_252), .Y(n_220) );
INVx3_ASAP7_75t_L g273 ( .A(n_221), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_221), .B(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_221), .B(n_316), .Y(n_315) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_222), .Y(n_260) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g358 ( .A(n_223), .Y(n_358) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AND2x2_ASAP7_75t_SL g255 ( .A(n_224), .B(n_225), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_236), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g275 ( .A1(n_230), .A2(n_255), .B(n_276), .C(n_277), .Y(n_275) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_230), .A2(n_310), .B(n_311), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
AND2x4_ASAP7_75t_L g262 ( .A(n_231), .B(n_235), .Y(n_262) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g284 ( .A(n_232), .Y(n_284) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g238 ( .A(n_233), .Y(n_238) );
INVx1_ASAP7_75t_L g302 ( .A(n_233), .Y(n_302) );
INVx1_ASAP7_75t_L g239 ( .A(n_234), .Y(n_239) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_234), .Y(n_244) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_234), .Y(n_246) );
INVx3_ASAP7_75t_L g281 ( .A(n_234), .Y(n_281) );
INVx4_ASAP7_75t_SL g251 ( .A(n_235), .Y(n_251) );
BUFx3_ASAP7_75t_L g285 ( .A(n_235), .Y(n_285) );
INVx5_ASAP7_75t_L g265 ( .A(n_237), .Y(n_265) );
AND2x6_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
BUFx3_ASAP7_75t_L g249 ( .A(n_238), .Y(n_249) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_238), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_245), .C(n_247), .Y(n_240) );
O2A1O1Ixp5_ASAP7_75t_L g312 ( .A1(n_242), .A2(n_247), .B(n_313), .C(n_314), .Y(n_312) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_242), .Y(n_535) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx4_ASAP7_75t_L g300 ( .A(n_244), .Y(n_300) );
INVx4_ASAP7_75t_L g267 ( .A(n_246), .Y(n_267) );
INVx2_ASAP7_75t_L g334 ( .A(n_246), .Y(n_334) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g323 ( .A(n_249), .Y(n_323) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_251), .A2(n_264), .B(n_265), .C(n_266), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_SL g295 ( .A1(n_251), .A2(n_265), .B(n_296), .C(n_297), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_SL g331 ( .A1(n_251), .A2(n_265), .B(n_332), .C(n_333), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_SL g361 ( .A1(n_251), .A2(n_265), .B(n_362), .C(n_363), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_251), .B(n_283), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g368 ( .A(n_254), .Y(n_368) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g308 ( .A(n_255), .Y(n_308) );
OA21x2_ASAP7_75t_L g329 ( .A1(n_255), .A2(n_330), .B(n_337), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_256), .B(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_257), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_257), .B(n_353), .Y(n_399) );
AND2x2_ASAP7_75t_L g492 ( .A(n_257), .B(n_432), .Y(n_492) );
OAI321xp33_ASAP7_75t_L g526 ( .A1(n_257), .A2(n_342), .A3(n_499), .B1(n_527), .B2(n_529), .C(n_530), .Y(n_526) );
NAND4xp25_ASAP7_75t_L g530 ( .A(n_257), .B(n_328), .C(n_439), .D(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_274), .Y(n_257) );
AND2x2_ASAP7_75t_L g394 ( .A(n_258), .B(n_340), .Y(n_394) );
AND2x2_ASAP7_75t_L g413 ( .A(n_258), .B(n_342), .Y(n_413) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g341 ( .A(n_259), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g369 ( .A(n_259), .B(n_274), .Y(n_369) );
AND2x2_ASAP7_75t_L g455 ( .A(n_259), .B(n_340), .Y(n_455) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B(n_272), .Y(n_259) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_260), .A2(n_294), .B(n_303), .Y(n_293) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_260), .A2(n_318), .B(n_324), .Y(n_317) );
BUFx2_ASAP7_75t_L g360 ( .A(n_262), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_267), .B(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx3_ASAP7_75t_SL g340 ( .A(n_274), .Y(n_340) );
AND2x2_ASAP7_75t_L g387 ( .A(n_274), .B(n_374), .Y(n_387) );
OR2x2_ASAP7_75t_L g420 ( .A(n_274), .B(n_342), .Y(n_420) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_274), .Y(n_427) );
AND2x2_ASAP7_75t_L g456 ( .A(n_274), .B(n_341), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_274), .B(n_429), .Y(n_471) );
AND2x2_ASAP7_75t_L g503 ( .A(n_274), .B(n_495), .Y(n_503) );
AND2x2_ASAP7_75t_L g512 ( .A(n_274), .B(n_354), .Y(n_512) );
OR2x6_ASAP7_75t_L g274 ( .A(n_275), .B(n_286), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B(n_282), .C(n_283), .Y(n_278) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_280), .A2(n_300), .B1(n_365), .B2(n_366), .Y(n_364) );
INVx5_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_281), .B(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_283), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_284), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_304), .Y(n_289) );
INVx1_ASAP7_75t_SL g480 ( .A(n_290), .Y(n_480) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g345 ( .A(n_291), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g327 ( .A(n_292), .B(n_306), .Y(n_327) );
AND2x2_ASAP7_75t_L g416 ( .A(n_292), .B(n_329), .Y(n_416) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g386 ( .A(n_293), .B(n_317), .Y(n_386) );
OR2x2_ASAP7_75t_L g397 ( .A(n_293), .B(n_329), .Y(n_397) );
AND2x2_ASAP7_75t_L g423 ( .A(n_293), .B(n_329), .Y(n_423) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_293), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_300), .B(n_322), .Y(n_321) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_304), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_304), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g396 ( .A(n_305), .B(n_397), .Y(n_396) );
AOI322xp5_ASAP7_75t_L g482 ( .A1(n_305), .A2(n_386), .A3(n_392), .B1(n_423), .B2(n_473), .C1(n_483), .C2(n_485), .Y(n_482) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_317), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_306), .B(n_328), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_306), .B(n_329), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_306), .B(n_346), .Y(n_403) );
AND2x2_ASAP7_75t_L g457 ( .A(n_306), .B(n_423), .Y(n_457) );
INVx1_ASAP7_75t_L g461 ( .A(n_306), .Y(n_461) );
AND2x2_ASAP7_75t_L g473 ( .A(n_306), .B(n_317), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_306), .B(n_345), .Y(n_505) );
INVx4_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g370 ( .A(n_307), .B(n_317), .Y(n_370) );
BUFx3_ASAP7_75t_L g384 ( .A(n_307), .Y(n_384) );
AND3x2_ASAP7_75t_L g466 ( .A(n_307), .B(n_446), .C(n_467), .Y(n_466) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B(n_315), .Y(n_307) );
NAND3xp33_ASAP7_75t_L g326 ( .A(n_317), .B(n_327), .C(n_328), .Y(n_326) );
INVx1_ASAP7_75t_SL g346 ( .A(n_317), .Y(n_346) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_317), .Y(n_451) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g445 ( .A(n_327), .B(n_446), .Y(n_445) );
INVxp67_ASAP7_75t_L g452 ( .A(n_327), .Y(n_452) );
AND2x2_ASAP7_75t_L g490 ( .A(n_328), .B(n_468), .Y(n_490) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx3_ASAP7_75t_L g371 ( .A(n_329), .Y(n_371) );
AND2x2_ASAP7_75t_L g446 ( .A(n_329), .B(n_346), .Y(n_446) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
OR2x2_ASAP7_75t_L g390 ( .A(n_340), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g509 ( .A(n_340), .B(n_409), .Y(n_509) );
AND2x2_ASAP7_75t_L g523 ( .A(n_340), .B(n_342), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_341), .B(n_354), .Y(n_464) );
AND2x2_ASAP7_75t_L g511 ( .A(n_341), .B(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g374 ( .A(n_342), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g391 ( .A(n_342), .B(n_354), .Y(n_391) );
INVx1_ASAP7_75t_L g401 ( .A(n_342), .Y(n_401) );
AND2x2_ASAP7_75t_L g432 ( .A(n_342), .B(n_354), .Y(n_432) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI221xp5_ASAP7_75t_L g474 ( .A1(n_344), .A2(n_475), .B1(n_479), .B2(n_481), .C(n_482), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_345), .B(n_347), .Y(n_344) );
AND2x2_ASAP7_75t_L g378 ( .A(n_345), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_348), .B(n_385), .Y(n_528) );
AOI322xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_370), .A3(n_371), .B1(n_372), .B2(n_378), .C1(n_380), .C2(n_387), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_369), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g408 ( .A(n_353), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_353), .B(n_419), .Y(n_418) );
O2A1O1Ixp33_ASAP7_75t_L g442 ( .A1(n_353), .A2(n_369), .B(n_443), .C(n_444), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_353), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_353), .B(n_413), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_353), .B(n_495), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_353), .B(n_523), .Y(n_522) );
BUFx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_354), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_354), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g484 ( .A(n_354), .B(n_371), .Y(n_484) );
OA21x2_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_359), .B(n_367), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AO21x2_ASAP7_75t_L g375 ( .A1(n_356), .A2(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g376 ( .A(n_359), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_367), .Y(n_377) );
INVx1_ASAP7_75t_L g459 ( .A(n_369), .Y(n_459) );
OAI31xp33_ASAP7_75t_L g469 ( .A1(n_369), .A2(n_394), .A3(n_470), .B(n_472), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_369), .B(n_375), .Y(n_521) );
INVx1_ASAP7_75t_SL g382 ( .A(n_370), .Y(n_382) );
AND2x2_ASAP7_75t_L g415 ( .A(n_370), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g496 ( .A(n_370), .B(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g381 ( .A(n_371), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g406 ( .A(n_371), .Y(n_406) );
AND2x2_ASAP7_75t_L g433 ( .A(n_371), .B(n_386), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_371), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g525 ( .A(n_371), .B(n_473), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_373), .B(n_443), .Y(n_516) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g412 ( .A(n_375), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g430 ( .A(n_375), .Y(n_430) );
NAND2xp33_ASAP7_75t_SL g380 ( .A(n_381), .B(n_383), .Y(n_380) );
OAI211xp5_ASAP7_75t_SL g424 ( .A1(n_382), .A2(n_425), .B(n_431), .C(n_447), .Y(n_424) );
OR2x2_ASAP7_75t_L g499 ( .A(n_382), .B(n_480), .Y(n_499) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
CKINVDCx16_ASAP7_75t_R g436 ( .A(n_384), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_384), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g405 ( .A(n_386), .B(n_406), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_392), .B(n_395), .C(n_398), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g439 ( .A(n_391), .Y(n_439) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_394), .B(n_432), .Y(n_437) );
INVx1_ASAP7_75t_L g443 ( .A(n_394), .Y(n_443) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g402 ( .A(n_397), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g435 ( .A(n_397), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g497 ( .A(n_397), .Y(n_497) );
AOI21xp33_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_400), .B(n_402), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_400), .A2(n_411), .B(n_414), .Y(n_410) );
AOI211xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B(n_410), .C(n_417), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_405), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_408), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g421 ( .A(n_409), .Y(n_421) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_411), .A2(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_416), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g441 ( .A(n_416), .Y(n_441) );
AOI21xp33_ASAP7_75t_SL g417 ( .A1(n_418), .A2(n_421), .B(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g472 ( .A(n_423), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_429), .B(n_455), .Y(n_481) );
AND2x2_ASAP7_75t_L g494 ( .A(n_429), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g508 ( .A(n_429), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g518 ( .A(n_429), .B(n_456), .Y(n_518) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI211xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_434), .C(n_442), .Y(n_431) );
INVx1_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_438), .B2(n_440), .Y(n_434) );
OR2x2_ASAP7_75t_L g440 ( .A(n_436), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_436), .B(n_497), .Y(n_519) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g513 ( .A(n_446), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_453), .B1(n_456), .B2(n_457), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g531 ( .A(n_451), .Y(n_531) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g477 ( .A(n_455), .Y(n_477) );
OAI211xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_460), .B(n_462), .C(n_469), .Y(n_458) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVxp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVxp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_477), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NOR5xp2_ASAP7_75t_L g487 ( .A(n_488), .B(n_506), .C(n_514), .D(n_520), .E(n_526), .Y(n_487) );
OAI211xp5_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_491), .B(n_493), .C(n_500), .Y(n_488) );
INVxp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_496), .B(n_498), .Y(n_493) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_503), .B(n_504), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_503), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AOI21xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_510), .B(n_513), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_SL g529 ( .A(n_509), .Y(n_529) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_517), .B(n_519), .Y(n_514) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g546 ( .A(n_535), .Y(n_546) );
OAI322xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_540), .A3(n_542), .B1(n_543), .B2(n_548), .C1(n_549), .C2(n_550), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_551), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
endmodule