module fake_aes_5069_n_22 (n_1, n_2, n_4, n_3, n_5, n_0, n_22);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_22;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_6;
wire n_7;
INVx1_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
NAND2xp33_ASAP7_75t_L g7 ( .A(n_0), .B(n_5), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_2), .Y(n_8) );
OR2x6_ASAP7_75t_L g9 ( .A(n_2), .B(n_4), .Y(n_9) );
AOI21xp5_ASAP7_75t_L g10 ( .A1(n_8), .A2(n_0), .B(n_1), .Y(n_10) );
O2A1O1Ixp5_ASAP7_75t_L g11 ( .A1(n_8), .A2(n_0), .B(n_1), .C(n_2), .Y(n_11) );
NOR2x1_ASAP7_75t_L g12 ( .A(n_6), .B(n_1), .Y(n_12) );
AND2x4_ASAP7_75t_L g13 ( .A(n_12), .B(n_9), .Y(n_13) );
NAND3xp33_ASAP7_75t_SL g14 ( .A(n_11), .B(n_9), .C(n_7), .Y(n_14) );
INVxp67_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_13), .B(n_9), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_16), .B(n_14), .Y(n_17) );
OAI21xp5_ASAP7_75t_SL g18 ( .A1(n_17), .A2(n_16), .B(n_15), .Y(n_18) );
AOI211xp5_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_7), .B(n_10), .C(n_3), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_18), .B(n_3), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
AOI21xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_4), .B(n_20), .Y(n_22) );
endmodule