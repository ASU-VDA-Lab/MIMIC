module fake_netlist_1_882_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_0), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
INVx1_ASAP7_75t_SL g16 ( .A(n_3), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_10), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_11), .B(n_0), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_14), .B(n_1), .Y(n_20) );
INVx2_ASAP7_75t_SL g21 ( .A(n_13), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_17), .Y(n_22) );
INVx1_ASAP7_75t_SL g23 ( .A(n_12), .Y(n_23) );
OAI21xp5_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_17), .B(n_15), .Y(n_24) );
A2O1A1Ixp33_ASAP7_75t_L g25 ( .A1(n_18), .A2(n_16), .B(n_3), .C(n_2), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_20), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_26) );
AND2x4_ASAP7_75t_L g27 ( .A(n_21), .B(n_9), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
INVx3_ASAP7_75t_SL g30 ( .A(n_25), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVxp67_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_32), .B(n_30), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_31), .B(n_24), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_34), .Y(n_35) );
NAND3xp33_ASAP7_75t_L g36 ( .A(n_33), .B(n_26), .C(n_22), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
NOR3xp33_ASAP7_75t_L g38 ( .A(n_37), .B(n_19), .C(n_36), .Y(n_38) );
AOI22xp33_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_37), .B1(n_18), .B2(n_23), .Y(n_39) );
endmodule