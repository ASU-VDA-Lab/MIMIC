module fake_jpeg_5552_n_336 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_5),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_45),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_7),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_46),
.A2(n_20),
.B(n_25),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_6),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_14),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_55),
.Y(n_78)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_30),
.B1(n_24),
.B2(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_23),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_62),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_66),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_35),
.B1(n_24),
.B2(n_30),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_93),
.C(n_26),
.Y(n_110)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_67),
.B(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_30),
.B1(n_33),
.B2(n_31),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_79),
.B1(n_86),
.B2(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_81),
.Y(n_128)
);

INVx5_ASAP7_75t_SL g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_17),
.B1(n_33),
.B2(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_37),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_82),
.B(n_87),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_84),
.B(n_96),
.Y(n_132)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_15),
.B1(n_25),
.B2(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_39),
.B(n_28),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_97),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_90),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_14),
.B(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_17),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_102),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_57),
.A2(n_15),
.B1(n_20),
.B2(n_21),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_18),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_48),
.A2(n_36),
.B1(n_27),
.B2(n_26),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_114),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_131),
.Y(n_151)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_118),
.Y(n_155)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_72),
.Y(n_146)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_27),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_104),
.Y(n_157)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_133),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_23),
.C(n_1),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

BUFx16f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_137),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_23),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_139),
.A2(n_86),
.B(n_101),
.Y(n_153)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_145),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_141),
.B(n_143),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_146),
.B(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_148),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_150),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_64),
.B1(n_63),
.B2(n_75),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_159),
.B1(n_107),
.B2(n_120),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_153),
.A2(n_8),
.B(n_13),
.Y(n_209)
);

CKINVDCx12_ASAP7_75t_R g154 ( 
.A(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_158),
.Y(n_181)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_111),
.A2(n_100),
.B1(n_63),
.B2(n_79),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_58),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_173),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_110),
.B1(n_127),
.B2(n_132),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_166),
.Y(n_196)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_100),
.B1(n_75),
.B2(n_68),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_123),
.B1(n_114),
.B2(n_131),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_170),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_119),
.B(n_88),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_172),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_60),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_90),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_112),
.B(n_9),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_113),
.B(n_0),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_151),
.Y(n_206)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_113),
.B(n_91),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

BUFx4f_ASAP7_75t_SL g180 ( 
.A(n_176),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_192),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_145),
.B(n_125),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_182),
.B(n_206),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_173),
.A2(n_122),
.B(n_109),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_183),
.A2(n_210),
.B(n_142),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_184),
.A2(n_204),
.B1(n_201),
.B2(n_203),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_138),
.B1(n_139),
.B2(n_91),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_188),
.A2(n_143),
.B1(n_99),
.B2(n_144),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_200),
.B1(n_155),
.B2(n_166),
.Y(n_224)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_128),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_197),
.C(n_204),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_139),
.B(n_138),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_210),
.B(n_177),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_71),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_146),
.A2(n_118),
.B1(n_71),
.B2(n_99),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_203),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_8),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_207),
.Y(n_241)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_183),
.B(n_189),
.Y(n_238)
);

NAND2x1p5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_0),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_115),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_151),
.B(n_10),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_161),
.C(n_147),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_115),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_220),
.B(n_189),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_228),
.C(n_233),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_210),
.A2(n_168),
.B(n_167),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_185),
.A2(n_150),
.B1(n_149),
.B2(n_141),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_222),
.A2(n_208),
.B(n_227),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_231),
.B(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_237),
.Y(n_248)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_227),
.B1(n_236),
.B2(n_243),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_185),
.A2(n_144),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_0),
.C(n_1),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_177),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_213),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_205),
.A2(n_2),
.B(n_3),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_180),
.A2(n_2),
.B(n_4),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_2),
.C(n_10),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_12),
.C(n_13),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_187),
.C(n_179),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_180),
.A2(n_191),
.B1(n_188),
.B2(n_200),
.Y(n_236)
);

OA21x2_ASAP7_75t_L g237 ( 
.A1(n_184),
.A2(n_199),
.B(n_209),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_240),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_186),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_239),
.Y(n_256)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_247),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_199),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_249),
.A2(n_252),
.B(n_254),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_194),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

OA22x2_ASAP7_75t_L g251 ( 
.A1(n_226),
.A2(n_199),
.B1(n_198),
.B2(n_208),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_251),
.A2(n_218),
.B1(n_235),
.B2(n_240),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_178),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_258),
.B(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_215),
.B(n_190),
.C(n_181),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_264),
.C(n_217),
.Y(n_268)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_262),
.A2(n_265),
.B(n_266),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_222),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_215),
.B(n_202),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_241),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_232),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_271),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_216),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_263),
.A2(n_238),
.B1(n_237),
.B2(n_220),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_233),
.C(n_228),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_279),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_237),
.B1(n_234),
.B2(n_225),
.Y(n_278)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_261),
.C(n_260),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_285),
.B(n_245),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_262),
.A2(n_218),
.B1(n_231),
.B2(n_248),
.Y(n_283)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_257),
.A2(n_251),
.B1(n_266),
.B2(n_252),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_284),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_251),
.A2(n_267),
.B1(n_249),
.B2(n_254),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_273),
.B(n_246),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_288),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_251),
.Y(n_288)
);

BUFx12_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_270),
.A2(n_245),
.B(n_249),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_294),
.B1(n_296),
.B2(n_284),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

OAI31xp33_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_254),
.A3(n_267),
.B(n_255),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_298),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_268),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_304),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_289),
.B(n_256),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_298),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_271),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_309),
.Y(n_314)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_272),
.C(n_269),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_306),
.A2(n_299),
.B1(n_287),
.B2(n_295),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_279),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_285),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_276),
.C(n_253),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_273),
.B(n_278),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_283),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_312),
.A2(n_316),
.B1(n_318),
.B2(n_320),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_317),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_300),
.A2(n_288),
.B1(n_290),
.B2(n_275),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_302),
.A2(n_290),
.B1(n_274),
.B2(n_280),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_292),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_319),
.B(n_307),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_306),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_313),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_320),
.A2(n_310),
.B1(n_256),
.B2(n_307),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_323),
.B(n_326),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_314),
.C(n_308),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_258),
.B1(n_305),
.B2(n_253),
.Y(n_326)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_328),
.Y(n_332)
);

NAND4xp25_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_330),
.C(n_321),
.D(n_322),
.Y(n_331)
);

XOR2x2_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_314),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_325),
.B(n_327),
.C(n_244),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_332),
.B(n_244),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_244),
.Y(n_336)
);


endmodule