module fake_netlist_5_2106_n_1926 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1926);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1926;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_368;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g193 ( 
.A(n_89),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_19),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_133),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_19),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_150),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_81),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_61),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_44),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_103),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_52),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_114),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_122),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_17),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_105),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_96),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_34),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_146),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_156),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_119),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_71),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_113),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_138),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_145),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_44),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_10),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_124),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_110),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_161),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_144),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_136),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_140),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_27),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_36),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_168),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_8),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_62),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_123),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_11),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_34),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_93),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_91),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_153),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_121),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_109),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_137),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_48),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_84),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_29),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_6),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_126),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_106),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_22),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_54),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_22),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_66),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_149),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_54),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_180),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_175),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_139),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_25),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_21),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_177),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_2),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_117),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_154),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_125),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_38),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_151),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_12),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_172),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_118),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_72),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_8),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_189),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_57),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_97),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_43),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_53),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_26),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_24),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_10),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_40),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_18),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_73),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_132),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_186),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_169),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_11),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_170),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_13),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_86),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_77),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_38),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_62),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_184),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_141),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_56),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_129),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_135),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_176),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_12),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_59),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_116),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_112),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_167),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_39),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_181),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_39),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_14),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_18),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_163),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_165),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_3),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_15),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_55),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_66),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_171),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_32),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_130),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_142),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_5),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_65),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_183),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_155),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_64),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_53),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_48),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_57),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_9),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_82),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_43),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_69),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_67),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_76),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_17),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_128),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_31),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_131),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_69),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_55),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_61),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_152),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_6),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_191),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_80),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_72),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_16),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_7),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_88),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_64),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_178),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_2),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_68),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_190),
.Y(n_354)
);

BUFx2_ASAP7_75t_SL g355 ( 
.A(n_31),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_87),
.Y(n_356)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_147),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_158),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_73),
.Y(n_359)
);

BUFx10_ASAP7_75t_L g360 ( 
.A(n_115),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_26),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_50),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_0),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_185),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_127),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_35),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_16),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_20),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_41),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_107),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_162),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_71),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_59),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_33),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_28),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_30),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_4),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_20),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_47),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_85),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_40),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_30),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_1),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_95),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_192),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_211),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_278),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_278),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_278),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_215),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_212),
.B(n_0),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_278),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_195),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_197),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_216),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_199),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_205),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_269),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_255),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_325),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_275),
.B(n_1),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_278),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_223),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_207),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_210),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_214),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_253),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_281),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_221),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_281),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_281),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_225),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_223),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_226),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_281),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_R g416 ( 
.A(n_342),
.B(n_104),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_228),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_281),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_364),
.B(n_193),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_229),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_349),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_365),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_232),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_239),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_208),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_208),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_337),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_326),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_337),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_337),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_337),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_242),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_248),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_364),
.B(n_193),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_194),
.B(n_3),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_383),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_257),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_200),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_337),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_259),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_352),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_352),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_194),
.B(n_4),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_352),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_266),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_352),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_271),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_381),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_274),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_252),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_296),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_260),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_298),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_355),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_326),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_300),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_313),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_303),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_213),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_313),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_R g467 ( 
.A(n_304),
.B(n_187),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_346),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_346),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_307),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_319),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_320),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_323),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_324),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_330),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_196),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_200),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_196),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_355),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_198),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_336),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_419),
.B(n_344),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_438),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_315),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_410),
.B(n_213),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_410),
.B(n_235),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_438),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_438),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_235),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_387),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_426),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_411),
.B(n_289),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_438),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_438),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_438),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_477),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_477),
.B(n_200),
.Y(n_498)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_398),
.Y(n_499)
);

NOR2x1_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_289),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_411),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_434),
.B(n_345),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_387),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_447),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_388),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_447),
.B(n_264),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_388),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_453),
.B(n_389),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_389),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_392),
.B(n_351),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_403),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_392),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_393),
.B(n_321),
.Y(n_513)
);

INVx6_ASAP7_75t_L g514 ( 
.A(n_398),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_453),
.B(n_359),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_402),
.B(n_408),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_402),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_408),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_415),
.B(n_361),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_415),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_428),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_418),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_418),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_427),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_427),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

CKINVDCx8_ASAP7_75t_R g528 ( 
.A(n_461),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_429),
.B(n_430),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_430),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_431),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_431),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_439),
.B(n_264),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_439),
.B(n_276),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_452),
.B(n_340),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_400),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_441),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_442),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_442),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_444),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_444),
.B(n_356),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_445),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_445),
.B(n_358),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_449),
.B(n_276),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_449),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_450),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_450),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_455),
.A2(n_203),
.B(n_201),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_456),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_386),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_461),
.B(n_243),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_456),
.B(n_370),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_460),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_460),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_435),
.B(n_380),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_476),
.B(n_285),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_463),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_476),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_501),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_547),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_552),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_SL g564 ( 
.A1(n_557),
.A2(n_401),
.B1(n_407),
.B2(n_436),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_513),
.B(n_394),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_487),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_501),
.Y(n_567)
);

OAI22x1_ASAP7_75t_L g568 ( 
.A1(n_536),
.A2(n_517),
.B1(n_522),
.B2(n_511),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_485),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_487),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_537),
.B(n_396),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_547),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_487),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_547),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_L g575 ( 
.A(n_557),
.B(n_416),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_506),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_482),
.B(n_397),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_506),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_506),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_482),
.B(n_502),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_502),
.B(n_404),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_501),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_510),
.B(n_405),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_485),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_487),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_528),
.B(n_432),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_537),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_510),
.B(n_406),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_549),
.B(n_443),
.C(n_391),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_515),
.B(n_409),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_487),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_515),
.A2(n_367),
.B1(n_335),
.B2(n_362),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_489),
.B(n_412),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_542),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_489),
.B(n_414),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_506),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_507),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_508),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_485),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_507),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_542),
.B(n_417),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_490),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_544),
.B(n_554),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_487),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_528),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_485),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_490),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_507),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_503),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_489),
.A2(n_206),
.B1(n_361),
.B2(n_222),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_536),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_503),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_486),
.B(n_201),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_505),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_487),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_505),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_508),
.B(n_459),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_509),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_544),
.B(n_420),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_508),
.B(n_520),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_528),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_511),
.B(n_423),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_517),
.B(n_424),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_522),
.B(n_433),
.Y(n_624)
);

AND3x2_ASAP7_75t_L g625 ( 
.A(n_491),
.B(n_291),
.C(n_285),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_504),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_554),
.B(n_440),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_SL g628 ( 
.A(n_553),
.B(n_437),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_519),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_486),
.B(n_446),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_499),
.B(n_448),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_509),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_518),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_486),
.B(n_203),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_498),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_519),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_519),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_518),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_499),
.B(n_451),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_530),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_491),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_523),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_523),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_484),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_530),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_530),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_498),
.Y(n_647)
);

BUFx4f_ASAP7_75t_L g648 ( 
.A(n_549),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_524),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_531),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_504),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_486),
.B(n_454),
.Y(n_652)
);

AND2x6_ASAP7_75t_L g653 ( 
.A(n_500),
.B(n_291),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_524),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_499),
.B(n_471),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_525),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_525),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_526),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_558),
.A2(n_206),
.B1(n_222),
.B2(n_198),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_526),
.Y(n_660)
);

INVxp33_ASAP7_75t_L g661 ( 
.A(n_484),
.Y(n_661)
);

OR2x6_ASAP7_75t_L g662 ( 
.A(n_499),
.B(n_218),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_527),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_531),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_520),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_499),
.B(n_472),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_504),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g668 ( 
.A(n_520),
.B(n_390),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_492),
.B(n_473),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_504),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_531),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_492),
.B(n_474),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_492),
.B(n_479),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_527),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_514),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_540),
.Y(n_676)
);

BUFx4f_ASAP7_75t_L g677 ( 
.A(n_549),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_539),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_514),
.B(n_475),
.Y(n_679)
);

CKINVDCx6p67_ASAP7_75t_R g680 ( 
.A(n_492),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_539),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_540),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_500),
.B(n_481),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_514),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_541),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_541),
.B(n_238),
.Y(n_686)
);

BUFx4f_ASAP7_75t_L g687 ( 
.A(n_549),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_504),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_514),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_514),
.Y(n_690)
);

OAI21xp33_ASAP7_75t_L g691 ( 
.A1(n_560),
.A2(n_277),
.B(n_273),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_543),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_539),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_555),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_560),
.B(n_463),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_543),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_516),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_555),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_546),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_558),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_L g701 ( 
.A(n_498),
.B(n_467),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_558),
.B(n_466),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_546),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_548),
.B(n_241),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_558),
.A2(n_302),
.B1(n_277),
.B2(n_283),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_548),
.B(n_268),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_550),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_533),
.B(n_400),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_549),
.A2(n_302),
.B1(n_283),
.B2(n_288),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_550),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_551),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_551),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_533),
.B(n_466),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_576),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_580),
.B(n_533),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_668),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_594),
.A2(n_462),
.B1(n_464),
.B2(n_470),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_593),
.B(n_458),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_675),
.B(n_218),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_576),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_581),
.B(n_533),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_577),
.B(n_457),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_603),
.B(n_534),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_587),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_583),
.B(n_588),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_709),
.B(n_357),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_675),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_684),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_587),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_601),
.B(n_395),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_589),
.A2(n_295),
.B(n_338),
.C(n_292),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_598),
.B(n_286),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_619),
.B(n_399),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_569),
.Y(n_734)
);

OR2x2_ASAP7_75t_SL g735 ( 
.A(n_665),
.B(n_273),
.Y(n_735)
);

AND2x6_ASAP7_75t_SL g736 ( 
.A(n_622),
.B(n_288),
.Y(n_736)
);

NAND2x1p5_ASAP7_75t_L g737 ( 
.A(n_635),
.B(n_219),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_598),
.A2(n_421),
.B1(n_422),
.B2(n_338),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_L g739 ( 
.A(n_653),
.B(n_357),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_578),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_635),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_627),
.B(n_562),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_579),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_562),
.B(n_534),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_700),
.B(n_312),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_623),
.B(n_256),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_579),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_596),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_572),
.B(n_534),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_620),
.A2(n_316),
.B(n_290),
.C(n_374),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_641),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_596),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_572),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_624),
.B(n_202),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_684),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_574),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_569),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_569),
.B(n_219),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_668),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_602),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_684),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_574),
.B(n_534),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_602),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_620),
.B(n_545),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_631),
.B(n_384),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_584),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_617),
.B(n_545),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_584),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_589),
.A2(n_292),
.B(n_295),
.C(n_354),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_584),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_639),
.B(n_243),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_575),
.B(n_545),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_655),
.B(n_243),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_666),
.B(n_371),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_565),
.B(n_204),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_607),
.B(n_545),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_607),
.B(n_556),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_609),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_617),
.B(n_478),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_605),
.B(n_621),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_609),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_612),
.B(n_556),
.Y(n_782)
);

INVxp67_ASAP7_75t_SL g783 ( 
.A(n_599),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_612),
.Y(n_784)
);

O2A1O1Ixp5_ASAP7_75t_L g785 ( 
.A1(n_648),
.A2(n_538),
.B(n_334),
.C(n_262),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_599),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_611),
.B(n_217),
.C(n_209),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_614),
.B(n_538),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_599),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_614),
.B(n_538),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_610),
.B(n_231),
.C(n_230),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_635),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_616),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_679),
.B(n_371),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_595),
.B(n_233),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_606),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_606),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_613),
.A2(n_270),
.B1(n_385),
.B2(n_220),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_606),
.Y(n_799)
);

O2A1O1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_691),
.A2(n_290),
.B(n_316),
.C(n_332),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_641),
.Y(n_801)
);

NAND2x1p5_ASAP7_75t_L g802 ( 
.A(n_635),
.B(n_220),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_564),
.B(n_371),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_684),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_702),
.B(n_478),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_616),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_564),
.B(n_265),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_690),
.B(n_265),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_618),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_618),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_632),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_690),
.B(n_630),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_632),
.Y(n_813)
);

CKINVDCx16_ASAP7_75t_R g814 ( 
.A(n_586),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_669),
.B(n_265),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_633),
.B(n_538),
.Y(n_816)
);

NOR2x1p5_ASAP7_75t_L g817 ( 
.A(n_563),
.B(n_234),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_633),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_638),
.B(n_559),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_713),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_L g821 ( 
.A(n_653),
.B(n_357),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_613),
.B(n_224),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_697),
.B(n_265),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_638),
.B(n_559),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_L g825 ( 
.A(n_689),
.B(n_516),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_673),
.B(n_360),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_642),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_713),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_642),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_643),
.Y(n_830)
);

AO22x2_ASAP7_75t_L g831 ( 
.A1(n_613),
.A2(n_270),
.B1(n_287),
.B2(n_299),
.Y(n_831)
);

NOR3xp33_ASAP7_75t_L g832 ( 
.A(n_644),
.B(n_237),
.C(n_236),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_643),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_649),
.B(n_559),
.Y(n_834)
);

AOI22x1_ASAP7_75t_L g835 ( 
.A1(n_613),
.A2(n_287),
.B1(n_262),
.B2(n_258),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_566),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_649),
.B(n_559),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_571),
.B(n_590),
.Y(n_838)
);

BUFx12f_ASAP7_75t_SL g839 ( 
.A(n_662),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_654),
.B(n_559),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_654),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_702),
.B(n_673),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_656),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_695),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_652),
.B(n_244),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_683),
.B(n_360),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_634),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_656),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_657),
.B(n_559),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_657),
.B(n_559),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_658),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_672),
.B(n_246),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_658),
.B(n_529),
.Y(n_853)
);

NAND2x1_ASAP7_75t_L g854 ( 
.A(n_570),
.B(n_498),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_662),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_660),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_708),
.B(n_247),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_660),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_648),
.A2(n_224),
.B(n_334),
.C(n_227),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_686),
.B(n_251),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_634),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_634),
.A2(n_354),
.B1(n_227),
.B2(n_240),
.Y(n_862)
);

NAND2xp33_ASAP7_75t_L g863 ( 
.A(n_653),
.B(n_357),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_628),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_663),
.B(n_529),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_663),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_674),
.B(n_676),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_674),
.B(n_483),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_704),
.B(n_254),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_706),
.B(n_261),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_634),
.A2(n_258),
.B1(n_240),
.B2(n_245),
.Y(n_871)
);

BUFx6f_ASAP7_75t_SL g872 ( 
.A(n_662),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_676),
.B(n_483),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_682),
.B(n_483),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_566),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_682),
.B(n_488),
.Y(n_876)
);

NOR2xp67_ASAP7_75t_SL g877 ( 
.A(n_635),
.B(n_200),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_648),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_662),
.B(n_245),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_685),
.Y(n_880)
);

NOR2xp67_ASAP7_75t_L g881 ( 
.A(n_568),
.B(n_75),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_685),
.B(n_488),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_592),
.B(n_263),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_677),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_568),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_725),
.B(n_692),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_714),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_724),
.B(n_592),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_751),
.B(n_661),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_715),
.B(n_692),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_751),
.Y(n_891)
);

AO21x1_ASAP7_75t_L g892 ( 
.A1(n_746),
.A2(n_250),
.B(n_249),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_836),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_754),
.A2(n_775),
.B(n_742),
.C(n_883),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_836),
.Y(n_895)
);

INVx5_ASAP7_75t_L g896 ( 
.A(n_836),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_724),
.B(n_677),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_836),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_721),
.A2(n_687),
.B1(n_677),
.B2(n_680),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_723),
.A2(n_687),
.B(n_701),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_764),
.B(n_696),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_764),
.B(n_767),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_878),
.A2(n_687),
.B(n_566),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_767),
.B(n_696),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_722),
.B(n_699),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_730),
.B(n_699),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_729),
.B(n_703),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_878),
.A2(n_566),
.B(n_635),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_769),
.A2(n_731),
.B(n_785),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_842),
.B(n_703),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_727),
.B(n_842),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_778),
.B(n_707),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_884),
.A2(n_712),
.B(n_710),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_884),
.A2(n_566),
.B(n_647),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_750),
.A2(n_828),
.B(n_820),
.C(n_844),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_729),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_836),
.Y(n_917)
);

AOI21xp33_ASAP7_75t_L g918 ( 
.A1(n_795),
.A2(n_869),
.B(n_860),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_867),
.A2(n_778),
.B(n_809),
.C(n_781),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_781),
.B(n_707),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_809),
.B(n_811),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_811),
.B(n_710),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_SL g923 ( 
.A(n_814),
.B(n_680),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_812),
.A2(n_647),
.B(n_651),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_772),
.A2(n_647),
.B(n_651),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_870),
.A2(n_712),
.B(n_711),
.C(n_249),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_720),
.A2(n_711),
.B(n_662),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_741),
.A2(n_647),
.B(n_651),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_720),
.A2(n_573),
.B(n_570),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_813),
.A2(n_818),
.B(n_848),
.C(n_843),
.Y(n_930)
);

BUFx8_ASAP7_75t_L g931 ( 
.A(n_872),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_741),
.A2(n_647),
.B(n_651),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_813),
.B(n_695),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_818),
.B(n_843),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_797),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_838),
.A2(n_250),
.B(n_299),
.C(n_305),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_741),
.A2(n_792),
.B(n_847),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_779),
.B(n_625),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_848),
.B(n_570),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_779),
.B(n_805),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_805),
.B(n_659),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_733),
.B(n_691),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_744),
.A2(n_573),
.B(n_570),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_749),
.A2(n_585),
.B(n_573),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_792),
.A2(n_647),
.B(n_651),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_845),
.A2(n_385),
.B(n_305),
.C(n_311),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_792),
.A2(n_585),
.B(n_573),
.Y(n_947)
);

AOI21xp33_ASAP7_75t_L g948 ( 
.A1(n_852),
.A2(n_705),
.B(n_311),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_797),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_847),
.A2(n_861),
.B(n_755),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_L g951 ( 
.A(n_797),
.B(n_653),
.Y(n_951)
);

BUFx4f_ASAP7_75t_L g952 ( 
.A(n_719),
.Y(n_952)
);

OAI21xp33_ASAP7_75t_L g953 ( 
.A1(n_732),
.A2(n_857),
.B(n_745),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_861),
.A2(n_591),
.B(n_585),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_728),
.A2(n_591),
.B(n_585),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_SL g956 ( 
.A1(n_859),
.A2(n_591),
.B(n_615),
.C(n_604),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_728),
.A2(n_604),
.B(n_591),
.Y(n_957)
);

AND2x2_ASAP7_75t_SL g958 ( 
.A(n_739),
.B(n_200),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_762),
.A2(n_600),
.B(n_597),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_726),
.A2(n_653),
.B1(n_378),
.B2(n_332),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_755),
.A2(n_615),
.B(n_604),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_780),
.B(n_360),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_866),
.B(n_880),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_740),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_727),
.B(n_360),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_718),
.B(n_604),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_866),
.B(n_880),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_717),
.B(n_480),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_726),
.A2(n_698),
.B(n_694),
.C(n_693),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_801),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_826),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_853),
.B(n_615),
.Y(n_972)
);

AO21x2_ASAP7_75t_L g973 ( 
.A1(n_753),
.A2(n_600),
.B(n_597),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_761),
.A2(n_615),
.B(n_626),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_738),
.B(n_267),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_735),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_735),
.Y(n_977)
);

O2A1O1Ixp5_ASAP7_75t_L g978 ( 
.A1(n_760),
.A2(n_698),
.B(n_694),
.C(n_693),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_865),
.B(n_626),
.Y(n_979)
);

CKINVDCx10_ASAP7_75t_R g980 ( 
.A(n_716),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_885),
.B(n_272),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_825),
.B(n_317),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_743),
.A2(n_688),
.B(n_626),
.C(n_667),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_760),
.B(n_626),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_763),
.B(n_667),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_763),
.B(n_667),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_864),
.B(n_279),
.Y(n_987)
);

AO21x1_ASAP7_75t_L g988 ( 
.A1(n_739),
.A2(n_350),
.B(n_347),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_776),
.A2(n_640),
.B(n_636),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_784),
.B(n_667),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_747),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_784),
.B(n_670),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_747),
.A2(n_688),
.B(n_670),
.C(n_678),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_793),
.B(n_670),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_793),
.B(n_670),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_761),
.A2(n_688),
.B(n_640),
.Y(n_996)
);

OAI321xp33_ASAP7_75t_L g997 ( 
.A1(n_807),
.A2(n_374),
.A3(n_382),
.B1(n_347),
.B2(n_350),
.C(n_353),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_797),
.B(n_317),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_806),
.B(n_688),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_797),
.B(n_480),
.Y(n_1000)
);

NAND2xp33_ASAP7_75t_L g1001 ( 
.A(n_864),
.B(n_653),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_753),
.A2(n_681),
.B(n_678),
.C(n_671),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_759),
.B(n_280),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_817),
.B(n_325),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_804),
.A2(n_681),
.B(n_671),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_806),
.B(n_636),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_810),
.B(n_645),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_804),
.A2(n_664),
.B(n_645),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_787),
.B(n_325),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_748),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_766),
.A2(n_664),
.B(n_646),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_810),
.B(n_646),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_748),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_719),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_855),
.B(n_770),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_823),
.B(n_282),
.Y(n_1016)
);

INVxp67_ASAP7_75t_SL g1017 ( 
.A(n_770),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_771),
.B(n_284),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_770),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_752),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_855),
.A2(n_650),
.B1(n_608),
.B2(n_637),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_827),
.B(n_650),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_827),
.B(n_829),
.Y(n_1023)
);

AND2x6_ASAP7_75t_L g1024 ( 
.A(n_879),
.B(n_317),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_766),
.A2(n_582),
.B(n_567),
.Y(n_1025)
);

AO21x1_ASAP7_75t_L g1026 ( 
.A1(n_821),
.A2(n_366),
.B(n_353),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_752),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_768),
.A2(n_799),
.B(n_783),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_829),
.B(n_653),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_768),
.A2(n_582),
.B(n_567),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_830),
.B(n_608),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_799),
.A2(n_637),
.B(n_629),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_773),
.B(n_293),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_734),
.A2(n_637),
.B1(n_629),
.B2(n_608),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_788),
.A2(n_816),
.B(n_790),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_830),
.B(n_629),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_833),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_757),
.B(n_366),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_756),
.A2(n_561),
.B(n_493),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_719),
.A2(n_561),
.B1(n_317),
.B2(n_369),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_719),
.A2(n_561),
.B1(n_317),
.B2(n_368),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_833),
.B(n_357),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_841),
.B(n_851),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_819),
.A2(n_495),
.B(n_488),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_868),
.A2(n_494),
.B(n_493),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_774),
.B(n_294),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_841),
.B(n_357),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_882),
.A2(n_493),
.B(n_494),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_786),
.B(n_378),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_851),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_873),
.A2(n_876),
.B(n_874),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_832),
.B(n_325),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_824),
.A2(n_494),
.B(n_495),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_879),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_856),
.B(n_496),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_789),
.A2(n_498),
.B1(n_357),
.B2(n_497),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_756),
.A2(n_495),
.B(n_496),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_856),
.B(n_496),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_858),
.B(n_357),
.Y(n_1059)
);

O2A1O1Ixp5_ASAP7_75t_L g1060 ( 
.A1(n_858),
.A2(n_777),
.B(n_782),
.C(n_837),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_758),
.B(n_497),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_834),
.A2(n_497),
.B(n_555),
.Y(n_1062)
);

AOI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_794),
.A2(n_318),
.B(n_314),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_815),
.B(n_297),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_758),
.B(n_504),
.Y(n_1065)
);

O2A1O1Ixp5_ASAP7_75t_L g1066 ( 
.A1(n_840),
.A2(n_468),
.B(n_469),
.C(n_382),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_849),
.A2(n_498),
.B(n_306),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_758),
.B(n_504),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_822),
.B(n_512),
.Y(n_1069)
);

NAND2xp33_ASAP7_75t_L g1070 ( 
.A(n_796),
.B(n_737),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_850),
.A2(n_532),
.B(n_521),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_875),
.A2(n_532),
.B(n_521),
.Y(n_1072)
);

AO21x1_ASAP7_75t_L g1073 ( 
.A1(n_821),
.A2(n_468),
.B(n_469),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_822),
.A2(n_498),
.B1(n_357),
.B2(n_521),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_887),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_940),
.B(n_881),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_911),
.B(n_803),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_918),
.A2(n_879),
.B(n_822),
.C(n_846),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_942),
.A2(n_839),
.B1(n_872),
.B2(n_798),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_894),
.A2(n_765),
.B1(n_872),
.B2(n_808),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_891),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_935),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_896),
.A2(n_875),
.B(n_863),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_R g1084 ( 
.A(n_923),
.B(n_839),
.Y(n_1084)
);

OAI22x1_ASAP7_75t_L g1085 ( 
.A1(n_975),
.A2(n_835),
.B1(n_736),
.B2(n_791),
.Y(n_1085)
);

O2A1O1Ixp5_ASAP7_75t_L g1086 ( 
.A1(n_942),
.A2(n_875),
.B(n_877),
.C(n_854),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_896),
.A2(n_863),
.B(n_802),
.Y(n_1087)
);

OR2x6_ASAP7_75t_L g1088 ( 
.A(n_911),
.B(n_831),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_948),
.A2(n_800),
.B(n_862),
.C(n_871),
.Y(n_1089)
);

O2A1O1Ixp5_ASAP7_75t_L g1090 ( 
.A1(n_906),
.A2(n_877),
.B(n_854),
.C(n_835),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_886),
.B(n_831),
.Y(n_1091)
);

O2A1O1Ixp5_ASAP7_75t_L g1092 ( 
.A1(n_906),
.A2(n_831),
.B(n_802),
.C(n_737),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_893),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_953),
.A2(n_348),
.B(n_308),
.C(n_309),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_935),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_915),
.A2(n_372),
.B(n_310),
.C(n_322),
.Y(n_1096)
);

NOR2x1_ASAP7_75t_L g1097 ( 
.A(n_970),
.B(n_512),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_902),
.B(n_831),
.Y(n_1098)
);

AOI22x1_ASAP7_75t_L g1099 ( 
.A1(n_1051),
.A2(n_802),
.B1(n_737),
.B2(n_373),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_SL g1100 ( 
.A1(n_1018),
.A2(n_498),
.B(n_79),
.C(n_164),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_905),
.B(n_301),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_893),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_941),
.B(n_910),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_896),
.A2(n_535),
.B(n_532),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_889),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_L g1106 ( 
.A(n_976),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_SL g1107 ( 
.A(n_896),
.B(n_327),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_SL g1108 ( 
.A1(n_975),
.A2(n_379),
.B1(n_377),
.B2(n_376),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_904),
.B(n_328),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_900),
.A2(n_535),
.B(n_532),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_899),
.A2(n_535),
.B(n_532),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_971),
.A2(n_938),
.B1(n_1033),
.B2(n_1018),
.Y(n_1112)
);

INVx6_ASAP7_75t_L g1113 ( 
.A(n_931),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_L g1114 ( 
.A(n_1015),
.B(n_512),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_SL g1115 ( 
.A1(n_1016),
.A2(n_375),
.B1(n_363),
.B2(n_343),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_913),
.A2(n_535),
.B(n_532),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_1003),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_890),
.A2(n_903),
.B(n_1070),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_1033),
.A2(n_498),
.B(n_134),
.C(n_120),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1054),
.B(n_108),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_901),
.B(n_341),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_933),
.B(n_339),
.Y(n_1122)
);

INVxp67_ASAP7_75t_SL g1123 ( 
.A(n_1017),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_979),
.A2(n_535),
.B(n_532),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1017),
.B(n_333),
.Y(n_1125)
);

NOR3xp33_ASAP7_75t_L g1126 ( 
.A(n_987),
.B(n_331),
.C(n_329),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_916),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_972),
.A2(n_535),
.B(n_521),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_L g1129 ( 
.A(n_897),
.B(n_535),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_SL g1130 ( 
.A1(n_1046),
.A2(n_179),
.B(n_174),
.C(n_160),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_935),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_987),
.B(n_5),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_916),
.B(n_7),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1000),
.B(n_521),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_971),
.B(n_888),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_952),
.B(n_521),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_909),
.A2(n_521),
.B(n_512),
.Y(n_1137)
);

AO22x1_ASAP7_75t_L g1138 ( 
.A1(n_1016),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_921),
.B(n_512),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_SL g1140 ( 
.A1(n_977),
.A2(n_15),
.B1(n_21),
.B2(n_23),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1019),
.A2(n_512),
.B(n_159),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1019),
.A2(n_512),
.B(n_148),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_934),
.B(n_143),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1020),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1046),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1014),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_952),
.B(n_101),
.Y(n_1147)
);

CKINVDCx14_ASAP7_75t_R g1148 ( 
.A(n_1009),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_946),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1060),
.A2(n_100),
.B(n_99),
.Y(n_1150)
);

AOI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_997),
.A2(n_32),
.B(n_33),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_968),
.B(n_98),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_935),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_943),
.A2(n_94),
.B(n_92),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_944),
.A2(n_90),
.B(n_83),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_951),
.A2(n_78),
.B(n_36),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1000),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_964),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_927),
.A2(n_35),
.B(n_37),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_958),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_966),
.B(n_42),
.Y(n_1161)
);

NAND2x1p5_ASAP7_75t_L g1162 ( 
.A(n_949),
.B(n_45),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_936),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_949),
.B(n_46),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1050),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_R g1166 ( 
.A(n_980),
.B(n_74),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1028),
.A2(n_74),
.B(n_50),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1004),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_931),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_966),
.B(n_49),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1010),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_963),
.B(n_49),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_967),
.B(n_912),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1064),
.A2(n_51),
.B(n_52),
.C(n_56),
.Y(n_1174)
);

O2A1O1Ixp5_ASAP7_75t_L g1175 ( 
.A1(n_982),
.A2(n_51),
.B(n_58),
.C(n_60),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1038),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_965),
.A2(n_58),
.B(n_60),
.C(n_63),
.Y(n_1177)
);

INVx5_ASAP7_75t_L g1178 ( 
.A(n_893),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1050),
.Y(n_1179)
);

OR2x6_ASAP7_75t_L g1180 ( 
.A(n_949),
.B(n_63),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_958),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1064),
.A2(n_70),
.B1(n_1052),
.B2(n_981),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_960),
.A2(n_922),
.B1(n_920),
.B2(n_1023),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1027),
.B(n_70),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_949),
.B(n_1001),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_929),
.A2(n_1043),
.B(n_1068),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1065),
.A2(n_937),
.B(n_1035),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1045),
.A2(n_1044),
.B(n_978),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_893),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1063),
.B(n_919),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1038),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_895),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1049),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_895),
.Y(n_1194)
);

NOR3xp33_ASAP7_75t_SL g1195 ( 
.A(n_981),
.B(n_962),
.C(n_907),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_925),
.A2(n_1069),
.B(n_1039),
.Y(n_1196)
);

AOI221xp5_ASAP7_75t_L g1197 ( 
.A1(n_1049),
.A2(n_960),
.B1(n_892),
.B2(n_930),
.C(n_926),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1061),
.A2(n_1029),
.B(n_1057),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_950),
.A2(n_986),
.B(n_984),
.Y(n_1199)
);

INVx5_ASAP7_75t_L g1200 ( 
.A(n_895),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_991),
.B(n_1013),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1040),
.A2(n_1041),
.B(n_983),
.C(n_993),
.Y(n_1202)
);

BUFx12f_ASAP7_75t_L g1203 ( 
.A(n_1024),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1037),
.B(n_939),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_985),
.A2(n_990),
.B(n_995),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_895),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_978),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1055),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_898),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1006),
.B(n_1022),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_988),
.B(n_1026),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1058),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1007),
.B(n_1012),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_992),
.A2(n_999),
.B(n_994),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_898),
.B(n_917),
.Y(n_1215)
);

BUFx4f_ASAP7_75t_L g1216 ( 
.A(n_898),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_973),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_898),
.B(n_917),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1021),
.A2(n_1047),
.B(n_1059),
.C(n_1042),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1031),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1036),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_908),
.A2(n_914),
.B(n_1060),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_917),
.B(n_973),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_SL g1224 ( 
.A(n_917),
.B(n_1024),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_956),
.A2(n_998),
.B(n_1002),
.C(n_1066),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1067),
.B(n_1066),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1034),
.Y(n_1227)
);

BUFx12f_ASAP7_75t_L g1228 ( 
.A(n_1024),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1011),
.B(n_1032),
.Y(n_1229)
);

NOR3xp33_ASAP7_75t_SL g1230 ( 
.A(n_974),
.B(n_961),
.C(n_955),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_996),
.A2(n_947),
.B(n_954),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_969),
.A2(n_1073),
.B(n_1025),
.C(n_1030),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1005),
.B(n_1008),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_928),
.A2(n_932),
.B(n_945),
.Y(n_1234)
);

AOI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1111),
.A2(n_1222),
.B(n_1118),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1187),
.A2(n_957),
.B(n_924),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1075),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1217),
.A2(n_1071),
.A3(n_1062),
.B(n_1048),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1112),
.B(n_1024),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_L g1240 ( 
.A(n_1182),
.B(n_1074),
.C(n_1053),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1223),
.A2(n_1072),
.A3(n_989),
.B(n_959),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_SL g1242 ( 
.A1(n_1078),
.A2(n_1056),
.B(n_1024),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1132),
.A2(n_1135),
.B1(n_1145),
.B2(n_1103),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1117),
.B(n_1076),
.Y(n_1244)
);

AO22x2_ASAP7_75t_L g1245 ( 
.A1(n_1160),
.A2(n_1181),
.B1(n_1159),
.B2(n_1170),
.Y(n_1245)
);

INVx5_ASAP7_75t_SL g1246 ( 
.A(n_1180),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1168),
.B(n_1101),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1089),
.A2(n_1195),
.B(n_1080),
.C(n_1096),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1190),
.A2(n_1197),
.B(n_1173),
.C(n_1155),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1173),
.B(n_1109),
.Y(n_1250)
);

INVx8_ASAP7_75t_L g1251 ( 
.A(n_1178),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1216),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1205),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1147),
.A2(n_1181),
.B(n_1160),
.C(n_1130),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1188),
.A2(n_1110),
.B(n_1234),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1199),
.A2(n_1231),
.B(n_1214),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1127),
.B(n_1081),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1191),
.B(n_1121),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1196),
.A2(n_1207),
.A3(n_1183),
.B(n_1229),
.Y(n_1259)
);

AO22x2_ASAP7_75t_L g1260 ( 
.A1(n_1161),
.A2(n_1150),
.B1(n_1091),
.B2(n_1098),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1106),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1150),
.A2(n_1226),
.B(n_1086),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1210),
.A2(n_1213),
.B(n_1087),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_1183),
.A2(n_1154),
.A3(n_1116),
.B(n_1091),
.Y(n_1264)
);

OAI21xp33_ASAP7_75t_L g1265 ( 
.A1(n_1126),
.A2(n_1133),
.B(n_1174),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1079),
.A2(n_1123),
.B1(n_1180),
.B2(n_1088),
.Y(n_1266)
);

AOI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1233),
.A2(n_1139),
.B(n_1143),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1124),
.A2(n_1128),
.B(n_1083),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1216),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1137),
.A2(n_1232),
.B(n_1143),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1122),
.B(n_1176),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_1146),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1137),
.A2(n_1139),
.B(n_1202),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1204),
.A2(n_1219),
.B(n_1225),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1148),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1104),
.A2(n_1129),
.B(n_1099),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1158),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1092),
.A2(n_1090),
.B(n_1098),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1204),
.A2(n_1178),
.B(n_1200),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1178),
.A2(n_1200),
.B(n_1220),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1113),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1178),
.A2(n_1200),
.B(n_1221),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1200),
.A2(n_1136),
.B(n_1134),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1085),
.A2(n_1184),
.A3(n_1172),
.B(n_1167),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1208),
.B(n_1212),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1180),
.A2(n_1088),
.B1(n_1172),
.B2(n_1171),
.Y(n_1286)
);

NOR2x1_ASAP7_75t_SL g1287 ( 
.A(n_1088),
.B(n_1192),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1108),
.A2(n_1115),
.B1(n_1140),
.B2(n_1084),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1211),
.A2(n_1230),
.B(n_1227),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1106),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1224),
.A2(n_1141),
.B(n_1142),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1120),
.B(n_1193),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1177),
.A2(n_1094),
.B(n_1149),
.C(n_1163),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1114),
.A2(n_1215),
.B(n_1201),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1184),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1152),
.A2(n_1156),
.B(n_1125),
.Y(n_1296)
);

NAND3x1_ASAP7_75t_L g1297 ( 
.A(n_1077),
.B(n_1097),
.C(n_1138),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1144),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1151),
.A2(n_1175),
.B(n_1157),
.C(n_1100),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1113),
.A2(n_1169),
.B1(n_1164),
.B2(n_1162),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1151),
.A2(n_1120),
.B(n_1179),
.C(n_1165),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1209),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1093),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1162),
.B(n_1164),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1218),
.B(n_1185),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1107),
.A2(n_1119),
.B(n_1082),
.C(n_1095),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1218),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1113),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1095),
.B(n_1153),
.Y(n_1309)
);

AO21x1_ASAP7_75t_L g1310 ( 
.A1(n_1131),
.A2(n_1192),
.B(n_1153),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_SL g1311 ( 
.A1(n_1206),
.A2(n_1228),
.B(n_1203),
.C(n_1131),
.Y(n_1311)
);

AOI21xp33_ASAP7_75t_L g1312 ( 
.A1(n_1093),
.A2(n_1102),
.B(n_1189),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1093),
.A2(n_1102),
.A3(n_1189),
.B(n_1194),
.Y(n_1313)
);

INVxp33_ASAP7_75t_L g1314 ( 
.A(n_1166),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1102),
.A2(n_1189),
.B(n_1194),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1081),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1118),
.A2(n_755),
.B(n_728),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1218),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1112),
.B(n_722),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1186),
.A2(n_894),
.B(n_1198),
.Y(n_1320)
);

OA22x2_ASAP7_75t_L g1321 ( 
.A1(n_1145),
.A2(n_592),
.B1(n_1140),
.B2(n_1112),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1123),
.Y(n_1322)
);

AOI22x1_ASAP7_75t_L g1323 ( 
.A1(n_1085),
.A2(n_1159),
.B1(n_1118),
.B2(n_1155),
.Y(n_1323)
);

AOI221x1_ASAP7_75t_L g1324 ( 
.A1(n_1159),
.A2(n_918),
.B1(n_894),
.B2(n_1150),
.C(n_1160),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1188),
.A2(n_1045),
.B(n_1110),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1186),
.A2(n_894),
.B(n_1198),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1118),
.A2(n_755),
.B(n_728),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1188),
.A2(n_1045),
.B(n_1110),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1105),
.B(n_889),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1081),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1103),
.B(n_940),
.Y(n_1331)
);

AOI221xp5_ASAP7_75t_L g1332 ( 
.A1(n_1182),
.A2(n_746),
.B1(n_883),
.B2(n_975),
.C(n_564),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1103),
.B(n_940),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1103),
.B(n_940),
.Y(n_1334)
);

NAND3x1_ASAP7_75t_L g1335 ( 
.A(n_1132),
.B(n_883),
.C(n_746),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1118),
.A2(n_755),
.B(n_728),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1222),
.A2(n_1217),
.A3(n_769),
.B(n_731),
.Y(n_1337)
);

AOI211x1_ASAP7_75t_L g1338 ( 
.A1(n_1138),
.A2(n_1151),
.B(n_1103),
.C(n_1160),
.Y(n_1338)
);

AO32x2_ASAP7_75t_L g1339 ( 
.A1(n_1160),
.A2(n_1181),
.A3(n_1145),
.B1(n_1183),
.B2(n_1140),
.Y(n_1339)
);

AOI221x1_ASAP7_75t_L g1340 ( 
.A1(n_1159),
.A2(n_918),
.B1(n_894),
.B2(n_1150),
.C(n_1160),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1118),
.A2(n_755),
.B(n_728),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1173),
.A2(n_894),
.B1(n_958),
.B2(n_942),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1118),
.A2(n_755),
.B(n_728),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1188),
.A2(n_1045),
.B(n_1110),
.Y(n_1344)
);

NOR2xp67_ASAP7_75t_L g1345 ( 
.A(n_1080),
.B(n_886),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_SL g1346 ( 
.A1(n_1159),
.A2(n_930),
.B(n_988),
.Y(n_1346)
);

AO31x2_ASAP7_75t_L g1347 ( 
.A1(n_1222),
.A2(n_1217),
.A3(n_769),
.B(n_731),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1112),
.B(n_722),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1186),
.A2(n_894),
.B(n_1198),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1105),
.B(n_889),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1188),
.A2(n_1045),
.B(n_1110),
.Y(n_1351)
);

AO31x2_ASAP7_75t_L g1352 ( 
.A1(n_1222),
.A2(n_1217),
.A3(n_769),
.B(n_731),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1186),
.A2(n_894),
.B(n_1198),
.Y(n_1353)
);

O2A1O1Ixp5_ASAP7_75t_L g1354 ( 
.A1(n_1190),
.A2(n_918),
.B(n_894),
.C(n_942),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1103),
.B(n_940),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1105),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1186),
.A2(n_894),
.B(n_1198),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1150),
.A2(n_1188),
.B(n_1137),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1188),
.A2(n_1045),
.B(n_1110),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1112),
.A2(n_814),
.B1(n_586),
.B2(n_746),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1222),
.A2(n_1217),
.A3(n_769),
.B(n_731),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1188),
.A2(n_1045),
.B(n_1110),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1188),
.A2(n_1045),
.B(n_1110),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_SL g1364 ( 
.A(n_1160),
.B(n_839),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_SL g1365 ( 
.A1(n_1078),
.A2(n_894),
.B(n_918),
.C(n_1096),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1105),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1076),
.B(n_976),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1120),
.B(n_911),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1188),
.A2(n_1045),
.B(n_1110),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1076),
.B(n_976),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1113),
.Y(n_1371)
);

AO31x2_ASAP7_75t_L g1372 ( 
.A1(n_1222),
.A2(n_1217),
.A3(n_769),
.B(n_731),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1081),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1188),
.A2(n_1045),
.B(n_1110),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1118),
.A2(n_755),
.B(n_728),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1118),
.A2(n_755),
.B(n_728),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1112),
.B(n_722),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1103),
.B(n_940),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_SL g1379 ( 
.A(n_1182),
.B(n_746),
.C(n_894),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1112),
.B(n_722),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1188),
.A2(n_1045),
.B(n_1110),
.Y(n_1381)
);

AO31x2_ASAP7_75t_L g1382 ( 
.A1(n_1222),
.A2(n_1217),
.A3(n_769),
.B(n_731),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1118),
.A2(n_755),
.B(n_728),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1081),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1112),
.B(n_722),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1105),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1222),
.A2(n_1217),
.A3(n_769),
.B(n_731),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1118),
.A2(n_755),
.B(n_728),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1319),
.A2(n_1377),
.B1(n_1380),
.B2(n_1348),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1366),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1277),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1332),
.A2(n_1288),
.B(n_1385),
.Y(n_1392)
);

AOI21xp33_ASAP7_75t_L g1393 ( 
.A1(n_1335),
.A2(n_1265),
.B(n_1360),
.Y(n_1393)
);

INVx8_ASAP7_75t_L g1394 ( 
.A(n_1251),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1379),
.A2(n_1321),
.B1(n_1265),
.B2(n_1245),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1371),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1281),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1250),
.B(n_1331),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1364),
.A2(n_1246),
.B1(n_1245),
.B2(n_1266),
.Y(n_1399)
);

BUFx10_ASAP7_75t_L g1400 ( 
.A(n_1257),
.Y(n_1400)
);

BUFx12f_ASAP7_75t_L g1401 ( 
.A(n_1275),
.Y(n_1401)
);

BUFx2_ASAP7_75t_SL g1402 ( 
.A(n_1316),
.Y(n_1402)
);

CKINVDCx11_ASAP7_75t_R g1403 ( 
.A(n_1290),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1251),
.Y(n_1404)
);

BUFx2_ASAP7_75t_SL g1405 ( 
.A(n_1330),
.Y(n_1405)
);

BUFx8_ASAP7_75t_SL g1406 ( 
.A(n_1386),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1252),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1243),
.A2(n_1258),
.B1(n_1271),
.B2(n_1244),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1252),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1243),
.A2(n_1342),
.B1(n_1345),
.B2(n_1295),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1342),
.A2(n_1345),
.B1(n_1364),
.B2(n_1239),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1333),
.A2(n_1334),
.B1(n_1355),
.B2(n_1378),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1323),
.A2(n_1266),
.B1(n_1260),
.B2(n_1289),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1246),
.A2(n_1286),
.B1(n_1247),
.B2(n_1367),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1260),
.A2(n_1289),
.B1(n_1240),
.B2(n_1286),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1373),
.Y(n_1416)
);

BUFx12f_ASAP7_75t_L g1417 ( 
.A(n_1261),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1248),
.A2(n_1322),
.B1(n_1249),
.B2(n_1356),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1370),
.A2(n_1368),
.B1(n_1292),
.B2(n_1300),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1259),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1324),
.A2(n_1340),
.B(n_1293),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1252),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1384),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1269),
.Y(n_1424)
);

AND2x4_ASAP7_75t_SL g1425 ( 
.A(n_1269),
.B(n_1368),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1259),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1240),
.A2(n_1270),
.B1(n_1285),
.B2(n_1339),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1308),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1259),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1339),
.A2(n_1287),
.B1(n_1304),
.B2(n_1281),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1298),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1297),
.A2(n_1365),
.B1(n_1272),
.B2(n_1305),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1339),
.A2(n_1346),
.B1(n_1357),
.B2(n_1326),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1302),
.B(n_1338),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1309),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1274),
.A2(n_1273),
.B1(n_1320),
.B2(n_1326),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1320),
.A2(n_1349),
.B1(n_1357),
.B2(n_1353),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1349),
.A2(n_1353),
.B1(n_1262),
.B2(n_1296),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1338),
.B(n_1307),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1269),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1318),
.B(n_1315),
.Y(n_1441)
);

OAI21xp33_ASAP7_75t_L g1442 ( 
.A1(n_1301),
.A2(n_1314),
.B(n_1262),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1303),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1313),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1278),
.A2(n_1263),
.B1(n_1291),
.B2(n_1358),
.Y(n_1445)
);

BUFx10_ASAP7_75t_L g1446 ( 
.A(n_1303),
.Y(n_1446)
);

INVx6_ASAP7_75t_L g1447 ( 
.A(n_1311),
.Y(n_1447)
);

INVx6_ASAP7_75t_L g1448 ( 
.A(n_1312),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1284),
.B(n_1354),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1313),
.Y(n_1450)
);

INVxp67_ASAP7_75t_SL g1451 ( 
.A(n_1310),
.Y(n_1451)
);

BUFx12f_ASAP7_75t_L g1452 ( 
.A(n_1313),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1283),
.A2(n_1282),
.B1(n_1280),
.B2(n_1279),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1294),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1278),
.A2(n_1358),
.B1(n_1253),
.B2(n_1254),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1306),
.A2(n_1253),
.B1(n_1388),
.B2(n_1383),
.Y(n_1456)
);

BUFx12f_ASAP7_75t_L g1457 ( 
.A(n_1284),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1315),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1317),
.A2(n_1341),
.B1(n_1343),
.B2(n_1376),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1284),
.B(n_1264),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1337),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1327),
.A2(n_1375),
.B1(n_1336),
.B2(n_1267),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1299),
.A2(n_1242),
.B1(n_1236),
.B2(n_1235),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_SL g1464 ( 
.A1(n_1256),
.A2(n_1276),
.B1(n_1268),
.B2(n_1255),
.Y(n_1464)
);

CKINVDCx11_ASAP7_75t_R g1465 ( 
.A(n_1264),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1325),
.A2(n_1359),
.B1(n_1381),
.B2(n_1362),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1328),
.A2(n_1374),
.B1(n_1369),
.B2(n_1344),
.Y(n_1467)
);

NAND2x1p5_ASAP7_75t_L g1468 ( 
.A(n_1351),
.B(n_1363),
.Y(n_1468)
);

CKINVDCx8_ASAP7_75t_R g1469 ( 
.A(n_1264),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1347),
.A2(n_1352),
.B1(n_1361),
.B2(n_1372),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1241),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1352),
.A2(n_1361),
.B1(n_1372),
.B2(n_1382),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1361),
.A2(n_1387),
.B1(n_1372),
.B2(n_1382),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1241),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1387),
.Y(n_1475)
);

INVx8_ASAP7_75t_L g1476 ( 
.A(n_1238),
.Y(n_1476)
);

CKINVDCx6p67_ASAP7_75t_R g1477 ( 
.A(n_1238),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1367),
.B(n_1370),
.Y(n_1478)
);

BUFx8_ASAP7_75t_SL g1479 ( 
.A(n_1371),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1480)
);

BUFx4f_ASAP7_75t_SL g1481 ( 
.A(n_1371),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1367),
.B(n_1370),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1485)
);

CKINVDCx11_ASAP7_75t_R g1486 ( 
.A(n_1371),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1366),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1319),
.A2(n_1377),
.B1(n_1380),
.B2(n_1348),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1489)
);

OAI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1321),
.A2(n_1243),
.B1(n_1332),
.B2(n_1319),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1316),
.Y(n_1493)
);

INVx8_ASAP7_75t_L g1494 ( 
.A(n_1251),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1251),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1366),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1498)
);

CKINVDCx6p67_ASAP7_75t_R g1499 ( 
.A(n_1371),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1319),
.A2(n_1377),
.B1(n_1380),
.B2(n_1348),
.Y(n_1500)
);

BUFx12f_ASAP7_75t_L g1501 ( 
.A(n_1275),
.Y(n_1501)
);

BUFx12f_ASAP7_75t_L g1502 ( 
.A(n_1275),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1329),
.B(n_1350),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1316),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1237),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1319),
.A2(n_1377),
.B1(n_1380),
.B2(n_1348),
.Y(n_1506)
);

INVx6_ASAP7_75t_L g1507 ( 
.A(n_1252),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1319),
.A2(n_894),
.B(n_918),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1366),
.Y(n_1510)
);

CKINVDCx11_ASAP7_75t_R g1511 ( 
.A(n_1371),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1237),
.Y(n_1512)
);

AO22x1_ASAP7_75t_L g1513 ( 
.A1(n_1319),
.A2(n_1348),
.B1(n_1380),
.B2(n_1377),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1319),
.A2(n_894),
.B(n_918),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1332),
.A2(n_1385),
.B1(n_1380),
.B2(n_1319),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1452),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1461),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1475),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1474),
.B(n_1449),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1454),
.B(n_1441),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1444),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1448),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1450),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1448),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1421),
.A2(n_1455),
.B(n_1413),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1433),
.B(n_1460),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1458),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1395),
.B(n_1415),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1420),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1452),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1426),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1457),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1429),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1513),
.B(n_1389),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1471),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1471),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1457),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1469),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1488),
.A2(n_1500),
.B1(n_1506),
.B2(n_1490),
.C(n_1392),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1477),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1498),
.B(n_1508),
.Y(n_1541)
);

AO21x2_ASAP7_75t_L g1542 ( 
.A1(n_1462),
.A2(n_1456),
.B(n_1463),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1476),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1395),
.B(n_1415),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1470),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1472),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1427),
.B(n_1413),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1390),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1468),
.A2(n_1467),
.B(n_1466),
.Y(n_1549)
);

A2O1A1Ixp33_ASAP7_75t_L g1550 ( 
.A1(n_1480),
.A2(n_1515),
.B(n_1482),
.C(n_1484),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1437),
.B(n_1427),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1480),
.B(n_1482),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1503),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1394),
.Y(n_1554)
);

AO21x2_ASAP7_75t_L g1555 ( 
.A1(n_1509),
.A2(n_1514),
.B(n_1453),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1398),
.B(n_1484),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1466),
.A2(n_1467),
.B(n_1459),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1465),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1408),
.B(n_1478),
.Y(n_1559)
);

CKINVDCx6p67_ASAP7_75t_R g1560 ( 
.A(n_1486),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1451),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1394),
.B(n_1494),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1485),
.B(n_1489),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1494),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1439),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1432),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1485),
.A2(n_1515),
.B(n_1497),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1447),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1431),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1473),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1437),
.B(n_1411),
.Y(n_1571)
);

OR2x6_ASAP7_75t_L g1572 ( 
.A(n_1418),
.B(n_1442),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1391),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1495),
.B(n_1505),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1411),
.B(n_1410),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1447),
.B(n_1404),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1512),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1510),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1435),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1455),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1410),
.B(n_1399),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1434),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1447),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1436),
.B(n_1489),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1436),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1483),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1459),
.A2(n_1445),
.B(n_1438),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1464),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1491),
.B(n_1492),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1438),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1491),
.B(n_1492),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1419),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1402),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1445),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1443),
.Y(n_1595)
);

AOI222xp33_ASAP7_75t_L g1596 ( 
.A1(n_1497),
.A2(n_1412),
.B1(n_1481),
.B2(n_1423),
.C1(n_1502),
.C2(n_1501),
.Y(n_1596)
);

NAND4xp25_ASAP7_75t_L g1597 ( 
.A(n_1393),
.B(n_1412),
.C(n_1414),
.D(n_1430),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1527),
.B(n_1400),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1553),
.B(n_1400),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1572),
.B(n_1405),
.Y(n_1600)
);

A2O1A1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1539),
.A2(n_1425),
.B(n_1409),
.C(n_1440),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1567),
.A2(n_1504),
.B1(n_1493),
.B2(n_1397),
.C(n_1416),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1521),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1519),
.B(n_1504),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1519),
.B(n_1493),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1574),
.Y(n_1606)
);

OR2x6_ASAP7_75t_L g1607 ( 
.A(n_1572),
.B(n_1417),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1550),
.A2(n_1481),
.B1(n_1499),
.B2(n_1496),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1541),
.A2(n_1552),
.B1(n_1563),
.B2(n_1591),
.Y(n_1609)
);

NAND4xp25_ASAP7_75t_L g1610 ( 
.A(n_1559),
.B(n_1403),
.C(n_1406),
.D(n_1511),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1589),
.A2(n_1487),
.B(n_1428),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1548),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1522),
.Y(n_1613)
);

CKINVDCx6p67_ASAP7_75t_R g1614 ( 
.A(n_1560),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1565),
.B(n_1409),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1534),
.A2(n_1511),
.B(n_1507),
.C(n_1407),
.Y(n_1616)
);

AO32x2_ASAP7_75t_L g1617 ( 
.A1(n_1524),
.A2(n_1446),
.A3(n_1507),
.B1(n_1407),
.B2(n_1409),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1584),
.A2(n_1396),
.B1(n_1424),
.B2(n_1409),
.C(n_1422),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1558),
.B(n_1422),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1572),
.A2(n_1507),
.B(n_1501),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1586),
.B(n_1401),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1526),
.B(n_1401),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1526),
.B(n_1502),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1520),
.B(n_1479),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1581),
.A2(n_1575),
.B(n_1584),
.C(n_1597),
.Y(n_1625)
);

NAND4xp25_ASAP7_75t_L g1626 ( 
.A(n_1596),
.B(n_1556),
.C(n_1566),
.D(n_1544),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1549),
.A2(n_1557),
.B(n_1587),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1587),
.A2(n_1566),
.B(n_1575),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1592),
.B(n_1582),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1549),
.A2(n_1580),
.B(n_1588),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1595),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1571),
.A2(n_1544),
.B(n_1528),
.Y(n_1632)
);

OAI211xp5_ASAP7_75t_L g1633 ( 
.A1(n_1528),
.A2(n_1581),
.B(n_1547),
.C(n_1525),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1590),
.B(n_1585),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1561),
.Y(n_1635)
);

INVx4_ASAP7_75t_L g1636 ( 
.A(n_1576),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1571),
.A2(n_1585),
.B(n_1590),
.Y(n_1637)
);

OR2x6_ASAP7_75t_L g1638 ( 
.A(n_1532),
.B(n_1543),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1551),
.A2(n_1547),
.B1(n_1525),
.B2(n_1582),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1574),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1582),
.B(n_1555),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1555),
.A2(n_1542),
.B1(n_1537),
.B2(n_1593),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1523),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1555),
.A2(n_1542),
.B1(n_1538),
.B2(n_1595),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1551),
.A2(n_1561),
.B(n_1583),
.C(n_1568),
.Y(n_1645)
);

AO32x2_ASAP7_75t_L g1646 ( 
.A1(n_1580),
.A2(n_1525),
.A3(n_1545),
.B1(n_1546),
.B2(n_1570),
.Y(n_1646)
);

NAND3xp33_ASAP7_75t_L g1647 ( 
.A(n_1525),
.B(n_1588),
.C(n_1540),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1574),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1579),
.B(n_1569),
.Y(n_1649)
);

AO32x2_ASAP7_75t_L g1650 ( 
.A1(n_1545),
.A2(n_1546),
.A3(n_1570),
.B1(n_1523),
.B2(n_1518),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1617),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1628),
.B(n_1594),
.Y(n_1652)
);

OAI222xp33_ASAP7_75t_L g1653 ( 
.A1(n_1609),
.A2(n_1579),
.B1(n_1576),
.B2(n_1577),
.C1(n_1573),
.C2(n_1562),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1630),
.B(n_1594),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1603),
.Y(n_1655)
);

AOI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1609),
.A2(n_1560),
.B1(n_1574),
.B2(n_1568),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1606),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1603),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1617),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1630),
.B(n_1535),
.Y(n_1660)
);

INVx5_ASAP7_75t_L g1661 ( 
.A(n_1600),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1606),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1643),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1641),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1641),
.B(n_1579),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1634),
.B(n_1639),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1639),
.B(n_1536),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1634),
.B(n_1635),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1613),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1649),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1626),
.A2(n_1608),
.B1(n_1607),
.B2(n_1602),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1608),
.A2(n_1540),
.B1(n_1516),
.B2(n_1530),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1627),
.A2(n_1533),
.B(n_1531),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1650),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1638),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1644),
.B(n_1529),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1642),
.B(n_1629),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1647),
.B(n_1517),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1655),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1655),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1658),
.Y(n_1681)
);

AOI33xp33_ASAP7_75t_L g1682 ( 
.A1(n_1671),
.A2(n_1652),
.A3(n_1654),
.B1(n_1599),
.B2(n_1660),
.B3(n_1598),
.Y(n_1682)
);

AOI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1666),
.A2(n_1625),
.B1(n_1632),
.B2(n_1637),
.C(n_1633),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1669),
.Y(n_1684)
);

AOI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1666),
.A2(n_1625),
.B1(n_1633),
.B2(n_1602),
.C(n_1616),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1673),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1677),
.A2(n_1607),
.B1(n_1631),
.B2(n_1620),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1675),
.B(n_1640),
.Y(n_1688)
);

AOI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1677),
.A2(n_1616),
.B(n_1611),
.C(n_1601),
.Y(n_1689)
);

AND2x2_ASAP7_75t_SL g1690 ( 
.A(n_1651),
.B(n_1636),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1664),
.B(n_1629),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1661),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1664),
.B(n_1665),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1656),
.A2(n_1601),
.B1(n_1645),
.B2(n_1618),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1665),
.Y(n_1695)
);

AOI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1652),
.A2(n_1653),
.B1(n_1672),
.B2(n_1651),
.C(n_1659),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1673),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1673),
.Y(n_1698)
);

OR2x2_ASAP7_75t_SL g1699 ( 
.A(n_1651),
.B(n_1604),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1675),
.B(n_1648),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1661),
.Y(n_1701)
);

NOR2x1_ASAP7_75t_L g1702 ( 
.A(n_1678),
.B(n_1645),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1673),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1656),
.A2(n_1618),
.B1(n_1605),
.B2(n_1614),
.Y(n_1704)
);

AOI322xp5_ASAP7_75t_L g1705 ( 
.A1(n_1674),
.A2(n_1623),
.A3(n_1622),
.B1(n_1621),
.B2(n_1624),
.C1(n_1578),
.C2(n_1612),
.Y(n_1705)
);

XNOR2x1_ASAP7_75t_L g1706 ( 
.A(n_1678),
.B(n_1619),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1651),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1657),
.B(n_1646),
.Y(n_1708)
);

INVx4_ASAP7_75t_L g1709 ( 
.A(n_1661),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1669),
.B(n_1610),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1667),
.B(n_1615),
.Y(n_1711)
);

INVxp67_ASAP7_75t_SL g1712 ( 
.A(n_1660),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1676),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1667),
.B(n_1638),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1707),
.B(n_1651),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1707),
.B(n_1651),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1692),
.B(n_1659),
.Y(n_1717)
);

INVx6_ASAP7_75t_L g1718 ( 
.A(n_1692),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1707),
.B(n_1659),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1707),
.B(n_1659),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1686),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1699),
.B(n_1674),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1686),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1713),
.B(n_1670),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1686),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1708),
.B(n_1712),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1708),
.B(n_1659),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1713),
.B(n_1659),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1699),
.B(n_1674),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1697),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1679),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1693),
.B(n_1668),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1702),
.B(n_1654),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1702),
.B(n_1657),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1679),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1680),
.Y(n_1736)
);

INVx4_ASAP7_75t_SL g1737 ( 
.A(n_1680),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1692),
.B(n_1661),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1690),
.B(n_1662),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1695),
.B(n_1668),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1693),
.B(n_1663),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1714),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1697),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1681),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1681),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1733),
.B(n_1682),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1731),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1722),
.B(n_1691),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1739),
.B(n_1690),
.Y(n_1749)
);

INVxp67_ASAP7_75t_L g1750 ( 
.A(n_1733),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1731),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1735),
.Y(n_1752)
);

NOR2x1p5_ASAP7_75t_L g1753 ( 
.A(n_1722),
.B(n_1684),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1733),
.B(n_1683),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1721),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1722),
.B(n_1691),
.Y(n_1756)
);

OAI22xp33_ASAP7_75t_SL g1757 ( 
.A1(n_1718),
.A2(n_1704),
.B1(n_1694),
.B2(n_1701),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1742),
.B(n_1683),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1735),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1736),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1739),
.B(n_1692),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1739),
.B(n_1690),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1727),
.B(n_1688),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1736),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1734),
.A2(n_1696),
.B(n_1685),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1721),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1727),
.B(n_1688),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1721),
.Y(n_1768)
);

INVx2_ASAP7_75t_SL g1769 ( 
.A(n_1718),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1727),
.B(n_1700),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1721),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1728),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1744),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1729),
.B(n_1711),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1744),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1742),
.A2(n_1696),
.B1(n_1685),
.B2(n_1694),
.C(n_1689),
.Y(n_1776)
);

NAND2x1p5_ASAP7_75t_L g1777 ( 
.A(n_1734),
.B(n_1701),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1745),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1723),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1732),
.B(n_1740),
.Y(n_1780)
);

NAND2x1p5_ASAP7_75t_L g1781 ( 
.A(n_1734),
.B(n_1701),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1732),
.B(n_1706),
.Y(n_1782)
);

OAI21xp33_ASAP7_75t_L g1783 ( 
.A1(n_1732),
.A2(n_1705),
.B(n_1689),
.Y(n_1783)
);

OR2x6_ASAP7_75t_L g1784 ( 
.A(n_1718),
.B(n_1701),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1718),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1729),
.B(n_1711),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1745),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1737),
.B(n_1709),
.Y(n_1788)
);

INVxp67_ASAP7_75t_SL g1789 ( 
.A(n_1724),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1718),
.A2(n_1704),
.B1(n_1687),
.B2(n_1706),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1759),
.Y(n_1791)
);

AND2x4_ASAP7_75t_SL g1792 ( 
.A(n_1788),
.B(n_1784),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1749),
.B(n_1715),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1776),
.B(n_1726),
.Y(n_1794)
);

OAI21xp33_ASAP7_75t_L g1795 ( 
.A1(n_1783),
.A2(n_1705),
.B(n_1729),
.Y(n_1795)
);

CKINVDCx16_ASAP7_75t_R g1796 ( 
.A(n_1765),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1759),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1749),
.B(n_1715),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1760),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1755),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1788),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1762),
.B(n_1715),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1760),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1755),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1772),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1766),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1758),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1754),
.B(n_1726),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1773),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1790),
.A2(n_1718),
.B1(n_1738),
.B2(n_1710),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1766),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1750),
.Y(n_1812)
);

INVx3_ASAP7_75t_L g1813 ( 
.A(n_1788),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1768),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1773),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1746),
.A2(n_1706),
.B1(n_1661),
.B2(n_1728),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1775),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1782),
.B(n_1726),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1789),
.B(n_1741),
.Y(n_1819)
);

AOI221xp5_ASAP7_75t_L g1820 ( 
.A1(n_1757),
.A2(n_1728),
.B1(n_1717),
.B2(n_1741),
.C(n_1740),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1775),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1747),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1751),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1780),
.B(n_1724),
.Y(n_1824)
);

OA21x2_ASAP7_75t_L g1825 ( 
.A1(n_1768),
.A2(n_1703),
.B(n_1698),
.Y(n_1825)
);

NOR2x1_ASAP7_75t_L g1826 ( 
.A(n_1753),
.B(n_1717),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1762),
.B(n_1716),
.Y(n_1827)
);

AOI21xp33_ASAP7_75t_L g1828 ( 
.A1(n_1795),
.A2(n_1785),
.B(n_1769),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1791),
.Y(n_1829)
);

AOI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1796),
.A2(n_1795),
.B1(n_1794),
.B2(n_1826),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1796),
.A2(n_1784),
.B1(n_1781),
.B2(n_1777),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1793),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1820),
.B(n_1761),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1794),
.A2(n_1784),
.B(n_1769),
.Y(n_1834)
);

OAI21xp33_ASAP7_75t_L g1835 ( 
.A1(n_1807),
.A2(n_1820),
.B(n_1810),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1826),
.A2(n_1761),
.B1(n_1718),
.B2(n_1784),
.Y(n_1836)
);

NOR2xp67_ASAP7_75t_SL g1837 ( 
.A(n_1813),
.B(n_1709),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1793),
.Y(n_1838)
);

AOI221x1_ASAP7_75t_L g1839 ( 
.A1(n_1813),
.A2(n_1761),
.B1(n_1717),
.B2(n_1787),
.C(n_1778),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1807),
.A2(n_1756),
.B1(n_1748),
.B2(n_1717),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1813),
.B(n_1748),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1791),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1797),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1818),
.B(n_1756),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1797),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1798),
.B(n_1763),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1816),
.A2(n_1738),
.B1(n_1717),
.B2(n_1763),
.Y(n_1847)
);

OAI31xp33_ASAP7_75t_L g1848 ( 
.A1(n_1816),
.A2(n_1781),
.A3(n_1777),
.B(n_1738),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1799),
.Y(n_1849)
);

O2A1O1Ixp5_ASAP7_75t_L g1850 ( 
.A1(n_1818),
.A2(n_1717),
.B(n_1738),
.C(n_1786),
.Y(n_1850)
);

NOR2x1p5_ASAP7_75t_L g1851 ( 
.A(n_1808),
.B(n_1709),
.Y(n_1851)
);

AOI21xp33_ASAP7_75t_SL g1852 ( 
.A1(n_1808),
.A2(n_1781),
.B(n_1777),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1812),
.A2(n_1738),
.B1(n_1767),
.B2(n_1770),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1846),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1835),
.A2(n_1819),
.B(n_1805),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1832),
.B(n_1824),
.Y(n_1856)
);

INVxp67_ASAP7_75t_L g1857 ( 
.A(n_1841),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1833),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1830),
.B(n_1798),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1828),
.B(n_1802),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1834),
.B(n_1792),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1832),
.B(n_1801),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1838),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1833),
.A2(n_1801),
.B1(n_1819),
.B2(n_1827),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1846),
.Y(n_1865)
);

AOI21xp33_ASAP7_75t_L g1866 ( 
.A1(n_1831),
.A2(n_1801),
.B(n_1813),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1840),
.A2(n_1802),
.B1(n_1827),
.B2(n_1824),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1853),
.A2(n_1792),
.B1(n_1767),
.B2(n_1770),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1838),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1840),
.A2(n_1853),
.B1(n_1847),
.B2(n_1836),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1851),
.B(n_1792),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1829),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1842),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1854),
.Y(n_1874)
);

XOR2x2_ASAP7_75t_L g1875 ( 
.A(n_1864),
.B(n_1844),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1865),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1871),
.B(n_1844),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1863),
.Y(n_1878)
);

OAI31xp33_ASAP7_75t_L g1879 ( 
.A1(n_1864),
.A2(n_1848),
.A3(n_1839),
.B(n_1849),
.Y(n_1879)
);

NOR3xp33_ASAP7_75t_L g1880 ( 
.A(n_1858),
.B(n_1852),
.C(n_1850),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1862),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1857),
.B(n_1843),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1859),
.B(n_1837),
.Y(n_1883)
);

OAI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1855),
.A2(n_1823),
.B(n_1822),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1881),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1877),
.B(n_1869),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1882),
.B(n_1861),
.Y(n_1887)
);

NAND4xp25_ASAP7_75t_L g1888 ( 
.A(n_1879),
.B(n_1883),
.C(n_1880),
.D(n_1860),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1874),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1876),
.Y(n_1890)
);

NOR4xp25_ASAP7_75t_L g1891 ( 
.A(n_1882),
.B(n_1873),
.C(n_1872),
.D(n_1870),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1878),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1875),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1875),
.B(n_1862),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1884),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1891),
.A2(n_1883),
.B(n_1870),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1893),
.B(n_1867),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1887),
.Y(n_1898)
);

OAI211xp5_ASAP7_75t_L g1899 ( 
.A1(n_1888),
.A2(n_1866),
.B(n_1867),
.C(n_1868),
.Y(n_1899)
);

AOI322xp5_ASAP7_75t_L g1900 ( 
.A1(n_1894),
.A2(n_1845),
.A3(n_1803),
.B1(n_1799),
.B2(n_1809),
.C1(n_1821),
.C2(n_1817),
.Y(n_1900)
);

A2O1A1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1896),
.A2(n_1887),
.B(n_1895),
.C(n_1886),
.Y(n_1901)
);

OAI311xp33_ASAP7_75t_L g1902 ( 
.A1(n_1897),
.A2(n_1885),
.A3(n_1890),
.B1(n_1889),
.C1(n_1856),
.Y(n_1902)
);

OAI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1899),
.A2(n_1892),
.B1(n_1822),
.B2(n_1823),
.C(n_1803),
.Y(n_1903)
);

AOI222xp33_ASAP7_75t_L g1904 ( 
.A1(n_1898),
.A2(n_1809),
.B1(n_1821),
.B2(n_1817),
.C1(n_1815),
.C2(n_1814),
.Y(n_1904)
);

OAI211xp5_ASAP7_75t_L g1905 ( 
.A1(n_1900),
.A2(n_1815),
.B(n_1806),
.C(n_1814),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1899),
.A2(n_1738),
.B1(n_1814),
.B2(n_1811),
.Y(n_1906)
);

XNOR2x1_ASAP7_75t_L g1907 ( 
.A(n_1902),
.B(n_1774),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1901),
.B(n_1774),
.Y(n_1908)
);

NAND4xp75_ASAP7_75t_L g1909 ( 
.A(n_1906),
.B(n_1804),
.C(n_1800),
.D(n_1811),
.Y(n_1909)
);

OAI211xp5_ASAP7_75t_L g1910 ( 
.A1(n_1903),
.A2(n_1811),
.B(n_1806),
.C(n_1804),
.Y(n_1910)
);

NAND4xp75_ASAP7_75t_L g1911 ( 
.A(n_1905),
.B(n_1806),
.C(n_1800),
.D(n_1804),
.Y(n_1911)
);

NOR3xp33_ASAP7_75t_L g1912 ( 
.A(n_1908),
.B(n_1904),
.C(n_1800),
.Y(n_1912)
);

AOI211xp5_ASAP7_75t_L g1913 ( 
.A1(n_1910),
.A2(n_1786),
.B(n_1720),
.C(n_1716),
.Y(n_1913)
);

AND3x2_ASAP7_75t_L g1914 ( 
.A(n_1907),
.B(n_1909),
.C(n_1911),
.Y(n_1914)
);

OAI22x1_ASAP7_75t_L g1915 ( 
.A1(n_1914),
.A2(n_1752),
.B1(n_1764),
.B2(n_1720),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1912),
.B1(n_1913),
.B2(n_1720),
.Y(n_1916)
);

AO21x2_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1779),
.B(n_1771),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1916),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1918),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1917),
.A2(n_1779),
.B(n_1771),
.Y(n_1920)
);

OAI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1919),
.A2(n_1920),
.B(n_1917),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1921),
.B(n_1716),
.Y(n_1922)
);

XNOR2x1_ASAP7_75t_L g1923 ( 
.A(n_1922),
.B(n_1554),
.Y(n_1923)
);

OAI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1923),
.A2(n_1825),
.B1(n_1725),
.B2(n_1743),
.Y(n_1924)
);

AOI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1924),
.A2(n_1723),
.B1(n_1725),
.B2(n_1730),
.C(n_1743),
.Y(n_1925)
);

AOI211xp5_ASAP7_75t_L g1926 ( 
.A1(n_1925),
.A2(n_1719),
.B(n_1554),
.C(n_1564),
.Y(n_1926)
);


endmodule