module real_jpeg_31458_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_620;
wire n_366;
wire n_332;
wire n_456;
wire n_578;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_278;
wire n_689;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_633;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_586;
wire n_120;
wire n_155;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_699;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_694;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_641;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_0),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_0),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_1),
.A2(n_51),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_1),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_1),
.A2(n_362),
.B1(n_437),
.B2(n_442),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_1),
.A2(n_222),
.B1(n_362),
.B2(n_586),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_1),
.A2(n_362),
.B1(n_639),
.B2(n_640),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_2),
.A2(n_383),
.B1(n_384),
.B2(n_386),
.Y(n_382)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_2),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_2),
.A2(n_386),
.B1(n_480),
.B2(n_483),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_2),
.A2(n_386),
.B1(n_586),
.B2(n_620),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_2),
.A2(n_386),
.B1(n_628),
.B2(n_629),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_4),
.A2(n_248),
.B1(n_252),
.B2(n_253),
.Y(n_247)
);

INVx2_ASAP7_75t_R g252 ( 
.A(n_4),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_4),
.A2(n_252),
.B1(n_388),
.B2(n_391),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_4),
.A2(n_252),
.B1(n_538),
.B2(n_541),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_4),
.A2(n_252),
.B1(n_603),
.B2(n_607),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_5),
.A2(n_158),
.B1(n_159),
.B2(n_161),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_5),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_5),
.A2(n_158),
.B1(n_260),
.B2(n_264),
.Y(n_259)
);

AOI21x1_ASAP7_75t_L g366 ( 
.A1(n_5),
.A2(n_367),
.B(n_371),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_5),
.A2(n_158),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_6),
.A2(n_357),
.B(n_359),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_6),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_6),
.B(n_455),
.Y(n_454)
);

OAI32xp33_ASAP7_75t_L g546 ( 
.A1(n_6),
.A2(n_187),
.A3(n_547),
.B1(n_550),
.B2(n_556),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_6),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_6),
.B(n_208),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_SL g645 ( 
.A1(n_6),
.A2(n_229),
.B1(n_638),
.B2(n_646),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_6),
.A2(n_557),
.B1(n_664),
.B2(n_669),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_7),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

INVx2_ASAP7_75t_R g170 ( 
.A(n_7),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_7),
.A2(n_170),
.B1(n_374),
.B2(n_377),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_7),
.A2(n_170),
.B1(n_179),
.B2(n_472),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_7),
.A2(n_170),
.B1(n_564),
.B2(n_568),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_9),
.Y(n_195)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_10),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_10),
.Y(n_571)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_11),
.Y(n_116)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_11),
.Y(n_125)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_11),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_12),
.A2(n_65),
.B1(n_68),
.B2(n_75),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_12),
.A2(n_75),
.B1(n_105),
.B2(n_108),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_12),
.A2(n_75),
.B1(n_218),
.B2(n_221),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_12),
.A2(n_75),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_13),
.A2(n_179),
.B1(n_181),
.B2(n_184),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_13),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_13),
.A2(n_184),
.B1(n_240),
.B2(n_244),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_13),
.A2(n_168),
.B1(n_184),
.B2(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_13),
.A2(n_184),
.B1(n_417),
.B2(n_420),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_14),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_14),
.Y(n_700)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_15),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_16),
.A2(n_49),
.B1(n_56),
.B2(n_61),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_16),
.A2(n_61),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_16),
.A2(n_61),
.B1(n_106),
.B2(n_231),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_16),
.A2(n_61),
.B1(n_287),
.B2(n_292),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_17),
.Y(n_119)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_17),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_17),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_17),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_18),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_18),
.Y(n_198)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_18),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_19),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_19),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_19),
.A2(n_136),
.B1(n_181),
.B2(n_204),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_19),
.A2(n_136),
.B1(n_309),
.B2(n_312),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_19),
.A2(n_136),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

OAI311xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_83),
.A3(n_691),
.B1(n_695),
.C1(n_698),
.Y(n_20)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_21),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_23),
.B(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_23),
.B(n_342),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_48),
.B1(n_62),
.B2(n_64),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_24),
.A2(n_78),
.B1(n_247),
.B2(n_255),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_24),
.A2(n_78),
.B1(n_274),
.B2(n_308),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g355 ( 
.A1(n_24),
.A2(n_62),
.B1(n_356),
.B2(n_361),
.Y(n_355)
);

OAI22x1_ASAP7_75t_L g502 ( 
.A1(n_24),
.A2(n_62),
.B1(n_247),
.B2(n_479),
.Y(n_502)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2x1p5_ASAP7_75t_L g166 ( 
.A(n_25),
.B(n_167),
.Y(n_166)
);

NAND2xp33_ASAP7_75t_SL g279 ( 
.A(n_25),
.B(n_157),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_25),
.A2(n_154),
.B1(n_478),
.B2(n_485),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_37),
.Y(n_25)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_28),
.Y(n_266)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_29),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g294 ( 
.A(n_29),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_29),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_29),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_32),
.Y(n_401)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_32),
.Y(n_410)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_34),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_34),
.Y(n_390)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_39),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_40),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_40),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_40),
.Y(n_482)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_45),
.Y(n_169)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_48),
.A2(n_62),
.B1(n_80),
.B2(n_308),
.Y(n_336)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_53),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_53),
.Y(n_311)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_54),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_62),
.Y(n_455)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_78),
.B(n_80),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g432 ( 
.A1(n_69),
.A2(n_397),
.A3(n_402),
.B1(n_406),
.B2(n_414),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_73),
.Y(n_358)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_83),
.B(n_696),
.Y(n_695)
);

OAI221xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_340),
.B1(n_343),
.B2(n_348),
.C(n_689),
.Y(n_83)
);

OA21x2_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_325),
.B(n_339),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_301),
.B(n_324),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_268),
.Y(n_86)
);

NOR2xp67_ASAP7_75t_SL g346 ( 
.A(n_87),
.B(n_268),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_174),
.C(n_226),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_89),
.B(n_506),
.Y(n_505)
);

XNOR2x1_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_151),
.Y(n_89)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_90),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_111),
.Y(n_90)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_91),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_91),
.B(n_111),
.Y(n_496)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B(n_103),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx8_ASAP7_75t_L g463 ( 
.A(n_94),
.Y(n_463)
);

INVx4_ASAP7_75t_SL g646 ( 
.A(n_94),
.Y(n_646)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_95),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_95),
.A2(n_416),
.B1(n_423),
.B2(n_425),
.Y(n_415)
);

AO22x1_ASAP7_75t_L g562 ( 
.A1(n_95),
.A2(n_423),
.B1(n_449),
.B2(n_563),
.Y(n_562)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_96),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_96),
.A2(n_230),
.B1(n_426),
.B2(n_461),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_96),
.A2(n_627),
.B1(n_638),
.B2(n_641),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_100),
.Y(n_237)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_101),
.Y(n_419)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_101),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_102),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_102),
.Y(n_606)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_102),
.Y(n_610)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_104),
.A2(n_229),
.B1(n_230),
.B2(n_234),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_127),
.B1(n_128),
.B2(n_131),
.Y(n_126)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_110),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_132),
.B1(n_142),
.B2(n_144),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_112),
.A2(n_132),
.B1(n_142),
.B2(n_239),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g282 ( 
.A1(n_112),
.A2(n_142),
.B(n_217),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_112),
.A2(n_142),
.B1(n_366),
.B2(n_373),
.Y(n_365)
);

OAI22x1_ASAP7_75t_SL g464 ( 
.A1(n_112),
.A2(n_142),
.B1(n_239),
.B2(n_366),
.Y(n_464)
);

OAI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_112),
.A2(n_142),
.B1(n_373),
.B2(n_536),
.Y(n_535)
);

OAI22x1_ASAP7_75t_L g617 ( 
.A1(n_112),
.A2(n_142),
.B1(n_618),
.B2(n_619),
.Y(n_617)
);

AO21x2_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_120),
.B(n_126),
.Y(n_112)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_113),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_119),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_119),
.Y(n_543)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_119),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_126),
.Y(n_214)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_127),
.Y(n_430)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_130),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_134),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_199)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_140),
.Y(n_372)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_140),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_141),
.Y(n_376)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_142),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_142),
.B(n_557),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_144),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_147),
.Y(n_244)
);

BUFx6f_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_173),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_152),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_156),
.B(n_166),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g273 ( 
.A1(n_153),
.A2(n_274),
.B(n_279),
.Y(n_273)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_158),
.B(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_161),
.Y(n_312)
);

OAI32xp33_ASAP7_75t_L g396 ( 
.A1(n_161),
.A2(n_397),
.A3(n_402),
.B1(n_406),
.B2(n_414),
.Y(n_396)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_165),
.Y(n_251)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_165),
.Y(n_484)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_167),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_175),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_225),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_210),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_210),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_185),
.B1(n_203),
.B2(n_208),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_178),
.A2(n_208),
.B1(n_258),
.B2(n_267),
.Y(n_257)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_181),
.Y(n_318)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_182),
.Y(n_442)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_183),
.Y(n_413)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_185),
.Y(n_334)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_186),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_186),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_186),
.A2(n_285),
.B1(n_286),
.B2(n_316),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_186),
.A2(n_285),
.B1(n_387),
.B2(n_471),
.Y(n_470)
);

OAI22x1_ASAP7_75t_L g500 ( 
.A1(n_186),
.A2(n_259),
.B1(n_285),
.B2(n_471),
.Y(n_500)
);

AO21x2_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_192),
.B(n_199),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_188),
.Y(n_383)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_197),
.Y(n_322)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_198),
.Y(n_385)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_201),
.Y(n_370)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_201),
.Y(n_561)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_203),
.Y(n_284)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_206),
.Y(n_405)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_206),
.Y(n_476)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_206),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_207),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_207),
.Y(n_394)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_208),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_208),
.A2(n_333),
.B(n_335),
.Y(n_332)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g662 ( 
.A1(n_209),
.A2(n_381),
.B1(n_436),
.B2(n_663),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_215),
.B1(n_216),
.B2(n_224),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_211),
.A2(n_579),
.B1(n_584),
.B2(n_585),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_211),
.A2(n_224),
.B1(n_537),
.B2(n_673),
.Y(n_672)
);

OA21x2_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B(n_214),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g588 ( 
.A1(n_213),
.A2(n_589),
.B(n_592),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_214),
.Y(n_584)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_225),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_225),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_226),
.B(n_505),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_245),
.C(n_256),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_227),
.B(n_493),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_238),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_228),
.B(n_238),
.Y(n_517)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_232),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_232),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx6_ASAP7_75t_L g591 ( 
.A(n_233),
.Y(n_591)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_233),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_233),
.Y(n_653)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx4f_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_243),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_L g493 ( 
.A1(n_246),
.A2(n_256),
.B1(n_257),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_246),
.Y(n_494)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_254),
.Y(n_360)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_267),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_298),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_280),
.B1(n_281),
.B2(n_297),
.Y(n_269)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_298),
.C(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_272),
.A2(n_273),
.B1(n_280),
.B2(n_281),
.Y(n_303)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_273),
.B(n_283),
.C(n_295),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_273),
.B(n_323),
.C(n_338),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx11_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_295),
.B2(n_296),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_282),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_295),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_282),
.B(n_307),
.C(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_285),
.A2(n_381),
.B1(n_382),
.B2(n_387),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_285),
.A2(n_334),
.B1(n_382),
.B2(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_301),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_302),
.B(n_304),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_323),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_313),
.Y(n_306)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

NOR2x1_ASAP7_75t_R g325 ( 
.A(n_326),
.B(n_337),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_337),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_330),
.B2(n_331),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_332),
.C(n_336),
.Y(n_342)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_336),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND3xp33_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_344),
.C(n_345),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_527),
.B(n_684),
.Y(n_349)
);

NAND4xp25_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_489),
.C(n_507),
.D(n_520),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_456),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_352),
.B(n_456),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_395),
.C(n_434),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_353),
.B(n_530),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_364),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_355),
.B(n_365),
.C(n_380),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_358),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_359),
.Y(n_414)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_361),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_380),
.Y(n_364)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_394),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_395),
.B(n_434),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_415),
.B1(n_431),
.B2(n_433),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_396),
.B(n_433),
.Y(n_488)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_411),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_415),
.Y(n_433)
);

AO22x1_ASAP7_75t_SL g443 ( 
.A1(n_416),
.A2(n_444),
.B1(n_448),
.B2(n_449),
.Y(n_443)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_443),
.C(n_453),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_435),
.B(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_443),
.B(n_454),
.Y(n_533)
);

INVx3_ASAP7_75t_SL g444 ( 
.A(n_445),
.Y(n_444)
);

INVx8_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_447),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_447),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_447),
.Y(n_650)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_448),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_448),
.A2(n_462),
.B1(n_626),
.B2(n_633),
.Y(n_625)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_467),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_465),
.B2(n_466),
.Y(n_457)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_458),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g522 ( 
.A(n_458),
.Y(n_522)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_459),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_464),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_460),
.B(n_464),
.Y(n_503)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_466),
.B(n_468),
.C(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_488),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_477),
.B1(n_486),
.B2(n_487),
.Y(n_469)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_477),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_477),
.Y(n_515)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_486),
.Y(n_516)
);

INVxp33_ASAP7_75t_L g514 ( 
.A(n_488),
.Y(n_514)
);

A2O1A1O1Ixp25_ASAP7_75t_L g684 ( 
.A1(n_489),
.A2(n_507),
.B(n_685),
.C(n_687),
.D(n_688),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_504),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_490),
.B(n_504),
.Y(n_688)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_495),
.C(n_497),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_519),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_498),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

MAJx2_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_501),
.C(n_503),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_499),
.A2(n_500),
.B1(n_502),
.B2(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_502),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_518),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_508),
.B(n_518),
.Y(n_687)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_513),
.C(n_517),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_526),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.C(n_516),
.Y(n_513)
);

MAJx2_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_515),
.C(n_516),
.Y(n_524)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_517),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_523),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g685 ( 
.A(n_521),
.B(n_523),
.C(n_686),
.Y(n_685)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_525),
.Y(n_523)
);

AOI21x1_ASAP7_75t_L g527 ( 
.A1(n_528),
.A2(n_572),
.B(n_683),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_529),
.B(n_531),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_SL g683 ( 
.A(n_529),
.B(n_531),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_534),
.C(n_544),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g678 ( 
.A(n_532),
.B(n_679),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_534),
.A2(n_545),
.B(n_680),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g680 ( 
.A(n_535),
.B(n_545),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_543),
.Y(n_581)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_562),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_SL g660 ( 
.A(n_546),
.B(n_562),
.Y(n_660)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_553),
.Y(n_583)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_554),
.Y(n_586)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_558),
.Y(n_556)
);

OAI21xp33_ASAP7_75t_SL g579 ( 
.A1(n_557),
.A2(n_580),
.B(n_582),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_557),
.B(n_583),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_557),
.B(n_649),
.Y(n_648)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_563),
.Y(n_614)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_571),
.Y(n_595)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_571),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_573),
.A2(n_677),
.B(n_682),
.Y(n_572)
);

AOI21x1_ASAP7_75t_L g573 ( 
.A1(n_574),
.A2(n_657),
.B(n_676),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_575),
.A2(n_623),
.B(n_656),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_599),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_576),
.B(n_599),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_577),
.B(n_587),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_577),
.A2(n_578),
.B1(n_587),
.B2(n_588),
.Y(n_634)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_582),
.A2(n_593),
.B(n_596),
.Y(n_592)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_585),
.Y(n_618)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_594),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_600),
.B(n_615),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_600),
.B(n_617),
.C(n_621),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_601),
.A2(n_602),
.B1(n_611),
.B2(n_614),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_602),
.Y(n_633)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_605),
.Y(n_628)
);

INVx6_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_616),
.A2(n_617),
.B1(n_621),
.B2(n_622),
.Y(n_615)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_616),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_617),
.Y(n_622)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_619),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_624),
.A2(n_635),
.B(n_655),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_625),
.B(n_634),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_625),
.B(n_634),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_628),
.Y(n_640)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_636),
.A2(n_644),
.B(n_654),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_637),
.B(n_643),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_637),
.B(n_643),
.Y(n_654)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_642),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_645),
.B(n_647),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_R g647 ( 
.A(n_648),
.B(n_651),
.Y(n_647)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_652),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_658),
.B(n_659),
.Y(n_657)
);

NOR2x1_ASAP7_75t_SL g676 ( 
.A(n_658),
.B(n_659),
.Y(n_676)
);

XNOR2xp5_ASAP7_75t_L g659 ( 
.A(n_660),
.B(n_661),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g681 ( 
.A(n_660),
.B(n_672),
.C(n_675),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_662),
.A2(n_672),
.B1(n_674),
.B2(n_675),
.Y(n_661)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_662),
.Y(n_675)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_665),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_666),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_667),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_668),
.Y(n_667)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_670),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_671),
.Y(n_670)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_672),
.Y(n_674)
);

NOR2x1_ASAP7_75t_SL g677 ( 
.A(n_678),
.B(n_681),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_678),
.B(n_681),
.Y(n_682)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_690),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_691),
.B(n_697),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_691),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_692),
.B(n_694),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_693),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_699),
.B(n_700),
.Y(n_698)
);


endmodule