module real_jpeg_12398_n_12 (n_5, n_4, n_8, n_0, n_299, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_299;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_288;
wire n_78;
wire n_286;
wire n_176;
wire n_221;
wire n_215;
wire n_292;
wire n_249;
wire n_166;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_200;
wire n_184;
wire n_275;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_3),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_3),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_22),
.B1(n_27),
.B2(n_40),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_3),
.A2(n_40),
.B1(n_51),
.B2(n_56),
.Y(n_288)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_6),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_28),
.B1(n_51),
.B2(n_56),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_6),
.A2(n_28),
.B1(n_33),
.B2(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_6),
.A2(n_28),
.B1(n_58),
.B2(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_70),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_6),
.B(n_22),
.C(n_36),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_6),
.B(n_86),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_6),
.B(n_38),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_6),
.A2(n_59),
.B(n_72),
.C(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_6),
.B(n_57),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_9),
.A2(n_51),
.B1(n_56),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_9),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_9),
.A2(n_22),
.B1(n_27),
.B2(n_101),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_9),
.A2(n_33),
.B1(n_37),
.B2(n_101),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_101),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_10),
.A2(n_33),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_10),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_10),
.A2(n_22),
.B1(n_27),
.B2(n_43),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_10),
.A2(n_43),
.B1(n_51),
.B2(n_56),
.Y(n_110)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_277),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_122),
.B(n_275),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_102),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_16),
.B(n_102),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_62),
.C(n_79),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_17),
.A2(n_18),
.B1(n_62),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_19),
.A2(n_20),
.B(n_46),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_20),
.A2(n_45),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_20),
.B(n_180),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_20),
.A2(n_29),
.B1(n_45),
.B2(n_266),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_26),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_21),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_21),
.B(n_26),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_21),
.A2(n_211),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g38 ( 
.A1(n_22),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_22),
.B(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_25),
.B(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_25),
.B(n_83),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_25),
.A2(n_82),
.B(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_28),
.A2(n_37),
.B(n_73),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_28),
.B(n_54),
.C(n_59),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_29),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_39),
.B(n_41),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_30),
.A2(n_67),
.B(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_31),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_31),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_31),
.B(n_66),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_33),
.A2(n_37),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_33),
.B(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_38),
.B(n_139),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_39),
.A2(n_64),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_41),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_41),
.B(n_150),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_60),
.B(n_61),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_48),
.B(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_49),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_49),
.B(n_110),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_57),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_50)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_54),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_56),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_57),
.B(n_100),
.Y(n_217)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_59),
.B1(n_72),
.B2(n_73),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_60),
.A2(n_239),
.B(n_288),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_62),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_68),
.B(n_78),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_68),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_64),
.B(n_149),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_65),
.B(n_138),
.Y(n_187)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_74),
.Y(n_68)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_70),
.B(n_177),
.Y(n_176)
);

NAND2x1_ASAP7_75t_SL g228 ( 
.A(n_70),
.B(n_94),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_70),
.A2(n_93),
.B(n_94),
.Y(n_240)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_77),
.Y(n_90)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_74),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_74),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_75),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_105),
.B1(n_106),
.B2(n_121),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_78),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_78),
.B(n_103),
.C(n_105),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_79),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_89),
.C(n_95),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_80),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_81),
.B(n_87),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_82),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_89),
.A2(n_95),
.B1(n_96),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_89),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_90),
.B(n_193),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_92),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_99),
.B(n_109),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_114),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_107),
.B(n_116),
.C(n_117),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_107),
.A2(n_108),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_112),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_115),
.A2(n_116),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_115),
.B(n_215),
.C(n_220),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_115),
.A2(n_116),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_269),
.B(n_274),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_256),
.B(n_268),
.Y(n_123)
);

AOI321xp33_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_223),
.A3(n_249),
.B1(n_254),
.B2(n_255),
.C(n_299),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_200),
.B(n_222),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_184),
.B(n_199),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_171),
.B(n_183),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_151),
.B(n_170),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_144),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_144),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_135),
.B1(n_136),
.B2(n_143),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_131),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_141),
.C(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_164),
.B(n_169),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_159),
.B(n_163),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_162),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_198),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_198),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_189),
.C(n_191),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_196),
.C(n_197),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_213),
.B2(n_214),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_206),
.C(n_213),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_212),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_244),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_244),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_232),
.C(n_243),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.C(n_230),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_226),
.B(n_227),
.CI(n_230),
.CON(n_246),
.SN(n_246)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_228),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_243),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_240),
.C(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_236),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.C(n_248),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_246),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_246),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_248),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_253),
.Y(n_254)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_258),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_267),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_265),
.C(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_295),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_280),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_289),
.B1(n_290),
.B2(n_294),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_287),
.Y(n_294)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);


endmodule