module fake_jpeg_25702_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_14),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_70),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_59),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_62),
.C(n_58),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_79),
.Y(n_90)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_78),
.Y(n_101)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_96),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_63),
.B1(n_54),
.B2(n_48),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_95),
.B1(n_64),
.B2(n_60),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_50),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_52),
.B1(n_45),
.B2(n_47),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_100),
.B1(n_102),
.B2(n_49),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_63),
.B1(n_56),
.B2(n_49),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_0),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_43),
.B1(n_51),
.B2(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_55),
.B1(n_56),
.B2(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_105),
.Y(n_117)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_102),
.B1(n_95),
.B2(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_94),
.B1(n_53),
.B2(n_2),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_0),
.Y(n_130)
);

AOI32xp33_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_98),
.A3(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_35),
.B(n_32),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_131),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_115),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_110),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_136),
.B(n_137),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_91),
.B1(n_110),
.B2(n_87),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_8),
.B1(n_40),
.B2(n_39),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_1),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_134),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_37),
.B(n_36),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_119),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_2),
.C(n_3),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_28),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_141),
.B(n_146),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_3),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_4),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_128),
.B1(n_125),
.B2(n_127),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_147),
.C(n_143),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_144),
.A2(n_25),
.B1(n_12),
.B2(n_9),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_139),
.B(n_7),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_152),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_142),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_149),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_148),
.B(n_138),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_156),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_145),
.Y(n_158)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_158),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_145),
.B(n_6),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_4),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);


endmodule