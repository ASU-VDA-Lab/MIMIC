module fake_jpeg_19754_n_108 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_1),
.B(n_4),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_37),
.B1(n_38),
.B2(n_36),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_43),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_26),
.B(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_20),
.B1(n_14),
.B2(n_19),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_15),
.B1(n_22),
.B2(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_18),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_48),
.C(n_43),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_6),
.C(n_7),
.Y(n_74)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_56),
.Y(n_71)
);

AOI32xp33_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_35),
.A3(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_31),
.B(n_34),
.C(n_23),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_67),
.B(n_34),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_22),
.B(n_21),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_68),
.B(n_9),
.Y(n_79)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_64),
.B1(n_52),
.B2(n_58),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_1),
.B1(n_12),
.B2(n_7),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_66),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_34),
.B1(n_19),
.B2(n_14),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_16),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_58),
.B1(n_66),
.B2(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_64),
.B1(n_58),
.B2(n_10),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_80),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_54),
.B(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_73),
.Y(n_92)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_87),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_72),
.B1(n_76),
.B2(n_71),
.Y(n_89)
);

XNOR2x1_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_80),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_82),
.B(n_79),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_90),
.A2(n_88),
.B(n_83),
.C(n_78),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_95),
.B(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_98),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_92),
.C(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_98),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_100),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_106),
.Y(n_108)
);


endmodule