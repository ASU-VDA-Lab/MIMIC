module fake_netlist_6_4960_n_672 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_77, n_92, n_42, n_8, n_90, n_24, n_54, n_0, n_87, n_32, n_66, n_85, n_78, n_84, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_80, n_41, n_86, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_672);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_77;
input n_92;
input n_42;
input n_8;
input n_90;
input n_24;
input n_54;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_78;
input n_84;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_80;
input n_41;
input n_86;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_672;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_255;
wire n_400;
wire n_284;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_108;
wire n_639;
wire n_327;
wire n_369;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_300;
wire n_248;
wire n_517;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_621;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_111;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_603;
wire n_119;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_101;
wire n_167;
wire n_631;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_656;
wire n_96;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_647;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_109;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_122;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_112;
wire n_172;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_107;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_570;
wire n_406;
wire n_483;
wire n_102;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_630;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_164;
wire n_100;
wire n_307;
wire n_121;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_124;
wire n_548;
wire n_94;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_523;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_319;
wire n_139;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_123;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_113;
wire n_618;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_99;
wire n_257;
wire n_655;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_120;
wire n_301;
wire n_274;
wire n_636;
wire n_151;
wire n_110;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVxp33_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_17),
.Y(n_102)
);

INVxp33_ASAP7_75t_SL g103 ( 
.A(n_34),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

INVxp67_ASAP7_75t_SL g111 ( 
.A(n_33),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_19),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_20),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_9),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

NOR2xp67_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_64),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_46),
.B(n_85),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_29),
.Y(n_123)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_59),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_27),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_40),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_54),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_0),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_38),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_9),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_22),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_35),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_31),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_32),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_63),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_16),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_39),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_82),
.Y(n_149)
);

INVxp33_ASAP7_75t_SL g150 ( 
.A(n_8),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_81),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_12),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_8),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_42),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_17),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_76),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_26),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_14),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_13),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_47),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_41),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_28),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_48),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_12),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_65),
.B(n_74),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_3),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_0),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_15),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_23),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_36),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_73),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_10),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_53),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_6),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_10),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_11),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_1),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_150),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_109),
.B(n_2),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_160),
.B(n_4),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_93),
.B(n_5),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_93),
.B(n_7),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_137),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_104),
.B(n_174),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_133),
.A2(n_11),
.B1(n_14),
.B2(n_16),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_141),
.B(n_18),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_106),
.B(n_24),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_133),
.B(n_37),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_134),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_156),
.B(n_49),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_134),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_101),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_136),
.B(n_57),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_114),
.B(n_67),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_114),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_102),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_117),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_106),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_154),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_97),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_118),
.B(n_75),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_118),
.B(n_80),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_157),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_122),
.B(n_91),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_150),
.A2(n_167),
.B1(n_175),
.B2(n_169),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_171),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_125),
.B(n_129),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_125),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_141),
.B(n_103),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_100),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_136),
.B(n_151),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_105),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_107),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_153),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_151),
.B(n_132),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_108),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_115),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_116),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_119),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_126),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_110),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_94),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_123),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_110),
.A2(n_143),
.B1(n_103),
.B2(n_178),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_143),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_138),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_112),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_251),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_203),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g263 ( 
.A(n_211),
.B(n_217),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_212),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_181),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_251),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_256),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_95),
.Y(n_271)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_98),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_253),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_212),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_230),
.Y(n_280)
);

AO22x2_ASAP7_75t_L g281 ( 
.A1(n_205),
.A2(n_210),
.B1(n_182),
.B2(n_191),
.Y(n_281)
);

AND2x6_ASAP7_75t_L g282 ( 
.A(n_217),
.B(n_168),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_230),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_203),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_187),
.B(n_94),
.Y(n_285)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_210),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_96),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_230),
.Y(n_289)
);

AO22x2_ASAP7_75t_L g290 ( 
.A1(n_210),
.A2(n_148),
.B1(n_161),
.B2(n_155),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_256),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_210),
.B(n_207),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_190),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

OR2x6_ASAP7_75t_L g295 ( 
.A(n_189),
.B(n_120),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_203),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_203),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_244),
.B(n_147),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_212),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_182),
.B(n_178),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_190),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_184),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_201),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_199),
.B(n_96),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_225),
.B(n_173),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_191),
.B(n_192),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_234),
.B(n_158),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_235),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_235),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_213),
.B(n_158),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_225),
.B(n_145),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_208),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_184),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_235),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_199),
.B(n_99),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_220),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_255),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_293),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_276),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_258),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_216),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_293),
.B(n_216),
.Y(n_325)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_282),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_275),
.B(n_247),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_263),
.B(n_243),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

NAND2x1p5_ASAP7_75t_L g330 ( 
.A(n_264),
.B(n_152),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_275),
.B(n_311),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_257),
.Y(n_333)
);

O2A1O1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_301),
.A2(n_257),
.B(n_250),
.C(n_249),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_260),
.Y(n_336)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_280),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_263),
.B(n_287),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_264),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_215),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_271),
.B(n_247),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_279),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_304),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_261),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_260),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_283),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_260),
.Y(n_352)
);

NAND3xp33_ASAP7_75t_L g353 ( 
.A(n_285),
.B(n_240),
.C(n_249),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_305),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_268),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_269),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_221),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_260),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_262),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_292),
.B(n_285),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_267),
.B(n_242),
.Y(n_361)
);

OR2x6_ASAP7_75t_L g362 ( 
.A(n_291),
.B(n_186),
.Y(n_362)
);

BUFx12f_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_262),
.Y(n_364)
);

OR2x6_ASAP7_75t_L g365 ( 
.A(n_295),
.B(n_186),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_267),
.Y(n_366)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_282),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_270),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_270),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_318),
.A2(n_231),
.B1(n_159),
.B2(n_149),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_314),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_287),
.B(n_243),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_308),
.B(n_259),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_288),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_289),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_329),
.Y(n_376)
);

AOI21xp33_ASAP7_75t_L g377 ( 
.A1(n_332),
.A2(n_333),
.B(n_360),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

AOI221xp5_ASAP7_75t_L g379 ( 
.A1(n_332),
.A2(n_327),
.B1(n_281),
.B2(n_231),
.C(n_370),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_329),
.Y(n_380)
);

OR2x6_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_281),
.Y(n_381)
);

AND2x4_ASAP7_75t_SL g382 ( 
.A(n_366),
.B(n_316),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_319),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_354),
.A2(n_286),
.B(n_272),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_348),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_344),
.B(n_300),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_282),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_319),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_327),
.B(n_295),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_324),
.B(n_300),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_335),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_320),
.B(n_317),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_360),
.A2(n_282),
.B1(n_295),
.B2(n_259),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_333),
.A2(n_281),
.B1(n_290),
.B2(n_308),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_355),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_366),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_372),
.A2(n_290),
.B1(n_286),
.B2(n_303),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_335),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_341),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_356),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_343),
.Y(n_406)
);

O2A1O1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_373),
.A2(n_331),
.B(n_334),
.C(n_340),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_347),
.A2(n_290),
.B1(n_286),
.B2(n_272),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_361),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_351),
.Y(n_411)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_336),
.Y(n_412)
);

BUFx6f_ASAP7_75t_SL g413 ( 
.A(n_365),
.Y(n_413)
);

NOR2x1_ASAP7_75t_SL g414 ( 
.A(n_326),
.B(n_218),
.Y(n_414)
);

BUFx2_ASAP7_75t_R g415 ( 
.A(n_342),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_325),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_331),
.B(n_322),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_370),
.A2(n_298),
.B1(n_198),
.B2(n_196),
.Y(n_419)
);

A2O1A1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_325),
.A2(n_229),
.B(n_226),
.C(n_227),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_326),
.B(n_312),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_322),
.B(n_221),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_326),
.A2(n_309),
.B(n_277),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_369),
.B(n_215),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_357),
.A2(n_243),
.B1(n_235),
.B2(n_163),
.Y(n_427)
);

BUFx6f_ASAP7_75t_SL g428 ( 
.A(n_365),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_342),
.B(n_223),
.Y(n_429)
);

OAI21xp33_ASAP7_75t_SL g430 ( 
.A1(n_369),
.A2(n_240),
.B(n_242),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_326),
.B(n_159),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_R g432 ( 
.A(n_358),
.B(n_127),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_321),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_323),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_337),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_365),
.A2(n_202),
.B1(n_196),
.B2(n_198),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_330),
.Y(n_438)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_336),
.Y(n_439)
);

OR2x6_ASAP7_75t_L g440 ( 
.A(n_362),
.B(n_223),
.Y(n_440)
);

OAI221xp5_ASAP7_75t_L g441 ( 
.A1(n_353),
.A2(n_250),
.B1(n_246),
.B2(n_204),
.C(n_202),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_337),
.B(n_149),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_362),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_330),
.Y(n_444)
);

NAND2x1p5_ASAP7_75t_L g445 ( 
.A(n_337),
.B(n_277),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_345),
.A2(n_111),
.B1(n_124),
.B2(n_121),
.Y(n_446)
);

AOI222xp33_ASAP7_75t_L g447 ( 
.A1(n_362),
.A2(n_209),
.B1(n_206),
.B2(n_200),
.C1(n_197),
.C2(n_233),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_346),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_337),
.B(n_315),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_350),
.Y(n_450)
);

NAND2x1_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_425),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_379),
.A2(n_367),
.B1(n_204),
.B2(n_246),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

AO31x2_ASAP7_75t_L g454 ( 
.A1(n_388),
.A2(n_165),
.A3(n_139),
.B(n_140),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_401),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g456 ( 
.A1(n_392),
.A2(n_367),
.B1(n_127),
.B2(n_164),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_392),
.A2(n_367),
.B1(n_144),
.B2(n_166),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_377),
.B(n_367),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_233),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_387),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_450),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_377),
.A2(n_375),
.B1(n_374),
.B2(n_339),
.Y(n_462)
);

NAND2x1p5_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_309),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_388),
.A2(n_371),
.B(n_294),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_401),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_380),
.Y(n_466)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_449),
.A2(n_371),
.B(n_310),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_400),
.B(n_209),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_409),
.B(n_206),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_379),
.A2(n_236),
.B1(n_238),
.B2(n_237),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_426),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_378),
.A2(n_243),
.B1(n_248),
.B2(n_254),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_425),
.Y(n_474)
);

AOI221xp5_ASAP7_75t_L g475 ( 
.A1(n_419),
.A2(n_200),
.B1(n_197),
.B2(n_237),
.C(n_238),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_406),
.B(n_224),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_386),
.B(n_396),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_405),
.Y(n_478)
);

CKINVDCx8_ASAP7_75t_R g479 ( 
.A(n_399),
.Y(n_479)
);

O2A1O1Ixp33_ASAP7_75t_SL g480 ( 
.A1(n_420),
.A2(n_236),
.B(n_219),
.C(n_184),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_422),
.B(n_224),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_SL g485 ( 
.A1(n_394),
.A2(n_235),
.B1(n_248),
.B2(n_254),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_411),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_394),
.A2(n_248),
.B1(n_254),
.B2(n_232),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_449),
.A2(n_265),
.B(n_266),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_415),
.B(n_228),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_SL g490 ( 
.A1(n_418),
.A2(n_248),
.B1(n_254),
.B2(n_232),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_398),
.A2(n_254),
.B1(n_248),
.B2(n_278),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_407),
.B(n_397),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_382),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_419),
.A2(n_402),
.B1(n_381),
.B2(n_416),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_381),
.A2(n_266),
.B1(n_299),
.B2(n_278),
.Y(n_495)
);

AOI21xp33_ASAP7_75t_L g496 ( 
.A1(n_430),
.A2(n_219),
.B(n_299),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_SL g497 ( 
.A1(n_413),
.A2(n_228),
.B1(n_185),
.B2(n_194),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_383),
.Y(n_498)
);

AOI222xp33_ASAP7_75t_L g499 ( 
.A1(n_437),
.A2(n_194),
.B1(n_185),
.B2(n_195),
.C1(n_193),
.C2(n_183),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_436),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_415),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_429),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_389),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_429),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_381),
.A2(n_265),
.B1(n_219),
.B2(n_214),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_410),
.A2(n_364),
.B1(n_359),
.B2(n_352),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_408),
.A2(n_183),
.B1(n_188),
.B2(n_193),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_390),
.B(n_195),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_433),
.A2(n_214),
.B1(n_359),
.B2(n_364),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_434),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_395),
.B(n_188),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_403),
.B(n_214),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_437),
.A2(n_364),
.B1(n_359),
.B2(n_352),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_448),
.B(n_364),
.Y(n_515)
);

OAI222xp33_ASAP7_75t_L g516 ( 
.A1(n_440),
.A2(n_208),
.B1(n_359),
.B2(n_336),
.C1(n_352),
.C2(n_349),
.Y(n_516)
);

AOI221xp5_ASAP7_75t_L g517 ( 
.A1(n_441),
.A2(n_208),
.B1(n_352),
.B2(n_349),
.C(n_296),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_423),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_443),
.A2(n_208),
.B1(n_349),
.B2(n_284),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_427),
.A2(n_349),
.B1(n_208),
.B2(n_284),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_440),
.B(n_313),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_432),
.Y(n_522)
);

AOI221xp5_ASAP7_75t_L g523 ( 
.A1(n_441),
.A2(n_262),
.B1(n_284),
.B2(n_296),
.C(n_297),
.Y(n_523)
);

AOI221xp5_ASAP7_75t_L g524 ( 
.A1(n_494),
.A2(n_428),
.B1(n_413),
.B2(n_404),
.C(n_447),
.Y(n_524)
);

AOI221xp5_ASAP7_75t_L g525 ( 
.A1(n_459),
.A2(n_428),
.B1(n_447),
.B2(n_446),
.C(n_444),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_477),
.A2(n_440),
.B1(n_442),
.B2(n_431),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_492),
.A2(n_421),
.B1(n_384),
.B2(n_445),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_453),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_466),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_L g530 ( 
.A1(n_489),
.A2(n_421),
.B1(n_439),
.B2(n_423),
.Y(n_530)
);

AOI211xp5_ASAP7_75t_L g531 ( 
.A1(n_460),
.A2(n_424),
.B(n_284),
.C(n_296),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_492),
.A2(n_445),
.B1(n_412),
.B2(n_423),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_456),
.A2(n_412),
.B1(n_439),
.B2(n_297),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_472),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_484),
.B(n_414),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_L g536 ( 
.A1(n_489),
.A2(n_439),
.B1(n_412),
.B2(n_297),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_461),
.A2(n_412),
.B1(n_296),
.B2(n_297),
.Y(n_537)
);

AOI21xp33_ASAP7_75t_SL g538 ( 
.A1(n_468),
.A2(n_262),
.B(n_313),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_452),
.A2(n_313),
.B1(n_511),
.B2(n_503),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_471),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_467),
.A2(n_313),
.B(n_488),
.Y(n_541)
);

OAI22xp33_ASAP7_75t_L g542 ( 
.A1(n_522),
.A2(n_478),
.B1(n_498),
.B2(n_504),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_452),
.A2(n_504),
.B1(n_509),
.B2(n_476),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_515),
.B(n_512),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_509),
.A2(n_476),
.B1(n_457),
.B2(n_500),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_499),
.B(n_469),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_482),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_458),
.A2(n_514),
.B1(n_474),
.B2(n_506),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_455),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_486),
.A2(n_502),
.B1(n_505),
.B2(n_475),
.Y(n_551)
);

AOI221xp5_ASAP7_75t_L g552 ( 
.A1(n_475),
.A2(n_470),
.B1(n_507),
.B2(n_522),
.C(n_497),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_502),
.A2(n_458),
.B1(n_495),
.B2(n_491),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_513),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_SL g555 ( 
.A1(n_502),
.A2(n_508),
.B1(n_501),
.B2(n_455),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_455),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_481),
.B(n_465),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_470),
.A2(n_507),
.B1(n_462),
.B2(n_487),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_479),
.Y(n_559)
);

AOI221xp5_ASAP7_75t_L g560 ( 
.A1(n_501),
.A2(n_508),
.B1(n_496),
.B2(n_483),
.C(n_517),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_L g561 ( 
.A1(n_508),
.A2(n_465),
.B1(n_521),
.B2(n_481),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_485),
.A2(n_465),
.B1(n_490),
.B2(n_499),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_496),
.A2(n_473),
.B1(n_517),
.B2(n_523),
.Y(n_563)
);

A2O1A1Ixp33_ASAP7_75t_L g564 ( 
.A1(n_464),
.A2(n_519),
.B(n_523),
.C(n_451),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_464),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_454),
.B(n_510),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_493),
.Y(n_567)
);

OA21x2_ASAP7_75t_L g568 ( 
.A1(n_516),
.A2(n_520),
.B(n_454),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_534),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_547),
.B(n_454),
.Y(n_570)
);

AO21x2_ASAP7_75t_L g571 ( 
.A1(n_565),
.A2(n_480),
.B(n_463),
.Y(n_571)
);

AOI31xp33_ASAP7_75t_L g572 ( 
.A1(n_524),
.A2(n_463),
.A3(n_518),
.B(n_525),
.Y(n_572)
);

NOR3xp33_ASAP7_75t_L g573 ( 
.A(n_542),
.B(n_518),
.C(n_545),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_541),
.A2(n_565),
.B(n_564),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_547),
.B(n_545),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_544),
.B(n_540),
.Y(n_576)
);

NAND3xp33_ASAP7_75t_L g577 ( 
.A(n_552),
.B(n_560),
.C(n_558),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_558),
.B(n_546),
.C(n_526),
.Y(n_578)
);

NOR2x1_ASAP7_75t_R g579 ( 
.A(n_559),
.B(n_567),
.Y(n_579)
);

AOI221xp5_ASAP7_75t_L g580 ( 
.A1(n_563),
.A2(n_554),
.B1(n_562),
.B2(n_549),
.C(n_530),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_528),
.Y(n_581)
);

AOI33xp33_ASAP7_75t_L g582 ( 
.A1(n_555),
.A2(n_554),
.A3(n_539),
.B1(n_529),
.B2(n_548),
.B3(n_528),
.Y(n_582)
);

OAI211xp5_ASAP7_75t_SL g583 ( 
.A1(n_553),
.A2(n_551),
.B(n_529),
.C(n_548),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_543),
.Y(n_584)
);

OAI211xp5_ASAP7_75t_L g585 ( 
.A1(n_535),
.A2(n_559),
.B(n_556),
.C(n_557),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_527),
.A2(n_532),
.B(n_536),
.Y(n_586)
);

AOI222xp33_ASAP7_75t_L g587 ( 
.A1(n_567),
.A2(n_535),
.B1(n_561),
.B2(n_566),
.C1(n_543),
.C2(n_550),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_543),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_566),
.B(n_550),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_568),
.Y(n_590)
);

AO21x2_ASAP7_75t_L g591 ( 
.A1(n_541),
.A2(n_538),
.B(n_568),
.Y(n_591)
);

OAI211xp5_ASAP7_75t_L g592 ( 
.A1(n_538),
.A2(n_533),
.B(n_531),
.C(n_537),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_568),
.B(n_545),
.Y(n_593)
);

AOI33xp33_ASAP7_75t_L g594 ( 
.A1(n_547),
.A2(n_370),
.A3(n_318),
.B1(n_379),
.B2(n_494),
.B3(n_417),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_547),
.B(n_477),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_534),
.Y(n_596)
);

NAND4xp25_ASAP7_75t_SL g597 ( 
.A(n_552),
.B(n_379),
.C(n_447),
.D(n_318),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_534),
.Y(n_598)
);

NOR4xp25_ASAP7_75t_L g599 ( 
.A(n_552),
.B(n_377),
.C(n_332),
.D(n_379),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_589),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_589),
.B(n_576),
.Y(n_601)
);

OAI211xp5_ASAP7_75t_L g602 ( 
.A1(n_599),
.A2(n_577),
.B(n_578),
.C(n_580),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_577),
.B(n_575),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_590),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_581),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_578),
.B(n_594),
.C(n_573),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_596),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_575),
.B(n_595),
.Y(n_608)
);

AOI221xp5_ASAP7_75t_L g609 ( 
.A1(n_597),
.A2(n_595),
.B1(n_572),
.B2(n_570),
.C(n_586),
.Y(n_609)
);

INVxp33_ASAP7_75t_SL g610 ( 
.A(n_579),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_570),
.B(n_576),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_583),
.A2(n_587),
.B1(n_585),
.B2(n_569),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_582),
.B(n_598),
.C(n_592),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_574),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_584),
.B(n_588),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_574),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_584),
.B(n_593),
.Y(n_617)
);

AOI33xp33_ASAP7_75t_L g618 ( 
.A1(n_596),
.A2(n_370),
.A3(n_318),
.B1(n_379),
.B2(n_599),
.B3(n_494),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_593),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_579),
.B(n_593),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_614),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_617),
.B(n_593),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_611),
.B(n_591),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_608),
.B(n_571),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_614),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_607),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_611),
.B(n_601),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_601),
.B(n_600),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_605),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_608),
.B(n_571),
.Y(n_630)
);

NOR3xp33_ASAP7_75t_SL g631 ( 
.A(n_606),
.B(n_591),
.C(n_613),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_601),
.B(n_600),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_619),
.B(n_604),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_629),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_633),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_633),
.B(n_619),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_621),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_623),
.B(n_617),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_623),
.B(n_601),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_627),
.B(n_632),
.Y(n_640)
);

OAI21xp33_ASAP7_75t_L g641 ( 
.A1(n_631),
.A2(n_618),
.B(n_602),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_627),
.B(n_616),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_632),
.B(n_616),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_637),
.Y(n_644)
);

OAI211xp5_ASAP7_75t_L g645 ( 
.A1(n_641),
.A2(n_609),
.B(n_612),
.C(n_606),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_635),
.A2(n_603),
.B(n_620),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_640),
.B(n_610),
.Y(n_647)
);

NAND4xp25_ASAP7_75t_SL g648 ( 
.A(n_638),
.B(n_612),
.C(n_613),
.D(n_603),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_635),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_640),
.B(n_607),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_637),
.B(n_624),
.Y(n_651)
);

AOI222xp33_ASAP7_75t_L g652 ( 
.A1(n_634),
.A2(n_628),
.B1(n_607),
.B2(n_630),
.C1(n_622),
.C2(n_629),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_651),
.B(n_636),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_649),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_645),
.A2(n_636),
.B(n_626),
.Y(n_655)
);

O2A1O1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_646),
.A2(n_626),
.B(n_605),
.C(n_628),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_651),
.B(n_638),
.Y(n_657)
);

AO22x1_ASAP7_75t_L g658 ( 
.A1(n_655),
.A2(n_650),
.B1(n_644),
.B2(n_647),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_657),
.B(n_648),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_653),
.Y(n_660)
);

OAI211xp5_ASAP7_75t_L g661 ( 
.A1(n_659),
.A2(n_656),
.B(n_652),
.C(n_654),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_660),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_662),
.Y(n_663)
);

AND2x4_ASAP7_75t_SL g664 ( 
.A(n_662),
.B(n_639),
.Y(n_664)
);

AO22x2_ASAP7_75t_L g665 ( 
.A1(n_663),
.A2(n_661),
.B1(n_658),
.B2(n_625),
.Y(n_665)
);

NAND3xp33_ASAP7_75t_SL g666 ( 
.A(n_664),
.B(n_639),
.C(n_642),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_664),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_665),
.A2(n_622),
.B1(n_642),
.B2(n_643),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_668),
.A2(n_667),
.B1(n_666),
.B2(n_622),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_669),
.B(n_643),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_670),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_671),
.A2(n_615),
.B(n_622),
.Y(n_672)
);


endmodule