module real_aes_1928_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_828, n_50, n_89, n_829, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_828;
input n_50;
input n_89;
input n_829;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g536 ( .A(n_0), .B(n_221), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_1), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g149 ( .A(n_2), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_3), .B(n_515), .Y(n_552) );
NAND2xp33_ASAP7_75t_SL g592 ( .A(n_4), .B(n_170), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_5), .B(n_205), .Y(n_212) );
INVx1_ASAP7_75t_L g585 ( .A(n_6), .Y(n_585) );
INVx1_ASAP7_75t_L g192 ( .A(n_7), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g825 ( .A(n_8), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_9), .Y(n_280) );
AND2x2_ASAP7_75t_L g550 ( .A(n_10), .B(n_173), .Y(n_550) );
INVx2_ASAP7_75t_L g141 ( .A(n_11), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_12), .A2(n_105), .B1(n_817), .B2(n_826), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_13), .Y(n_122) );
INVx1_ASAP7_75t_L g222 ( .A(n_14), .Y(n_222) );
AOI221x1_ASAP7_75t_L g588 ( .A1(n_15), .A2(n_138), .B1(n_517), .B2(n_589), .C(n_591), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_16), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g125 ( .A(n_17), .Y(n_125) );
INVx1_ASAP7_75t_L g219 ( .A(n_18), .Y(n_219) );
INVx1_ASAP7_75t_SL g234 ( .A(n_19), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_20), .B(n_164), .Y(n_208) );
AOI33xp33_ASAP7_75t_L g184 ( .A1(n_21), .A2(n_54), .A3(n_146), .B1(n_157), .B2(n_185), .B3(n_186), .Y(n_184) );
AOI221xp5_ASAP7_75t_SL g526 ( .A1(n_22), .A2(n_45), .B1(n_515), .B2(n_517), .C(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_23), .A2(n_517), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_24), .B(n_221), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_25), .A2(n_38), .B1(n_799), .B2(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_25), .Y(n_800) );
INVx1_ASAP7_75t_L g274 ( .A(n_26), .Y(n_274) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_27), .A2(n_92), .B(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g174 ( .A(n_27), .B(n_92), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_28), .B(n_224), .Y(n_520) );
INVxp67_ASAP7_75t_L g587 ( .A(n_29), .Y(n_587) );
AND2x2_ASAP7_75t_L g574 ( .A(n_30), .B(n_172), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_31), .B(n_144), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_32), .A2(n_517), .B(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_33), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_34), .B(n_377), .Y(n_376) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_34), .Y(n_500) );
OAI22x1_ASAP7_75t_R g802 ( .A1(n_34), .A2(n_40), .B1(n_500), .B2(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_35), .B(n_224), .Y(n_528) );
AND2x2_ASAP7_75t_L g151 ( .A(n_36), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g156 ( .A(n_36), .Y(n_156) );
AND2x2_ASAP7_75t_L g170 ( .A(n_36), .B(n_149), .Y(n_170) );
OR2x6_ASAP7_75t_L g123 ( .A(n_37), .B(n_124), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_38), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_39), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_40), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_41), .B(n_144), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_42), .A2(n_139), .B1(n_201), .B2(n_205), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_43), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_43), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_44), .B(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_46), .B(n_164), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_47), .A2(n_84), .B1(n_154), .B2(n_517), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_48), .B(n_221), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_49), .B(n_179), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_50), .B(n_164), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_51), .Y(n_204) );
AND2x2_ASAP7_75t_L g539 ( .A(n_52), .B(n_172), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_53), .B(n_172), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_55), .B(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g147 ( .A(n_56), .Y(n_147) );
INVx1_ASAP7_75t_L g166 ( .A(n_56), .Y(n_166) );
AND2x2_ASAP7_75t_L g171 ( .A(n_57), .B(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_58), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g190 ( .A1(n_59), .A2(n_77), .B1(n_144), .B2(n_154), .C(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_60), .B(n_144), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_61), .B(n_515), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_62), .B(n_139), .Y(n_282) );
AOI21xp5_ASAP7_75t_SL g242 ( .A1(n_63), .A2(n_154), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g565 ( .A(n_64), .B(n_172), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_65), .B(n_224), .Y(n_537) );
INVx1_ASAP7_75t_L g215 ( .A(n_66), .Y(n_215) );
AND2x2_ASAP7_75t_SL g521 ( .A(n_67), .B(n_173), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_68), .B(n_221), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_69), .A2(n_517), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g161 ( .A(n_70), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_71), .B(n_224), .Y(n_556) );
AND2x2_ASAP7_75t_SL g547 ( .A(n_72), .B(n_179), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_73), .A2(n_154), .B(n_160), .Y(n_153) );
OAI22xp5_ASAP7_75t_SL g116 ( .A1(n_74), .A2(n_96), .B1(n_117), .B2(n_118), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_74), .Y(n_117) );
INVx1_ASAP7_75t_L g152 ( .A(n_75), .Y(n_152) );
INVx1_ASAP7_75t_L g168 ( .A(n_75), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_76), .B(n_144), .Y(n_187) );
AND2x2_ASAP7_75t_L g236 ( .A(n_78), .B(n_138), .Y(n_236) );
INVx1_ASAP7_75t_L g216 ( .A(n_79), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_80), .A2(n_154), .B(n_233), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_81), .A2(n_154), .B(n_178), .C(n_207), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_82), .A2(n_87), .B1(n_144), .B2(n_515), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_83), .B(n_515), .Y(n_564) );
INVx1_ASAP7_75t_L g126 ( .A(n_85), .Y(n_126) );
AND2x2_ASAP7_75t_SL g240 ( .A(n_86), .B(n_138), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_88), .A2(n_154), .B1(n_182), .B2(n_183), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_89), .B(n_221), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_90), .B(n_221), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_91), .A2(n_517), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g244 ( .A(n_93), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_94), .B(n_224), .Y(n_562) );
AND2x2_ASAP7_75t_L g188 ( .A(n_95), .B(n_138), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_96), .Y(n_118) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_97), .A2(n_272), .B(n_273), .C(n_275), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_98), .B(n_515), .Y(n_538) );
INVxp67_ASAP7_75t_L g590 ( .A(n_99), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_100), .B(n_224), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_101), .A2(n_517), .B(n_518), .Y(n_516) );
BUFx2_ASAP7_75t_L g110 ( .A(n_102), .Y(n_110) );
BUFx2_ASAP7_75t_SL g796 ( .A(n_102), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_103), .B(n_164), .Y(n_245) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_794), .B(n_812), .Y(n_105) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_111), .C(n_785), .Y(n_106) );
CKINVDCx11_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2x1_ASAP7_75t_R g810 ( .A(n_110), .B(n_811), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_119), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_113), .A2(n_786), .B(n_789), .Y(n_785) );
INVxp33_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_127), .B1(n_502), .B2(n_506), .Y(n_119) );
OAI21x1_ASAP7_75t_L g786 ( .A1(n_120), .A2(n_787), .B(n_788), .Y(n_786) );
CKINVDCx11_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
AND2x6_ASAP7_75t_SL g121 ( .A(n_122), .B(n_123), .Y(n_121) );
OR2x6_ASAP7_75t_SL g504 ( .A(n_122), .B(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g793 ( .A(n_122), .B(n_123), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_122), .B(n_505), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_123), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
INVx2_ASAP7_75t_L g787 ( .A(n_127), .Y(n_787) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_497), .Y(n_127) );
NOR4xp25_ASAP7_75t_L g128 ( .A(n_129), .B(n_376), .C(n_400), .D(n_466), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_129), .A2(n_400), .B1(n_500), .B2(n_828), .Y(n_501) );
INVx2_ASAP7_75t_L g807 ( .A(n_129), .Y(n_807) );
NAND3x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_328), .C(n_362), .Y(n_129) );
NOR3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_287), .C(n_307), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_262), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_195), .B1(n_251), .B2(n_259), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_175), .Y(n_133) );
AND2x2_ASAP7_75t_L g426 ( .A(n_134), .B(n_356), .Y(n_426) );
INVx1_ASAP7_75t_L g433 ( .A(n_134), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_134), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_134), .B(n_296), .Y(n_485) );
OR2x2_ASAP7_75t_L g495 ( .A(n_134), .B(n_496), .Y(n_495) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_135), .B(n_253), .Y(n_316) );
AND2x4_ASAP7_75t_L g344 ( .A(n_135), .B(n_258), .Y(n_344) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g292 ( .A(n_136), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_136), .B(n_177), .Y(n_382) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_136), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_136), .B(n_269), .Y(n_419) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_142), .B(n_171), .Y(n_136) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_137), .A2(n_142), .B(n_171), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_137), .A2(n_138), .B1(n_271), .B2(n_276), .Y(n_270) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_139), .B(n_279), .Y(n_278) );
AOI21x1_ASAP7_75t_L g532 ( .A1(n_139), .A2(n_533), .B(n_539), .Y(n_532) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_140), .Y(n_179) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_141), .B(n_174), .Y(n_173) );
AND2x4_ASAP7_75t_L g205 ( .A(n_141), .B(n_174), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_153), .Y(n_142) );
INVx1_ASAP7_75t_L g283 ( .A(n_144), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_144), .A2(n_154), .B1(n_584), .B2(n_586), .Y(n_583) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_150), .Y(n_144) );
INVx1_ASAP7_75t_L g202 ( .A(n_145), .Y(n_202) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
OR2x6_ASAP7_75t_L g162 ( .A(n_146), .B(n_158), .Y(n_162) );
INVxp33_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g159 ( .A(n_147), .B(n_149), .Y(n_159) );
AND2x4_ASAP7_75t_L g224 ( .A(n_147), .B(n_167), .Y(n_224) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g203 ( .A(n_150), .Y(n_203) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g517 ( .A(n_151), .B(n_159), .Y(n_517) );
INVx2_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
AND2x6_ASAP7_75t_L g221 ( .A(n_152), .B(n_165), .Y(n_221) );
INVxp67_ASAP7_75t_L g281 ( .A(n_154), .Y(n_281) );
AND2x4_ASAP7_75t_L g154 ( .A(n_155), .B(n_159), .Y(n_154) );
NOR2x1p5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx1_ASAP7_75t_L g186 ( .A(n_157), .Y(n_186) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_163), .C(n_169), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_SL g191 ( .A1(n_162), .A2(n_169), .B(n_192), .C(n_193), .Y(n_191) );
INVx2_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_162), .A2(n_215), .B1(n_216), .B2(n_217), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g233 ( .A1(n_162), .A2(n_169), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_162), .A2(n_169), .B(n_244), .C(n_245), .Y(n_243) );
INVxp67_ASAP7_75t_L g272 ( .A(n_162), .Y(n_272) );
INVx1_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
AND2x4_ASAP7_75t_L g515 ( .A(n_164), .B(n_170), .Y(n_515) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_167), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g182 ( .A(n_169), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_169), .A2(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_169), .B(n_205), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_169), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_169), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_169), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_169), .A2(n_555), .B(n_556), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_169), .A2(n_562), .B(n_563), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_169), .A2(n_571), .B(n_572), .Y(n_570) );
INVx5_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_170), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_172), .Y(n_229) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_172), .A2(n_526), .B(n_530), .Y(n_525) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_175), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g490 ( .A(n_175), .B(n_327), .Y(n_490) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OR2x2_ASAP7_75t_L g480 ( .A(n_176), .B(n_419), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_189), .Y(n_176) );
INVx2_ASAP7_75t_L g258 ( .A(n_177), .Y(n_258) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_180), .B(n_188), .Y(n_177) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_178), .A2(n_180), .B(n_188), .Y(n_286) );
AOI21x1_ASAP7_75t_L g543 ( .A1(n_178), .A2(n_544), .B(n_547), .Y(n_543) );
INVx2_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_179), .A2(n_190), .B(n_194), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_179), .A2(n_514), .B(n_516), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_181), .B(n_187), .Y(n_180) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
INVx2_ASAP7_75t_L g268 ( .A(n_189), .Y(n_268) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_189), .Y(n_293) );
INVx1_ASAP7_75t_L g306 ( .A(n_189), .Y(n_306) );
INVxp67_ASAP7_75t_L g325 ( .A(n_189), .Y(n_325) );
AND2x4_ASAP7_75t_L g356 ( .A(n_189), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_237), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_226), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g398 ( .A(n_198), .B(n_385), .Y(n_398) );
AND2x2_ASAP7_75t_L g422 ( .A(n_198), .B(n_238), .Y(n_422) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_211), .Y(n_198) );
INVx2_ASAP7_75t_L g250 ( .A(n_199), .Y(n_250) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_199), .Y(n_265) );
INVx1_ASAP7_75t_L g322 ( .A(n_199), .Y(n_322) );
AND2x4_ASAP7_75t_L g331 ( .A(n_199), .B(n_249), .Y(n_331) );
AND2x2_ASAP7_75t_L g387 ( .A(n_199), .B(n_239), .Y(n_387) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_206), .Y(n_199) );
NOR3xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .C(n_204), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_205), .A2(n_242), .B(n_246), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_205), .A2(n_552), .B(n_553), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_205), .B(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_205), .B(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_205), .B(n_590), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_205), .B(n_217), .C(n_592), .Y(n_591) );
INVx3_ASAP7_75t_L g249 ( .A(n_211), .Y(n_249) );
AND2x2_ASAP7_75t_L g261 ( .A(n_211), .B(n_228), .Y(n_261) );
INVx2_ASAP7_75t_L g300 ( .A(n_211), .Y(n_300) );
NOR2x1_ASAP7_75t_SL g313 ( .A(n_211), .B(n_239), .Y(n_313) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_218), .B(n_225), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_217), .B(n_274), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B1(n_222), .B2(n_223), .Y(n_218) );
INVxp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVxp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g415 ( .A(n_226), .Y(n_415) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g338 ( .A(n_227), .Y(n_338) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_228), .Y(n_296) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_228), .Y(n_312) );
AND2x2_ASAP7_75t_L g320 ( .A(n_228), .B(n_249), .Y(n_320) );
INVx1_ASAP7_75t_L g360 ( .A(n_228), .Y(n_360) );
INVx1_ASAP7_75t_L g385 ( .A(n_228), .Y(n_385) );
OR2x2_ASAP7_75t_L g446 ( .A(n_228), .B(n_239), .Y(n_446) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_236), .Y(n_228) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_229), .A2(n_559), .B(n_565), .Y(n_558) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_229), .A2(n_568), .B(n_574), .Y(n_567) );
AO21x2_ASAP7_75t_L g612 ( .A1(n_229), .A2(n_568), .B(n_574), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
OA211x2_ASAP7_75t_L g467 ( .A1(n_237), .A2(n_468), .B(n_470), .C(n_477), .Y(n_467) );
OR2x6_ASAP7_75t_L g237 ( .A(n_238), .B(n_247), .Y(n_237) );
AND2x2_ASAP7_75t_L g388 ( .A(n_238), .B(n_261), .Y(n_388) );
AND2x2_ASAP7_75t_SL g406 ( .A(n_238), .B(n_248), .Y(n_406) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx4_ASAP7_75t_L g260 ( .A(n_239), .Y(n_260) );
INVx2_ASAP7_75t_L g302 ( .A(n_239), .Y(n_302) );
AND2x4_ASAP7_75t_L g365 ( .A(n_239), .B(n_322), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_239), .B(n_361), .Y(n_416) );
AND2x2_ASAP7_75t_L g459 ( .A(n_239), .B(n_300), .Y(n_459) );
OR2x6_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_248), .B(n_360), .Y(n_453) );
AND2x2_ASAP7_75t_L g473 ( .A(n_248), .B(n_296), .Y(n_473) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g361 ( .A(n_249), .Y(n_361) );
INVx1_ASAP7_75t_L g335 ( .A(n_250), .Y(n_335) );
NOR2xp67_ASAP7_75t_SL g251 ( .A(n_252), .B(n_255), .Y(n_251) );
INVx1_ASAP7_75t_L g429 ( .A(n_252), .Y(n_429) );
NOR2xp67_ASAP7_75t_L g476 ( .A(n_252), .B(n_430), .Y(n_476) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g449 ( .A(n_254), .B(n_291), .Y(n_449) );
OAI211xp5_ASAP7_75t_L g437 ( .A1(n_255), .A2(n_438), .B(n_441), .C(n_450), .Y(n_437) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_255), .A2(n_475), .B(n_482), .C(n_486), .Y(n_481) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g366 ( .A(n_256), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g285 ( .A(n_257), .Y(n_285) );
NOR2x1_ASAP7_75t_L g305 ( .A(n_257), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g341 ( .A(n_257), .B(n_291), .Y(n_341) );
NOR2xp67_ASAP7_75t_L g451 ( .A(n_257), .B(n_291), .Y(n_451) );
AND2x2_ASAP7_75t_L g324 ( .A(n_258), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g375 ( .A(n_258), .Y(n_375) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x4_ASAP7_75t_SL g264 ( .A(n_260), .B(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g321 ( .A(n_260), .B(n_322), .Y(n_321) );
NOR2x1_ASAP7_75t_L g350 ( .A(n_260), .B(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g369 ( .A(n_260), .B(n_370), .Y(n_369) );
NOR2xp67_ASAP7_75t_SL g452 ( .A(n_260), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_SL g263 ( .A(n_261), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_261), .B(n_334), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx2_ASAP7_75t_SL g460 ( .A(n_266), .Y(n_460) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_284), .Y(n_266) );
INVx3_ASAP7_75t_L g383 ( .A(n_267), .Y(n_383) );
AND2x2_ASAP7_75t_L g404 ( .A(n_267), .B(n_395), .Y(n_404) );
AND2x2_ASAP7_75t_L g462 ( .A(n_267), .B(n_344), .Y(n_462) );
AND2x4_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx2_ASAP7_75t_L g291 ( .A(n_269), .Y(n_291) );
INVx1_ASAP7_75t_L g327 ( .A(n_269), .Y(n_327) );
INVx1_ASAP7_75t_L g347 ( .A(n_269), .Y(n_347) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_277), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .B1(n_282), .B2(n_283), .Y(n_277) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g430 ( .A(n_284), .Y(n_430) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g290 ( .A(n_286), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g357 ( .A(n_286), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_294), .B1(n_297), .B2(n_303), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
AND2x2_ASAP7_75t_L g304 ( .A(n_290), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g315 ( .A(n_290), .Y(n_315) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g364 ( .A(n_295), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVxp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g384 ( .A(n_299), .B(n_385), .Y(n_384) );
NOR2x1_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g392 ( .A(n_300), .Y(n_392) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g440 ( .A(n_302), .B(n_331), .Y(n_440) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_304), .A2(n_398), .B(n_399), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_314), .B(n_317), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g363 ( .A(n_313), .B(n_337), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_314), .A2(n_421), .B1(n_423), .B2(n_425), .Y(n_420) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_323), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_SL g370 ( .A(n_320), .Y(n_370) );
AND2x2_ASAP7_75t_L g399 ( .A(n_321), .B(n_337), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_321), .B(n_359), .Y(n_431) );
AND2x2_ASAP7_75t_L g435 ( .A(n_321), .B(n_392), .Y(n_435) );
OAI21xp5_ASAP7_75t_SL g379 ( .A1(n_323), .A2(n_380), .B(n_384), .Y(n_379) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
AND2x2_ASAP7_75t_L g340 ( .A(n_324), .B(n_341), .Y(n_340) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_324), .B(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g409 ( .A(n_327), .Y(n_409) );
NOR2x1_ASAP7_75t_L g328 ( .A(n_329), .B(n_352), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_339), .B1(n_342), .B2(n_348), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx4_ASAP7_75t_L g351 ( .A(n_331), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_331), .B(n_337), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_331), .B(n_484), .Y(n_483) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_334), .A2(n_358), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g457 ( .A(n_334), .B(n_359), .Y(n_457) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g439 ( .A(n_336), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g475 ( .A(n_337), .B(n_459), .Y(n_475) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g355 ( .A(n_341), .B(n_356), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_341), .B(n_375), .Y(n_374) );
OAI22xp5_ASAP7_75t_SL g352 ( .A1(n_342), .A2(n_353), .B1(n_354), .B2(n_358), .Y(n_352) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g469 ( .A(n_346), .B(n_356), .Y(n_469) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g367 ( .A(n_347), .Y(n_367) );
AND2x2_ASAP7_75t_L g393 ( .A(n_347), .B(n_356), .Y(n_393) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_349), .B(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_350), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g444 ( .A(n_351), .Y(n_444) );
INVx1_ASAP7_75t_L g456 ( .A(n_353), .Y(n_456) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_355), .A2(n_399), .B1(n_478), .B2(n_479), .Y(n_477) );
AND2x2_ASAP7_75t_L g394 ( .A(n_356), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g465 ( .A(n_356), .B(n_418), .Y(n_465) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI211xp5_ASAP7_75t_SL g368 ( .A1(n_359), .A2(n_369), .B(n_371), .C(n_372), .Y(n_368) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_359), .B(n_365), .Y(n_478) );
AND2x4_ASAP7_75t_SL g359 ( .A(n_360), .B(n_361), .Y(n_359) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_360), .Y(n_412) );
O2A1O1Ixp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B(n_366), .C(n_368), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_363), .A2(n_391), .B1(n_393), .B2(n_394), .Y(n_390) );
INVx2_ASAP7_75t_L g371 ( .A(n_365), .Y(n_371) );
AND2x2_ASAP7_75t_L g391 ( .A(n_365), .B(n_392), .Y(n_391) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_365), .Y(n_458) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g499 ( .A(n_377), .Y(n_499) );
NAND4xp75_ASAP7_75t_L g804 ( .A(n_377), .B(n_805), .C(n_806), .D(n_807), .Y(n_804) );
NOR2x1_ASAP7_75t_SL g377 ( .A(n_378), .B(n_389), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_386), .Y(n_378) );
OAI21xp5_ASAP7_75t_L g386 ( .A1(n_380), .A2(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g410 ( .A(n_382), .Y(n_410) );
INVx1_ASAP7_75t_L g486 ( .A(n_383), .Y(n_486) );
AND2x2_ASAP7_75t_L g424 ( .A(n_387), .B(n_412), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_388), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_390), .B(n_397), .Y(n_389) );
AND2x2_ASAP7_75t_L g491 ( .A(n_393), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g805 ( .A(n_400), .Y(n_805) );
NAND2x1_ASAP7_75t_L g400 ( .A(n_401), .B(n_436), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_420), .C(n_427), .Y(n_401) );
OAI222xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_405), .B1(n_407), .B2(n_411), .C1(n_413), .C2(n_417), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NOR2x1_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g463 ( .A(n_422), .Y(n_463) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_431), .B1(n_432), .B2(n_434), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NOR2xp67_ASAP7_75t_SL g436 ( .A(n_437), .B(n_454), .Y(n_436) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_447), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_444), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g496 ( .A(n_449), .Y(n_496) );
NAND2xp33_ASAP7_75t_SL g450 ( .A(n_451), .B(n_452), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_460), .B1(n_461), .B2(n_463), .C(n_464), .Y(n_454) );
NOR4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .C(n_458), .D(n_459), .Y(n_455) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_466), .A2(n_499), .B(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g806 ( .A(n_466), .Y(n_806) );
NAND4xp75_ASAP7_75t_L g466 ( .A(n_467), .B(n_481), .C(n_487), .D(n_493), .Y(n_466) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_471), .B(n_476), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NOR2x1_ASAP7_75t_L g487 ( .A(n_488), .B(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
NAND2x1_ASAP7_75t_SL g788 ( .A(n_503), .B(n_506), .Y(n_788) );
CKINVDCx11_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_677), .Y(n_507) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_605), .C(n_655), .Y(n_508) );
OAI211xp5_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_540), .B(n_575), .C(n_594), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_522), .Y(n_510) );
AND2x2_ASAP7_75t_L g604 ( .A(n_511), .B(n_523), .Y(n_604) );
INVx1_ASAP7_75t_L g735 ( .A(n_511), .Y(n_735) );
NOR2x1p5_ASAP7_75t_L g767 ( .A(n_511), .B(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g580 ( .A(n_512), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g626 ( .A(n_512), .Y(n_626) );
OR2x2_ASAP7_75t_L g630 ( .A(n_512), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_512), .B(n_525), .Y(n_642) );
OR2x2_ASAP7_75t_L g664 ( .A(n_512), .B(n_525), .Y(n_664) );
AND2x4_ASAP7_75t_L g670 ( .A(n_512), .B(n_634), .Y(n_670) );
OR2x2_ASAP7_75t_L g687 ( .A(n_512), .B(n_582), .Y(n_687) );
INVx1_ASAP7_75t_L g722 ( .A(n_512), .Y(n_722) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_512), .Y(n_744) );
OR2x2_ASAP7_75t_L g758 ( .A(n_512), .B(n_691), .Y(n_758) );
AND2x4_ASAP7_75t_SL g762 ( .A(n_512), .B(n_582), .Y(n_762) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_521), .Y(n_512) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g714 ( .A(n_523), .B(n_670), .Y(n_714) );
AND2x2_ASAP7_75t_L g761 ( .A(n_523), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_531), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g579 ( .A(n_525), .Y(n_579) );
AND2x2_ASAP7_75t_L g624 ( .A(n_525), .B(n_531), .Y(n_624) );
INVx2_ASAP7_75t_L g631 ( .A(n_525), .Y(n_631) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_525), .Y(n_752) );
BUFx3_ASAP7_75t_L g768 ( .A(n_525), .Y(n_768) );
INVx2_ASAP7_75t_L g593 ( .A(n_531), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_531), .B(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g691 ( .A(n_531), .B(n_631), .Y(n_691) );
INVx1_ASAP7_75t_L g709 ( .A(n_531), .Y(n_709) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_531), .Y(n_725) );
INVx1_ASAP7_75t_L g747 ( .A(n_531), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_531), .B(n_626), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_531), .B(n_582), .Y(n_784) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_548), .Y(n_541) );
AND2x4_ASAP7_75t_L g598 ( .A(n_542), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g609 ( .A(n_542), .Y(n_609) );
AND2x2_ASAP7_75t_L g614 ( .A(n_542), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g649 ( .A(n_542), .B(n_557), .Y(n_649) );
AND2x2_ASAP7_75t_L g659 ( .A(n_542), .B(n_558), .Y(n_659) );
OR2x2_ASAP7_75t_L g739 ( .A(n_542), .B(n_654), .Y(n_739) );
OAI322xp33_ASAP7_75t_L g769 ( .A1(n_542), .A2(n_682), .A3(n_721), .B1(n_754), .B2(n_770), .C1(n_771), .C2(n_772), .Y(n_769) );
OR2x2_ASAP7_75t_L g770 ( .A(n_542), .B(n_752), .Y(n_770) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g603 ( .A(n_543), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_548), .A2(n_716), .B1(n_720), .B2(n_723), .Y(n_715) );
AOI211xp5_ASAP7_75t_L g775 ( .A1(n_548), .A2(n_776), .B(n_777), .C(n_780), .Y(n_775) );
AND2x4_ASAP7_75t_SL g548 ( .A(n_549), .B(n_557), .Y(n_548) );
AND2x4_ASAP7_75t_L g597 ( .A(n_549), .B(n_567), .Y(n_597) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_549), .Y(n_601) );
INVx5_ASAP7_75t_L g613 ( .A(n_549), .Y(n_613) );
INVx2_ASAP7_75t_L g622 ( .A(n_549), .Y(n_622) );
AND2x2_ASAP7_75t_L g645 ( .A(n_549), .B(n_558), .Y(n_645) );
AND2x2_ASAP7_75t_L g674 ( .A(n_549), .B(n_566), .Y(n_674) );
OR2x2_ASAP7_75t_L g683 ( .A(n_549), .B(n_603), .Y(n_683) );
OR2x2_ASAP7_75t_L g698 ( .A(n_549), .B(n_612), .Y(n_698) );
OR2x6_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_557), .B(n_576), .Y(n_575) );
INVx3_ASAP7_75t_SL g682 ( .A(n_557), .Y(n_682) );
AND2x2_ASAP7_75t_L g705 ( .A(n_557), .B(n_613), .Y(n_705) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_566), .Y(n_557) );
INVx2_ASAP7_75t_L g599 ( .A(n_558), .Y(n_599) );
AND2x2_ASAP7_75t_L g602 ( .A(n_558), .B(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g616 ( .A(n_558), .B(n_567), .Y(n_616) );
INVx1_ASAP7_75t_L g620 ( .A(n_558), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_558), .B(n_567), .Y(n_654) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_558), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_558), .B(n_613), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .Y(n_559) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_567), .Y(n_635) );
AND2x2_ASAP7_75t_L g719 ( .A(n_567), .B(n_603), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_573), .Y(n_568) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_577), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x6_ASAP7_75t_SL g783 ( .A(n_578), .B(n_784), .Y(n_783) );
INVxp67_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_579), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_579), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g731 ( .A(n_579), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_580), .A2(n_640), .B1(n_643), .B2(n_650), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_581), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g675 ( .A(n_581), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_581), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_SL g730 ( .A(n_581), .B(n_731), .Y(n_730) );
AND2x4_ASAP7_75t_L g581 ( .A(n_582), .B(n_593), .Y(n_581) );
AND2x2_ASAP7_75t_L g625 ( .A(n_582), .B(n_626), .Y(n_625) );
INVx3_ASAP7_75t_L g634 ( .A(n_582), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g692 ( .A1(n_582), .A2(n_641), .B1(n_693), .B2(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g700 ( .A(n_582), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_582), .B(n_694), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_582), .B(n_624), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_582), .B(n_631), .Y(n_773) );
AND2x4_ASAP7_75t_L g582 ( .A(n_583), .B(n_588), .Y(n_582) );
OAI21xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_600), .B(n_604), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
NAND4xp25_ASAP7_75t_SL g643 ( .A(n_596), .B(n_644), .C(n_646), .D(n_648), .Y(n_643) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_597), .B(n_704), .Y(n_733) );
AND2x2_ASAP7_75t_L g760 ( .A(n_597), .B(n_598), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_597), .B(n_620), .Y(n_771) );
INVx1_ASAP7_75t_L g636 ( .A(n_598), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_598), .A2(n_661), .B1(n_672), .B2(n_675), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_598), .B(n_611), .C(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_598), .B(n_613), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_598), .B(n_621), .Y(n_764) );
AND2x2_ASAP7_75t_L g696 ( .A(n_599), .B(n_603), .Y(n_696) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_599), .Y(n_757) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g652 ( .A(n_601), .Y(n_652) );
INVx1_ASAP7_75t_L g742 ( .A(n_602), .Y(n_742) );
AND2x2_ASAP7_75t_L g749 ( .A(n_602), .B(n_613), .Y(n_749) );
BUFx2_ASAP7_75t_L g704 ( .A(n_603), .Y(n_704) );
NAND3xp33_ASAP7_75t_SL g605 ( .A(n_606), .B(n_627), .C(n_639), .Y(n_605) );
OAI31xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_614), .A3(n_617), .B(n_623), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_607), .A2(n_661), .B1(n_665), .B2(n_666), .Y(n_660) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OR2x2_ASAP7_75t_L g646 ( .A(n_609), .B(n_647), .Y(n_646) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_609), .B(n_673), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g741 ( .A1(n_610), .A2(n_712), .B(n_742), .C(n_743), .Y(n_741) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_611), .B(n_757), .Y(n_756) );
AND2x4_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_612), .B(n_620), .Y(n_647) );
AND2x2_ASAP7_75t_L g665 ( .A(n_612), .B(n_645), .Y(n_665) );
AND2x2_ASAP7_75t_L g782 ( .A(n_615), .B(n_704), .Y(n_782) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g638 ( .A(n_616), .B(n_622), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_621), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_621), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g713 ( .A(n_621), .B(n_696), .Y(n_713) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_622), .B(n_696), .Y(n_702) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx2_ASAP7_75t_L g694 ( .A(n_624), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_625), .B(n_725), .Y(n_724) );
AOI32xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_635), .A3(n_636), .B1(n_637), .B2(n_829), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_628), .A2(n_713), .B1(n_749), .B2(n_750), .C(n_753), .Y(n_748) );
AND2x4_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_631), .Y(n_676) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g641 ( .A(n_633), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g746 ( .A(n_634), .B(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_635), .B(n_657), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_637), .A2(n_680), .B1(n_684), .B2(n_688), .C(n_692), .Y(n_679) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI211xp5_ASAP7_75t_L g655 ( .A1(n_642), .A2(n_656), .B(n_660), .C(n_671), .Y(n_655) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI322xp33_ASAP7_75t_L g753 ( .A1(n_648), .A2(n_658), .A3(n_707), .B1(n_754), .B2(n_755), .C1(n_756), .C2(n_758), .Y(n_753) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI21xp33_ASAP7_75t_L g780 ( .A1(n_651), .A2(n_781), .B(n_783), .Y(n_780) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_657), .A2(n_738), .B(n_740), .C(n_741), .Y(n_737) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g779 ( .A(n_664), .B(n_745), .Y(n_779) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_670), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g754 ( .A(n_670), .Y(n_754) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI31xp33_ASAP7_75t_L g710 ( .A1(n_674), .A2(n_711), .A3(n_713), .B(n_714), .Y(n_710) );
NOR2x1_ASAP7_75t_L g677 ( .A(n_678), .B(n_736), .Y(n_677) );
NAND5xp2_ASAP7_75t_L g678 ( .A(n_679), .B(n_699), .C(n_710), .D(n_715), .E(n_726), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
AOI21xp33_ASAP7_75t_L g777 ( .A1(n_682), .A2(n_778), .B(n_779), .Y(n_777) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g750 ( .A(n_686), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B(n_703), .C(n_706), .Y(n_699) );
INVxp33_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
OR2x2_ASAP7_75t_L g728 ( .A(n_704), .B(n_729), .Y(n_728) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_707), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_SL g716 ( .A(n_717), .B(n_719), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g778 ( .A(n_719), .Y(n_778) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_730), .B(n_732), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_728), .A2(n_733), .B(n_734), .Y(n_732) );
NAND4xp25_ASAP7_75t_L g736 ( .A(n_737), .B(n_748), .C(n_759), .D(n_775), .Y(n_736) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_746), .B(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g776 ( .A(n_758), .Y(n_776) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_763), .B2(n_765), .C(n_769), .Y(n_759) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OR2x2_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx1_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_797), .B(n_810), .Y(n_794) );
CKINVDCx8_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_801), .B1(n_808), .B2(n_809), .Y(n_797) );
INVx1_ASAP7_75t_L g809 ( .A(n_798), .Y(n_809) );
INVx2_ASAP7_75t_L g808 ( .A(n_801), .Y(n_808) );
XNOR2x1_ASAP7_75t_L g801 ( .A(n_802), .B(n_804), .Y(n_801) );
BUFx3_ASAP7_75t_L g816 ( .A(n_811), .Y(n_816) );
BUFx2_ASAP7_75t_L g822 ( .A(n_811), .Y(n_822) );
NOR2x1_ASAP7_75t_R g812 ( .A(n_813), .B(n_814), .Y(n_812) );
CKINVDCx11_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_819), .Y(n_826) );
INVx2_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_SL g820 ( .A(n_821), .B(n_823), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
endmodule