module fake_netlist_6_3821_n_3760 (n_992, n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_968, n_909, n_580, n_762, n_1030, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_1008, n_1027, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_1033, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_933, n_740, n_1038, n_578, n_703, n_1003, n_144, n_365, n_978, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_1044, n_951, n_783, n_106, n_725, n_952, n_999, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_994, n_677, n_969, n_988, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_974, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_1020, n_180, n_1009, n_1042, n_62, n_628, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_1032, n_845, n_255, n_807, n_1036, n_739, n_284, n_400, n_140, n_337, n_955, n_865, n_893, n_214, n_925, n_485, n_67, n_15, n_1026, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_935, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_963, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_1024, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_1018, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_1037, n_72, n_721, n_996, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_1015, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_56, n_763, n_1057, n_360, n_945, n_977, n_603, n_1005, n_119, n_991, n_957, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_971, n_946, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_987, n_641, n_822, n_693, n_1056, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_943, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_989, n_797, n_666, n_1016, n_371, n_795, n_770, n_940, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_1035, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_953, n_20, n_1004, n_1017, n_494, n_539, n_493, n_397, n_155, n_1022, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_1049, n_576, n_1028, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_976, n_490, n_803, n_290, n_220, n_809, n_1043, n_1011, n_118, n_224, n_48, n_926, n_927, n_25, n_93, n_839, n_986, n_80, n_734, n_708, n_196, n_919, n_402, n_352, n_917, n_668, n_478, n_626, n_990, n_574, n_779, n_9, n_800, n_929, n_460, n_107, n_907, n_854, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_921, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_293, n_1054, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_998, n_16, n_1046, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_924, n_298, n_18, n_492, n_972, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_962, n_1000, n_279, n_686, n_796, n_1041, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_936, n_184, n_552, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_984, n_411, n_503, n_716, n_152, n_623, n_1048, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_1021, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_958, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_942, n_792, n_880, n_476, n_981, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_985, n_589, n_860, n_481, n_788, n_819, n_939, n_997, n_821, n_325, n_938, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_964, n_982, n_561, n_33, n_477, n_549, n_980, n_533, n_954, n_408, n_932, n_806, n_864, n_879, n_959, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_979, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_993, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_1051, n_583, n_596, n_123, n_136, n_966, n_546, n_562, n_249, n_201, n_386, n_764, n_1039, n_556, n_159, n_1034, n_157, n_162, n_692, n_733, n_754, n_941, n_975, n_1031, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_970, n_560, n_1014, n_753, n_642, n_995, n_276, n_569, n_441, n_221, n_811, n_882, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_973, n_346, n_88, n_3, n_416, n_1053, n_530, n_277, n_520, n_1029, n_418, n_113, n_618, n_1055, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_967, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_1047, n_1010, n_355, n_426, n_317, n_149, n_1040, n_915, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_1052, n_502, n_328, n_672, n_534, n_488, n_429, n_1006, n_373, n_1012, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_1045, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_1002, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_1019, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_965, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_983, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_961, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_950, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_956, n_960, n_531, n_827, n_1001, n_60, n_361, n_508, n_663, n_856, n_1050, n_379, n_170, n_778, n_1025, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_1013, n_1023, n_194, n_664, n_171, n_949, n_678, n_192, n_57, n_169, n_1007, n_51, n_649, n_283, n_3760);

input n_992;
input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_968;
input n_909;
input n_580;
input n_762;
input n_1030;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_1008;
input n_1027;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_1033;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_933;
input n_740;
input n_1038;
input n_578;
input n_703;
input n_1003;
input n_144;
input n_365;
input n_978;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_1044;
input n_951;
input n_783;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_994;
input n_677;
input n_969;
input n_988;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_974;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_1020;
input n_180;
input n_1009;
input n_1042;
input n_62;
input n_628;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_1032;
input n_845;
input n_255;
input n_807;
input n_1036;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_955;
input n_865;
input n_893;
input n_214;
input n_925;
input n_485;
input n_67;
input n_15;
input n_1026;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_935;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_963;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_1024;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_1018;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_1037;
input n_72;
input n_721;
input n_996;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_1015;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_56;
input n_763;
input n_1057;
input n_360;
input n_945;
input n_977;
input n_603;
input n_1005;
input n_119;
input n_991;
input n_957;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_971;
input n_946;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_987;
input n_641;
input n_822;
input n_693;
input n_1056;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_943;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_989;
input n_797;
input n_666;
input n_1016;
input n_371;
input n_795;
input n_770;
input n_940;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_1035;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_953;
input n_20;
input n_1004;
input n_1017;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_1022;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_1049;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_976;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_1043;
input n_1011;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_25;
input n_93;
input n_839;
input n_986;
input n_80;
input n_734;
input n_708;
input n_196;
input n_919;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_990;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_921;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_293;
input n_1054;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_998;
input n_16;
input n_1046;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_18;
input n_492;
input n_972;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_962;
input n_1000;
input n_279;
input n_686;
input n_796;
input n_1041;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_984;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_1048;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_958;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_981;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_985;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_939;
input n_997;
input n_821;
input n_325;
input n_938;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_964;
input n_982;
input n_561;
input n_33;
input n_477;
input n_549;
input n_980;
input n_533;
input n_954;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_959;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_979;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_993;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_1051;
input n_583;
input n_596;
input n_123;
input n_136;
input n_966;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_1039;
input n_556;
input n_159;
input n_1034;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_970;
input n_560;
input n_1014;
input n_753;
input n_642;
input n_995;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_973;
input n_346;
input n_88;
input n_3;
input n_416;
input n_1053;
input n_530;
input n_277;
input n_520;
input n_1029;
input n_418;
input n_113;
input n_618;
input n_1055;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_967;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_1047;
input n_1010;
input n_355;
input n_426;
input n_317;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_1052;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_1006;
input n_373;
input n_1012;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_1045;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_1002;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_1019;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_965;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_983;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_961;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_950;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_956;
input n_960;
input n_531;
input n_827;
input n_1001;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_1050;
input n_379;
input n_170;
input n_778;
input n_1025;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_1013;
input n_1023;
input n_194;
input n_664;
input n_171;
input n_949;
input n_678;
input n_192;
input n_57;
input n_169;
input n_1007;
input n_51;
input n_649;
input n_283;

output n_3760;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1674;
wire n_1199;
wire n_3392;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_3152;
wire n_3579;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_1581;
wire n_1237;
wire n_1061;
wire n_2534;
wire n_2353;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_3741;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_3465;
wire n_1975;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_3706;
wire n_1160;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_1285;
wire n_2974;
wire n_2886;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_3232;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_3316;
wire n_2212;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_3107;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_3368;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_1446;
wire n_2591;
wire n_3507;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_1658;
wire n_2593;
wire n_3506;
wire n_3568;
wire n_3269;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_1193;
wire n_1967;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_1530;
wire n_3488;
wire n_1543;
wire n_2811;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_3317;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_3716;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1605;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_1726;
wire n_1950;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3247;
wire n_3069;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_3346;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3298;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_3691;
wire n_2624;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_1801;
wire n_1214;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2519;
wire n_2319;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_1630;
wire n_2887;
wire n_3500;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_3545;
wire n_1369;
wire n_3578;
wire n_2271;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3337;
wire n_3450;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1627;
wire n_1164;
wire n_1295;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_3614;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_1952;
wire n_3616;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_3436;
wire n_1932;
wire n_1101;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_2767;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_1514;
wire n_1863;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1139;
wire n_1714;
wire n_3179;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_2897;
wire n_2537;
wire n_2554;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_3608;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_2339;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3426;
wire n_3158;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3435;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3537;
wire n_2134;
wire n_1176;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_2231;
wire n_3609;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_3693;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_3200;
wire n_1665;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_3656;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_1073;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_2481;
wire n_3561;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2424;
wire n_2296;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_1142;
wire n_2849;
wire n_1774;
wire n_1475;
wire n_1398;
wire n_1201;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_3393;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_3641;
wire n_1314;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_2475;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_2990;
wire n_1773;
wire n_1775;
wire n_1286;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3364;
wire n_3323;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3425;
wire n_2384;
wire n_1745;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_3547;
wire n_1901;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_2829;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_1869;
wire n_3625;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_2201;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3194;
wire n_3113;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_2924;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1669;
wire n_1403;
wire n_1852;
wire n_3548;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_3475;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3262;
wire n_3544;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_3692;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_3597;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_1637;
wire n_2635;
wire n_3439;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_3712;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_3074;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_2154;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3469;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_3149;
wire n_3375;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_2128;
wire n_1794;
wire n_1650;
wire n_1962;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_3124;
wire n_1741;
wire n_1746;
wire n_1325;
wire n_1949;
wire n_3398;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_3711;
wire n_1727;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1800;
wire n_2241;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_3343;
wire n_3303;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_3652;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_1408;
wire n_3567;
wire n_1196;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_1848;
wire n_1785;
wire n_1114;
wire n_1147;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_3473;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1347;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_3215;
wire n_3336;
wire n_2952;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_2255;
wire n_2112;
wire n_1737;
wire n_1464;
wire n_2430;
wire n_3486;
wire n_1414;
wire n_3584;
wire n_2649;
wire n_2721;
wire n_3556;
wire n_2034;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_2444;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_1821;
wire n_1537;
wire n_1500;
wire n_2205;
wire n_3699;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_3378;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_3123;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_3038;
wire n_2033;
wire n_3086;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_3361;
wire n_3596;
wire n_3478;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_3310;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_3374;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_3552;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_2879;
wire n_3717;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_1170;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_3444;
wire n_2553;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_3527;
wire n_2512;
wire n_3433;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_1322;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_3504;
wire n_1449;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_69),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_994),
.Y(n_1059)
);

CKINVDCx16_ASAP7_75t_R g1060 ( 
.A(n_65),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_400),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_289),
.Y(n_1062)
);

CKINVDCx16_ASAP7_75t_R g1063 ( 
.A(n_387),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_255),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_390),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1012),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_930),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_1032),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_672),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_19),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_694),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_850),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_455),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_895),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_732),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_483),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_475),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_632),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_684),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1010),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_1027),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_430),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_916),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_416),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_329),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_827),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_270),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_676),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_981),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_60),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_691),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_656),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_347),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_501),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_403),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_565),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_570),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_6),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_779),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_66),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_261),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_414),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_552),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_849),
.Y(n_1104)
);

BUFx10_ASAP7_75t_L g1105 ( 
.A(n_239),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_301),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_914),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_181),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_974),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_697),
.Y(n_1110)
);

BUFx8_ASAP7_75t_SL g1111 ( 
.A(n_35),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_508),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_231),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_342),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_95),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_137),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_310),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_1015),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_71),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_874),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_704),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_9),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_815),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_936),
.Y(n_1124)
);

CKINVDCx14_ASAP7_75t_R g1125 ( 
.A(n_429),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_675),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_1024),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1052),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_789),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_821),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_681),
.Y(n_1131)
);

CKINVDCx16_ASAP7_75t_R g1132 ( 
.A(n_14),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_270),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_710),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_829),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_25),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_248),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_792),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_206),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1031),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_681),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_599),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_102),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_715),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_587),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_132),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1036),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_613),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_780),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_239),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_515),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_563),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_949),
.Y(n_1153)
);

BUFx10_ASAP7_75t_L g1154 ( 
.A(n_716),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_585),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_7),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_984),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_707),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_639),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_723),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_753),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_222),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_423),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_324),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_596),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_38),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_690),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_668),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_527),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1009),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_150),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_273),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1019),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_676),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_288),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_688),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_551),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_195),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_968),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_182),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_594),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_497),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_245),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_296),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_569),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_216),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_932),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1017),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_781),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_742),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_719),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_417),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_689),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_205),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_443),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_288),
.Y(n_1197)
);

BUFx10_ASAP7_75t_L g1198 ( 
.A(n_1025),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_828),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1041),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_519),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_18),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_251),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_566),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_364),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_0),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_699),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_43),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_112),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_695),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_476),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_650),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_686),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_261),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_837),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_937),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_131),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_204),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_245),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_592),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1049),
.Y(n_1221)
);

CKINVDCx14_ASAP7_75t_R g1222 ( 
.A(n_651),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_2),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_814),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_362),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_709),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_677),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_98),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_345),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_510),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_517),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_196),
.Y(n_1232)
);

BUFx10_ASAP7_75t_L g1233 ( 
.A(n_566),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_632),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_215),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1020),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_90),
.Y(n_1237)
);

CKINVDCx14_ASAP7_75t_R g1238 ( 
.A(n_929),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_982),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_75),
.Y(n_1240)
);

CKINVDCx16_ASAP7_75t_R g1241 ( 
.A(n_579),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_51),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1050),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1030),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_88),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_772),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_663),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_912),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_398),
.Y(n_1249)
);

BUFx8_ASAP7_75t_SL g1250 ( 
.A(n_1011),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_116),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_423),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_881),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_648),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_80),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_66),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_53),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_244),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_983),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_133),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_56),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_671),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_834),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_682),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_170),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_864),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_630),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_431),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_343),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_57),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1022),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_857),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_488),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_584),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_122),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1014),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_706),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_890),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_580),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_285),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1040),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_354),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_972),
.Y(n_1283)
);

INVxp67_ASAP7_75t_SL g1284 ( 
.A(n_686),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_541),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_647),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_57),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_692),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_861),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_683),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_444),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_963),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_711),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_562),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_458),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_227),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_322),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_766),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_700),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_891),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1039),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_451),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_523),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_194),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1008),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_999),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1035),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_2),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_915),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_705),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_689),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_389),
.Y(n_1312)
);

CKINVDCx16_ASAP7_75t_R g1313 ( 
.A(n_604),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_918),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_734),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_483),
.Y(n_1316)
);

BUFx10_ASAP7_75t_L g1317 ( 
.A(n_486),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_226),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_603),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_607),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_950),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_807),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_562),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_894),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_659),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_267),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_606),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_892),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_712),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_87),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1053),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_697),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_427),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_468),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_810),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_661),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_898),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_115),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_675),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_875),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_604),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_210),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_687),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_728),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_707),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_854),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_408),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_618),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_244),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_267),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_158),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_679),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_651),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_156),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_435),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_473),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_939),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_143),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_538),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_673),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_658),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_998),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1037),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_509),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1026),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_509),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_442),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_269),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_679),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_68),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_208),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_96),
.Y(n_1372)
);

BUFx10_ASAP7_75t_L g1373 ( 
.A(n_750),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_397),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_822),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1033),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_382),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_174),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_304),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_293),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_598),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_137),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_355),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_706),
.Y(n_1384)
);

BUFx8_ASAP7_75t_SL g1385 ( 
.A(n_402),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1002),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_674),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1003),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_971),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_53),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_3),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_209),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_843),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_500),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_117),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_147),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_696),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1023),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_714),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_96),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_796),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_577),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_473),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1038),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_450),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_223),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_656),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_811),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_616),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_553),
.Y(n_1410)
);

CKINVDCx16_ASAP7_75t_R g1411 ( 
.A(n_759),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_252),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_718),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_770),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_906),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_573),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_80),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1028),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_801),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_693),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_119),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_429),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1042),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_685),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_101),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_471),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_47),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_713),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1016),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_751),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_717),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_448),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_958),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1021),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_581),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_869),
.Y(n_1436)
);

BUFx10_ASAP7_75t_L g1437 ( 
.A(n_89),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_123),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_399),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_802),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_309),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_210),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_669),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_13),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_368),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_590),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_809),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_201),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_356),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_678),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_499),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_407),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_671),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1047),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_89),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1044),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_325),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_18),
.Y(n_1458)
);

BUFx2_ASAP7_75t_SL g1459 ( 
.A(n_499),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_709),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_204),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_586),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_594),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_805),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_114),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_708),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_699),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_350),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_153),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_10),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1045),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_397),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_867),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_373),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_442),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_339),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_717),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_907),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1043),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_851),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_714),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_533),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_85),
.Y(n_1483)
);

BUFx5_ASAP7_75t_L g1484 ( 
.A(n_273),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_237),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_670),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_704),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1018),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_762),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_209),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_413),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_897),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_127),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_22),
.Y(n_1494)
);

BUFx10_ASAP7_75t_L g1495 ( 
.A(n_40),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_970),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_147),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_235),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_923),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_698),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_78),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_957),
.Y(n_1502)
);

CKINVDCx14_ASAP7_75t_R g1503 ( 
.A(n_103),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_12),
.Y(n_1504)
);

INVxp67_ASAP7_75t_L g1505 ( 
.A(n_345),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_453),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_680),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_359),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_218),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_104),
.Y(n_1510)
);

CKINVDCx14_ASAP7_75t_R g1511 ( 
.A(n_196),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_569),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_783),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_702),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_527),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_739),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_388),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_476),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_12),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_705),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_703),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_778),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_101),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_106),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_73),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_383),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_229),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_586),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_687),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_116),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_183),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1054),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_398),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_701),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_579),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_746),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_931),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_372),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_93),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_81),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_302),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_877),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1046),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_198),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1029),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_361),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_501),
.Y(n_1547)
);

CKINVDCx16_ASAP7_75t_R g1548 ( 
.A(n_1034),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_733),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_225),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_366),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_295),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_948),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_492),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_385),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_460),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_342),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1013),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1051),
.Y(n_1559)
);

BUFx5_ASAP7_75t_L g1560 ( 
.A(n_597),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_187),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_259),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_591),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_954),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1059),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1484),
.Y(n_1566)
);

INVxp33_ASAP7_75t_SL g1567 ( 
.A(n_1461),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1250),
.Y(n_1568)
);

INVxp67_ASAP7_75t_SL g1569 ( 
.A(n_1107),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1484),
.Y(n_1570)
);

CKINVDCx14_ASAP7_75t_R g1571 ( 
.A(n_1125),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1111),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1484),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1484),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1385),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1118),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1484),
.Y(n_1577)
);

INVxp67_ASAP7_75t_SL g1578 ( 
.A(n_1068),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1560),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1560),
.Y(n_1580)
);

INVxp67_ASAP7_75t_SL g1581 ( 
.A(n_1074),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1127),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1060),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1067),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1272),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1222),
.B(n_0),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1560),
.Y(n_1587)
);

CKINVDCx20_ASAP7_75t_R g1588 ( 
.A(n_1328),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1072),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_1346),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1075),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1433),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1062),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1560),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1560),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1062),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1081),
.Y(n_1597)
);

NOR2xp67_ASAP7_75t_L g1598 ( 
.A(n_1356),
.B(n_1),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1062),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1122),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1488),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1122),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1122),
.Y(n_1603)
);

CKINVDCx16_ASAP7_75t_R g1604 ( 
.A(n_1063),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1089),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1133),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1104),
.Y(n_1607)
);

CKINVDCx14_ASAP7_75t_R g1608 ( 
.A(n_1503),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1133),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_1502),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1109),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1271),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1133),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1123),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1141),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1141),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1141),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_1283),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1177),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1177),
.Y(n_1620)
);

CKINVDCx16_ASAP7_75t_R g1621 ( 
.A(n_1132),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1177),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1249),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_R g1624 ( 
.A(n_1238),
.B(n_1048),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1249),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1130),
.Y(n_1626)
);

INVxp67_ASAP7_75t_SL g1627 ( 
.A(n_1309),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1511),
.B(n_4),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1249),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_1411),
.Y(n_1630)
);

CKINVDCx16_ASAP7_75t_R g1631 ( 
.A(n_1241),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1299),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_1548),
.Y(n_1633)
);

INVxp33_ASAP7_75t_L g1634 ( 
.A(n_1518),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1098),
.B(n_3),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1513),
.B(n_5),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1299),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1135),
.Y(n_1638)
);

CKINVDCx20_ASAP7_75t_R g1639 ( 
.A(n_1138),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1129),
.B(n_4),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1596),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1599),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1593),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1600),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1602),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1603),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1567),
.A2(n_1313),
.B1(n_1137),
.B2(n_1284),
.Y(n_1647)
);

AND3x1_ASAP7_75t_L g1648 ( 
.A(n_1636),
.B(n_1227),
.C(n_1169),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1606),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1593),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1583),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1639),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1609),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1613),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1615),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1616),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1617),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1619),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1620),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1622),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1623),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1625),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1629),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1632),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1637),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1584),
.B(n_1331),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1566),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1570),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1578),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1589),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1573),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1574),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1571),
.B(n_1064),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1577),
.A2(n_1580),
.B(n_1579),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1591),
.B(n_1436),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1597),
.B(n_1357),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1594),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1605),
.B(n_1440),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1581),
.B(n_1537),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1595),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1587),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1612),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1640),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1627),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1569),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1604),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1598),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1608),
.B(n_1092),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1635),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1607),
.B(n_1276),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1611),
.B(n_1614),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1586),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1628),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1621),
.B(n_1198),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1626),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1638),
.B(n_1300),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1624),
.B(n_1365),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1634),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1568),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1631),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1618),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1630),
.B(n_1263),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1633),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1671),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1671),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1649),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1667),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1668),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1672),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1697),
.B(n_1281),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1698),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1649),
.Y(n_1712)
);

NAND2x1p5_ASAP7_75t_L g1713 ( 
.A(n_1699),
.B(n_1322),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1657),
.Y(n_1714)
);

INVx4_ASAP7_75t_L g1715 ( 
.A(n_1692),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1689),
.B(n_1572),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1657),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1679),
.B(n_1213),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1690),
.B(n_1575),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1696),
.B(n_1565),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1643),
.B(n_1342),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_L g1722 ( 
.A(n_1685),
.B(n_1061),
.C(n_1058),
.Y(n_1722)
);

OAI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1647),
.A2(n_1207),
.B1(n_1291),
.B2(n_1162),
.Y(n_1723)
);

OR2x2_ASAP7_75t_SL g1724 ( 
.A(n_1693),
.B(n_1077),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1665),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1665),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1650),
.B(n_1319),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_SL g1728 ( 
.A(n_1692),
.B(n_1076),
.Y(n_1728)
);

BUFx10_ASAP7_75t_L g1729 ( 
.A(n_1700),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1677),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1693),
.B(n_1198),
.Y(n_1731)
);

OAI21xp33_ASAP7_75t_L g1732 ( 
.A1(n_1687),
.A2(n_1435),
.B(n_1428),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1641),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1680),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1642),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1664),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1686),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1681),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1656),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1644),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1683),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1651),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1682),
.B(n_1504),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1673),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1669),
.A2(n_1576),
.B1(n_1585),
.B2(n_1582),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1645),
.Y(n_1746)
);

INVx4_ASAP7_75t_L g1747 ( 
.A(n_1670),
.Y(n_1747)
);

INVxp33_ASAP7_75t_L g1748 ( 
.A(n_1688),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1683),
.B(n_1363),
.Y(n_1749)
);

NAND2xp33_ASAP7_75t_L g1750 ( 
.A(n_1666),
.B(n_1434),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1684),
.B(n_1414),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1658),
.Y(n_1752)
);

BUFx6f_ASAP7_75t_L g1753 ( 
.A(n_1674),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1646),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1676),
.B(n_1492),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1702),
.B(n_1373),
.Y(n_1756)
);

AO22x2_ASAP7_75t_L g1757 ( 
.A1(n_1694),
.A2(n_1459),
.B1(n_1413),
.B2(n_1371),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1653),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1678),
.B(n_1140),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1675),
.B(n_1105),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1695),
.B(n_1373),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1654),
.B(n_1655),
.Y(n_1762)
);

AND3x4_ASAP7_75t_L g1763 ( 
.A(n_1652),
.B(n_1405),
.C(n_1403),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1691),
.B(n_1149),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1648),
.B(n_1455),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1659),
.B(n_1663),
.Y(n_1766)
);

NAND2xp33_ASAP7_75t_L g1767 ( 
.A(n_1660),
.B(n_1434),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_1661),
.Y(n_1768)
);

OAI21xp33_ASAP7_75t_L g1769 ( 
.A1(n_1662),
.A2(n_1501),
.B(n_1420),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1701),
.B(n_1588),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1703),
.B(n_1590),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1671),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1698),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1671),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1671),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1679),
.B(n_1466),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1671),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1671),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1693),
.B(n_1157),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1739),
.Y(n_1780)
);

OR2x6_ASAP7_75t_SL g1781 ( 
.A(n_1716),
.B(n_1065),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1710),
.B(n_1066),
.Y(n_1782)
);

AO22x2_ASAP7_75t_L g1783 ( 
.A1(n_1763),
.A2(n_1547),
.B1(n_1483),
.B2(n_1079),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1755),
.B(n_1080),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1752),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1762),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1728),
.Y(n_1787)
);

BUFx8_ASAP7_75t_L g1788 ( 
.A(n_1737),
.Y(n_1788)
);

AO22x2_ASAP7_75t_L g1789 ( 
.A1(n_1756),
.A2(n_1085),
.B1(n_1091),
.B2(n_1071),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1733),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_1749),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1735),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1742),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1740),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1715),
.B(n_1592),
.Y(n_1795)
);

NAND2x1p5_ASAP7_75t_L g1796 ( 
.A(n_1741),
.B(n_1083),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1707),
.Y(n_1797)
);

INVx3_ASAP7_75t_L g1798 ( 
.A(n_1706),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1708),
.Y(n_1799)
);

INVx2_ASAP7_75t_SL g1800 ( 
.A(n_1718),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1709),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1730),
.Y(n_1802)
);

AO22x2_ASAP7_75t_L g1803 ( 
.A1(n_1765),
.A2(n_1095),
.B1(n_1100),
.B2(n_1094),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1760),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1759),
.B(n_1086),
.Y(n_1805)
);

OR2x6_ASAP7_75t_L g1806 ( 
.A(n_1747),
.B(n_1372),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1720),
.A2(n_1610),
.B1(n_1601),
.B2(n_1161),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_1744),
.Y(n_1808)
);

AO22x2_ASAP7_75t_L g1809 ( 
.A1(n_1731),
.A2(n_1102),
.B1(n_1115),
.B2(n_1101),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1711),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1748),
.B(n_1105),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1753),
.A2(n_1479),
.B1(n_1558),
.B2(n_1454),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1734),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1764),
.B(n_1099),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1746),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1738),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1719),
.A2(n_1171),
.B1(n_1174),
.B2(n_1160),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1766),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1754),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1773),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1745),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1722),
.A2(n_1188),
.B1(n_1189),
.B2(n_1180),
.Y(n_1822)
);

AO22x2_ASAP7_75t_L g1823 ( 
.A1(n_1723),
.A2(n_1327),
.B1(n_1378),
.B2(n_1172),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1743),
.B(n_1139),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1736),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1758),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1714),
.B(n_1705),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1704),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1753),
.B(n_1120),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1721),
.Y(n_1830)
);

AOI22x1_ASAP7_75t_L g1831 ( 
.A1(n_1757),
.A2(n_1128),
.B1(n_1147),
.B2(n_1124),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1758),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1772),
.Y(n_1833)
);

NAND2xp33_ASAP7_75t_L g1834 ( 
.A(n_1751),
.B(n_1191),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1774),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1727),
.B(n_1465),
.Y(n_1836)
);

AO22x2_ASAP7_75t_L g1837 ( 
.A1(n_1761),
.A2(n_1143),
.B1(n_1144),
.B2(n_1121),
.Y(n_1837)
);

BUFx3_ASAP7_75t_L g1838 ( 
.A(n_1778),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1768),
.Y(n_1839)
);

AO22x2_ASAP7_75t_L g1840 ( 
.A1(n_1776),
.A2(n_1158),
.B1(n_1194),
.B2(n_1148),
.Y(n_1840)
);

NAND2x1p5_ASAP7_75t_L g1841 ( 
.A(n_1706),
.B(n_1153),
.Y(n_1841)
);

NAND2xp33_ASAP7_75t_L g1842 ( 
.A(n_1778),
.B(n_1775),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1777),
.Y(n_1843)
);

AO22x2_ASAP7_75t_L g1844 ( 
.A1(n_1779),
.A2(n_1264),
.B1(n_1286),
.B2(n_1176),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1768),
.B(n_1190),
.Y(n_1845)
);

OR2x6_ASAP7_75t_L g1846 ( 
.A(n_1713),
.B(n_1505),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1770),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1769),
.A2(n_1215),
.B1(n_1221),
.B2(n_1199),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1732),
.A2(n_1216),
.B1(n_1239),
.B2(n_1200),
.Y(n_1849)
);

AND2x6_ASAP7_75t_L g1850 ( 
.A(n_1771),
.B(n_1248),
.Y(n_1850)
);

BUFx8_ASAP7_75t_L g1851 ( 
.A(n_1725),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1724),
.Y(n_1852)
);

AO22x2_ASAP7_75t_L g1853 ( 
.A1(n_1712),
.A2(n_1225),
.B1(n_1329),
.B2(n_1178),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1717),
.B(n_1253),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1725),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1726),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1726),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1750),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1767),
.B(n_1259),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1729),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1739),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1741),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1747),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1715),
.B(n_1152),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1739),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1739),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1710),
.B(n_1335),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1710),
.B(n_1337),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1762),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1715),
.B(n_1155),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1739),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1739),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1720),
.A2(n_1236),
.B1(n_1243),
.B2(n_1224),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1762),
.Y(n_1874)
);

AO22x2_ASAP7_75t_L g1875 ( 
.A1(n_1763),
.A2(n_1218),
.B1(n_1308),
.B2(n_1182),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1715),
.B(n_1163),
.Y(n_1876)
);

OAI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1769),
.A2(n_1167),
.B1(n_1196),
.B2(n_1192),
.C(n_1185),
.Y(n_1877)
);

NAND2x1p5_ASAP7_75t_L g1878 ( 
.A(n_1715),
.B(n_1362),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1739),
.Y(n_1879)
);

AOI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1720),
.A2(n_1246),
.B1(n_1266),
.B2(n_1244),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1710),
.B(n_1376),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1710),
.B(n_1389),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1710),
.B(n_1408),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1739),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1715),
.B(n_1197),
.Y(n_1885)
);

AO22x2_ASAP7_75t_L g1886 ( 
.A1(n_1763),
.A2(n_1303),
.B1(n_1452),
.B2(n_1294),
.Y(n_1886)
);

AO22x2_ASAP7_75t_L g1887 ( 
.A1(n_1763),
.A2(n_1374),
.B1(n_1394),
.B2(n_1360),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1739),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1739),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1739),
.Y(n_1890)
);

OAI22x1_ASAP7_75t_SL g1891 ( 
.A1(n_1747),
.A2(n_1097),
.B1(n_1164),
.B2(n_1087),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1715),
.B(n_1278),
.Y(n_1892)
);

AO22x2_ASAP7_75t_L g1893 ( 
.A1(n_1763),
.A2(n_1252),
.B1(n_1334),
.B2(n_1209),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1715),
.B(n_1553),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1739),
.Y(n_1895)
);

INVxp67_ASAP7_75t_L g1896 ( 
.A(n_1749),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1749),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1739),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1762),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1715),
.B(n_1242),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1755),
.B(n_1069),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1739),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1715),
.B(n_1559),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1762),
.Y(n_1904)
);

AO22x2_ASAP7_75t_L g1905 ( 
.A1(n_1763),
.A2(n_1421),
.B1(n_1494),
.B2(n_1351),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1710),
.B(n_1429),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1739),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1710),
.B(n_1464),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1778),
.Y(n_1909)
);

BUFx8_ASAP7_75t_L g1910 ( 
.A(n_1737),
.Y(n_1910)
);

AO22x2_ASAP7_75t_L g1911 ( 
.A1(n_1763),
.A2(n_1390),
.B1(n_1514),
.B2(n_1380),
.Y(n_1911)
);

BUFx3_ASAP7_75t_L g1912 ( 
.A(n_1741),
.Y(n_1912)
);

AO22x2_ASAP7_75t_L g1913 ( 
.A1(n_1763),
.A2(n_1458),
.B1(n_1438),
.B2(n_1265),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1739),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1728),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1710),
.B(n_1478),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1741),
.B(n_1139),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1739),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_SL g1919 ( 
.A(n_1765),
.Y(n_1919)
);

AO22x2_ASAP7_75t_L g1920 ( 
.A1(n_1763),
.A2(n_1354),
.B1(n_1475),
.B2(n_1297),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1739),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1791),
.B(n_1289),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1896),
.B(n_1897),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1818),
.B(n_1292),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1804),
.B(n_1847),
.Y(n_1925)
);

NAND2xp33_ASAP7_75t_SL g1926 ( 
.A(n_1863),
.B(n_1229),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1901),
.B(n_1298),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1869),
.B(n_1301),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1874),
.B(n_1305),
.Y(n_1929)
);

NAND2xp33_ASAP7_75t_SL g1930 ( 
.A(n_1787),
.B(n_1232),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1782),
.B(n_1867),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1899),
.B(n_1306),
.Y(n_1932)
);

NAND2xp33_ASAP7_75t_SL g1933 ( 
.A(n_1915),
.B(n_1256),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1904),
.B(n_1307),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1810),
.B(n_1314),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1826),
.B(n_1260),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1820),
.B(n_1315),
.Y(n_1937)
);

NAND2xp33_ASAP7_75t_SL g1938 ( 
.A(n_1852),
.B(n_1270),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1868),
.B(n_1522),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1786),
.B(n_1321),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1780),
.B(n_1785),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1797),
.B(n_1324),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1799),
.B(n_1340),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1824),
.B(n_1154),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1801),
.B(n_1344),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1802),
.B(n_1375),
.Y(n_1946)
);

NAND2xp33_ASAP7_75t_SL g1947 ( 
.A(n_1919),
.B(n_1336),
.Y(n_1947)
);

NAND2xp33_ASAP7_75t_SL g1948 ( 
.A(n_1909),
.B(n_1345),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1813),
.B(n_1386),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1861),
.B(n_1388),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1865),
.B(n_1866),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1871),
.B(n_1393),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1872),
.B(n_1398),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1879),
.B(n_1401),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1884),
.B(n_1404),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1888),
.B(n_1415),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1889),
.B(n_1418),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1890),
.B(n_1419),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1895),
.B(n_1423),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1881),
.B(n_1536),
.Y(n_1960)
);

NAND2xp33_ASAP7_75t_SL g1961 ( 
.A(n_1909),
.B(n_1352),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1898),
.B(n_1430),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1902),
.B(n_1447),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1907),
.B(n_1456),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1836),
.B(n_1154),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1882),
.B(n_1542),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1883),
.B(n_1549),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1906),
.B(n_1471),
.Y(n_1968)
);

NAND2xp33_ASAP7_75t_SL g1969 ( 
.A(n_1821),
.B(n_1364),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1914),
.B(n_1473),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1918),
.B(n_1480),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1921),
.B(n_1489),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1808),
.B(n_1496),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1784),
.B(n_1499),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1816),
.B(n_1516),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1908),
.B(n_1532),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1916),
.B(n_1543),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1811),
.B(n_1230),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1873),
.B(n_1545),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1880),
.B(n_1814),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1819),
.B(n_1564),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1793),
.B(n_1434),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1805),
.B(n_1299),
.Y(n_1983)
);

NAND2xp33_ASAP7_75t_SL g1984 ( 
.A(n_1860),
.B(n_1830),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1829),
.B(n_1406),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1790),
.B(n_1406),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1807),
.B(n_1400),
.Y(n_1987)
);

NAND2xp33_ASAP7_75t_SL g1988 ( 
.A(n_1800),
.B(n_1409),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1817),
.B(n_1422),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1822),
.B(n_1825),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1917),
.B(n_1432),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1832),
.B(n_1441),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1839),
.B(n_1460),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1792),
.B(n_1406),
.Y(n_1994)
);

NAND2xp33_ASAP7_75t_SL g1995 ( 
.A(n_1849),
.B(n_1070),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1846),
.B(n_1230),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1794),
.B(n_1073),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1846),
.B(n_1233),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1815),
.B(n_1078),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1795),
.B(n_1082),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1864),
.B(n_1088),
.Y(n_2001)
);

NAND2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1855),
.B(n_1090),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1827),
.B(n_1268),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1870),
.B(n_1096),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1850),
.B(n_1103),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_SL g2006 ( 
.A(n_1876),
.B(n_1106),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1885),
.B(n_1108),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1900),
.B(n_1110),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1850),
.B(n_1112),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1850),
.B(n_1113),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1848),
.B(n_1114),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1845),
.B(n_1116),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1831),
.B(n_1117),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1858),
.B(n_1119),
.Y(n_2014)
);

NAND2xp33_ASAP7_75t_SL g2015 ( 
.A(n_1856),
.B(n_1126),
.Y(n_2015)
);

NAND2xp33_ASAP7_75t_SL g2016 ( 
.A(n_1857),
.B(n_1131),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_SL g2017 ( 
.A(n_1798),
.B(n_1134),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1828),
.B(n_1136),
.Y(n_2018)
);

NAND2xp33_ASAP7_75t_SL g2019 ( 
.A(n_1833),
.B(n_1142),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1812),
.B(n_1145),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1835),
.B(n_1843),
.Y(n_2021)
);

NAND2xp33_ASAP7_75t_SL g2022 ( 
.A(n_1892),
.B(n_1146),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1854),
.B(n_1150),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1862),
.B(n_1279),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1878),
.B(n_1151),
.Y(n_2025)
);

NAND2xp33_ASAP7_75t_SL g2026 ( 
.A(n_1894),
.B(n_1156),
.Y(n_2026)
);

NAND2xp33_ASAP7_75t_SL g2027 ( 
.A(n_1903),
.B(n_1159),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1912),
.B(n_1165),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1838),
.B(n_1166),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1796),
.B(n_1168),
.Y(n_2030)
);

NAND2xp33_ASAP7_75t_SL g2031 ( 
.A(n_1789),
.B(n_1170),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1841),
.B(n_1173),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1806),
.B(n_1175),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1834),
.B(n_1179),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1788),
.B(n_1183),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1806),
.B(n_1233),
.Y(n_2036)
);

NAND2xp33_ASAP7_75t_SL g2037 ( 
.A(n_1859),
.B(n_1184),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1844),
.B(n_1186),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1853),
.B(n_1317),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1910),
.B(n_1193),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1851),
.B(n_1195),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1809),
.B(n_1201),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1837),
.B(n_1202),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1823),
.B(n_1203),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1781),
.B(n_1204),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1877),
.B(n_1803),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1875),
.B(n_1205),
.Y(n_2047)
);

NAND2xp33_ASAP7_75t_SL g2048 ( 
.A(n_1886),
.B(n_1206),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1887),
.B(n_1208),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1893),
.B(n_1210),
.Y(n_2050)
);

NAND2xp33_ASAP7_75t_SL g2051 ( 
.A(n_1905),
.B(n_1211),
.Y(n_2051)
);

XNOR2x2_ASAP7_75t_L g2052 ( 
.A(n_1911),
.B(n_1312),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1913),
.B(n_1212),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1920),
.B(n_1214),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1783),
.B(n_1217),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1840),
.B(n_1219),
.Y(n_2056)
);

NAND2xp33_ASAP7_75t_SL g2057 ( 
.A(n_1842),
.B(n_1220),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1891),
.B(n_1223),
.Y(n_2058)
);

NAND2xp33_ASAP7_75t_SL g2059 ( 
.A(n_1863),
.B(n_1226),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1818),
.B(n_1228),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1824),
.B(n_1317),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1824),
.B(n_1437),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1791),
.B(n_1234),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1791),
.B(n_1237),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1818),
.B(n_1240),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1818),
.B(n_1245),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_1791),
.B(n_1247),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1791),
.B(n_1251),
.Y(n_2068)
);

NAND2xp33_ASAP7_75t_SL g2069 ( 
.A(n_1863),
.B(n_1254),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_SL g2070 ( 
.A(n_1791),
.B(n_1255),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1791),
.B(n_1257),
.Y(n_2071)
);

NAND2xp33_ASAP7_75t_SL g2072 ( 
.A(n_1863),
.B(n_1258),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1791),
.B(n_1261),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1791),
.B(n_1262),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1791),
.B(n_1267),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1791),
.B(n_1269),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1791),
.B(n_1273),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1791),
.B(n_1274),
.Y(n_2078)
);

NAND2xp33_ASAP7_75t_SL g2079 ( 
.A(n_1863),
.B(n_1275),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1791),
.B(n_1277),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1791),
.B(n_1280),
.Y(n_2081)
);

NAND2xp33_ASAP7_75t_SL g2082 ( 
.A(n_1863),
.B(n_1282),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1791),
.B(n_1285),
.Y(n_2083)
);

NAND2xp33_ASAP7_75t_SL g2084 ( 
.A(n_1863),
.B(n_1287),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_SL g2085 ( 
.A(n_1791),
.B(n_1288),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_1824),
.B(n_1437),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1791),
.B(n_1290),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1818),
.B(n_1293),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1818),
.B(n_1295),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1791),
.B(n_1296),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1791),
.B(n_1304),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1791),
.B(n_1310),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1818),
.B(n_1311),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1791),
.B(n_1316),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1824),
.B(n_1495),
.Y(n_2095)
);

NAND2xp33_ASAP7_75t_SL g2096 ( 
.A(n_1863),
.B(n_1318),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1791),
.B(n_1320),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1791),
.B(n_1325),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1791),
.B(n_1326),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1818),
.B(n_1330),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1791),
.B(n_1332),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1791),
.B(n_1333),
.Y(n_2102)
);

NAND2xp33_ASAP7_75t_SL g2103 ( 
.A(n_1863),
.B(n_1338),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1791),
.B(n_1341),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1818),
.B(n_1343),
.Y(n_2105)
);

NAND2xp33_ASAP7_75t_SL g2106 ( 
.A(n_1863),
.B(n_1347),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1791),
.B(n_1348),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1826),
.B(n_1323),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1791),
.B(n_1350),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1791),
.B(n_1358),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1791),
.B(n_1366),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_1791),
.B(n_1367),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1791),
.B(n_1368),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1791),
.B(n_1369),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1791),
.B(n_1370),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1818),
.B(n_1377),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1791),
.B(n_1379),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1791),
.B(n_1381),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_1791),
.B(n_1382),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1791),
.B(n_1383),
.Y(n_2120)
);

NAND2xp33_ASAP7_75t_SL g2121 ( 
.A(n_1863),
.B(n_1384),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1791),
.B(n_1387),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1818),
.B(n_1392),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1931),
.B(n_1395),
.Y(n_2124)
);

AOI21x1_ASAP7_75t_L g2125 ( 
.A1(n_1985),
.A2(n_1349),
.B(n_1339),
.Y(n_2125)
);

OAI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_1980),
.A2(n_1402),
.B1(n_1407),
.B2(n_1399),
.Y(n_2126)
);

OAI21xp5_ASAP7_75t_SL g2127 ( 
.A1(n_1987),
.A2(n_1551),
.B(n_1550),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2060),
.B(n_1410),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2065),
.B(n_1412),
.Y(n_2129)
);

OAI22x1_ASAP7_75t_L g2130 ( 
.A1(n_1989),
.A2(n_1424),
.B1(n_1425),
.B2(n_1417),
.Y(n_2130)
);

A2O1A1Ixp33_ASAP7_75t_L g2131 ( 
.A1(n_2046),
.A2(n_1359),
.B(n_1361),
.C(n_1353),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_SL g2132 ( 
.A1(n_2033),
.A2(n_1482),
.B1(n_1497),
.B2(n_1449),
.Y(n_2132)
);

AOI21xp5_ASAP7_75t_L g2133 ( 
.A1(n_1990),
.A2(n_1397),
.B(n_1396),
.Y(n_2133)
);

OAI21x1_ASAP7_75t_L g2134 ( 
.A1(n_1986),
.A2(n_1431),
.B(n_1416),
.Y(n_2134)
);

O2A1O1Ixp5_ASAP7_75t_L g2135 ( 
.A1(n_2013),
.A2(n_1443),
.B(n_1446),
.C(n_1439),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_1941),
.A2(n_1470),
.B(n_1468),
.Y(n_2136)
);

OAI21xp5_ASAP7_75t_SL g2137 ( 
.A1(n_1991),
.A2(n_1508),
.B(n_1490),
.Y(n_2137)
);

AOI21xp5_ASAP7_75t_SL g2138 ( 
.A1(n_2014),
.A2(n_721),
.B(n_720),
.Y(n_2138)
);

O2A1O1Ixp33_ASAP7_75t_L g2139 ( 
.A1(n_1925),
.A2(n_1510),
.B(n_1519),
.C(n_1509),
.Y(n_2139)
);

AND2x4_ASAP7_75t_L g2140 ( 
.A(n_2003),
.B(n_1528),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2066),
.B(n_1426),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1936),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1936),
.Y(n_2143)
);

OAI21x1_ASAP7_75t_L g2144 ( 
.A1(n_1951),
.A2(n_1539),
.B(n_1535),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_2024),
.Y(n_2145)
);

CKINVDCx11_ASAP7_75t_R g2146 ( 
.A(n_2024),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_1924),
.A2(n_1546),
.B(n_1540),
.Y(n_2147)
);

AO21x2_ASAP7_75t_L g2148 ( 
.A1(n_1927),
.A2(n_1976),
.B(n_1974),
.Y(n_2148)
);

AOI21x1_ASAP7_75t_L g2149 ( 
.A1(n_1983),
.A2(n_1552),
.B(n_1093),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2108),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2108),
.Y(n_2151)
);

BUFx12f_ASAP7_75t_L g2152 ( 
.A(n_2003),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2088),
.B(n_1427),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2021),
.Y(n_2154)
);

AOI21xp5_ASAP7_75t_L g2155 ( 
.A1(n_1928),
.A2(n_1181),
.B(n_1084),
.Y(n_2155)
);

OAI21x1_ASAP7_75t_L g2156 ( 
.A1(n_1929),
.A2(n_1231),
.B(n_1187),
.Y(n_2156)
);

AO21x2_ASAP7_75t_L g2157 ( 
.A1(n_1977),
.A2(n_1302),
.B(n_1235),
.Y(n_2157)
);

INVx1_ASAP7_75t_SL g2158 ( 
.A(n_1948),
.Y(n_2158)
);

AO21x1_ASAP7_75t_L g2159 ( 
.A1(n_2031),
.A2(n_1391),
.B(n_1355),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1944),
.B(n_1495),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2089),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2093),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1947),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2100),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2105),
.B(n_1442),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2116),
.B(n_1444),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2123),
.B(n_1445),
.Y(n_2167)
);

NOR3xp33_ASAP7_75t_L g2168 ( 
.A(n_1926),
.B(n_1450),
.C(n_1448),
.Y(n_2168)
);

AOI31xp67_ASAP7_75t_L g2169 ( 
.A1(n_1939),
.A2(n_1544),
.A3(n_1555),
.B(n_1463),
.Y(n_2169)
);

OAI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_2011),
.A2(n_1562),
.B(n_1453),
.Y(n_2170)
);

AOI21xp5_ASAP7_75t_L g2171 ( 
.A1(n_1932),
.A2(n_1934),
.B(n_1940),
.Y(n_2171)
);

INVx4_ASAP7_75t_L g2172 ( 
.A(n_1996),
.Y(n_2172)
);

AOI21x1_ASAP7_75t_L g2173 ( 
.A1(n_1960),
.A2(n_724),
.B(n_722),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_1968),
.A2(n_726),
.B(n_725),
.Y(n_2174)
);

INVx1_ASAP7_75t_SL g2175 ( 
.A(n_1961),
.Y(n_2175)
);

AO21x2_ASAP7_75t_L g2176 ( 
.A1(n_1966),
.A2(n_729),
.B(n_727),
.Y(n_2176)
);

OAI21x1_ASAP7_75t_L g2177 ( 
.A1(n_1967),
.A2(n_731),
.B(n_730),
.Y(n_2177)
);

O2A1O1Ixp5_ASAP7_75t_L g2178 ( 
.A1(n_1979),
.A2(n_736),
.B(n_737),
.C(n_735),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_1923),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2061),
.B(n_1451),
.Y(n_2180)
);

OAI21x1_ASAP7_75t_L g2181 ( 
.A1(n_1981),
.A2(n_740),
.B(n_738),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_1969),
.B(n_1930),
.Y(n_2182)
);

AOI21xp5_ASAP7_75t_L g2183 ( 
.A1(n_1942),
.A2(n_743),
.B(n_741),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2062),
.B(n_2086),
.Y(n_2184)
);

AO32x2_ASAP7_75t_L g2185 ( 
.A1(n_2052),
.A2(n_7),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1978),
.B(n_1457),
.Y(n_2186)
);

OAI21x1_ASAP7_75t_L g2187 ( 
.A1(n_1943),
.A2(n_745),
.B(n_744),
.Y(n_2187)
);

BUFx6f_ASAP7_75t_L g2188 ( 
.A(n_1998),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2095),
.B(n_1462),
.Y(n_2189)
);

OAI21x1_ASAP7_75t_L g2190 ( 
.A1(n_1945),
.A2(n_748),
.B(n_747),
.Y(n_2190)
);

INVx4_ASAP7_75t_SL g2191 ( 
.A(n_2036),
.Y(n_2191)
);

OA21x2_ASAP7_75t_L g2192 ( 
.A1(n_1997),
.A2(n_1469),
.B(n_1467),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1965),
.B(n_1922),
.Y(n_2193)
);

A2O1A1Ixp33_ASAP7_75t_L g2194 ( 
.A1(n_1995),
.A2(n_2005),
.B(n_2010),
.C(n_2009),
.Y(n_2194)
);

OAI21x1_ASAP7_75t_L g2195 ( 
.A1(n_1946),
.A2(n_752),
.B(n_749),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_1933),
.B(n_1472),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2063),
.B(n_1474),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_L g2198 ( 
.A1(n_1949),
.A2(n_1952),
.B(n_1950),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2064),
.B(n_2067),
.Y(n_2199)
);

INVx1_ASAP7_75t_SL g2200 ( 
.A(n_2002),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_2034),
.B(n_1476),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_2059),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1994),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1999),
.Y(n_2204)
);

BUFx4_ASAP7_75t_SL g2205 ( 
.A(n_1938),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2020),
.Y(n_2206)
);

AO31x2_ASAP7_75t_L g2207 ( 
.A1(n_2038),
.A2(n_755),
.A3(n_756),
.B(n_754),
.Y(n_2207)
);

OAI21xp5_ASAP7_75t_L g2208 ( 
.A1(n_1953),
.A2(n_1481),
.B(n_1477),
.Y(n_2208)
);

AOI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_1954),
.A2(n_758),
.B(n_757),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2018),
.Y(n_2210)
);

OAI21x1_ASAP7_75t_L g2211 ( 
.A1(n_1955),
.A2(n_761),
.B(n_760),
.Y(n_2211)
);

OAI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_1956),
.A2(n_1486),
.B(n_1485),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_1992),
.B(n_1487),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2044),
.Y(n_2214)
);

O2A1O1Ixp5_ASAP7_75t_L g2215 ( 
.A1(n_2000),
.A2(n_764),
.B(n_765),
.C(n_763),
.Y(n_2215)
);

NOR2xp67_ASAP7_75t_L g2216 ( 
.A(n_2068),
.B(n_767),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1957),
.Y(n_2217)
);

OAI21x1_ASAP7_75t_SL g2218 ( 
.A1(n_2056),
.A2(n_769),
.B(n_768),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1958),
.Y(n_2219)
);

INVx6_ASAP7_75t_L g2220 ( 
.A(n_2039),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2070),
.B(n_2071),
.Y(n_2221)
);

OAI21xp5_ASAP7_75t_L g2222 ( 
.A1(n_1959),
.A2(n_1493),
.B(n_1491),
.Y(n_2222)
);

AOI21xp5_ASAP7_75t_L g2223 ( 
.A1(n_1962),
.A2(n_773),
.B(n_771),
.Y(n_2223)
);

OAI21x1_ASAP7_75t_L g2224 ( 
.A1(n_1963),
.A2(n_775),
.B(n_774),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1964),
.Y(n_2225)
);

OAI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_1970),
.A2(n_1500),
.B(n_1498),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1971),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_1988),
.B(n_1506),
.Y(n_2228)
);

AO31x2_ASAP7_75t_L g2229 ( 
.A1(n_2043),
.A2(n_777),
.A3(n_782),
.B(n_776),
.Y(n_2229)
);

NOR3xp33_ASAP7_75t_L g2230 ( 
.A(n_1993),
.B(n_1512),
.C(n_1507),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1972),
.Y(n_2231)
);

OAI21x1_ASAP7_75t_L g2232 ( 
.A1(n_1975),
.A2(n_785),
.B(n_784),
.Y(n_2232)
);

BUFx6f_ASAP7_75t_L g2233 ( 
.A(n_2028),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_1937),
.A2(n_787),
.B(n_786),
.Y(n_2234)
);

AO31x2_ASAP7_75t_L g2235 ( 
.A1(n_2042),
.A2(n_790),
.A3(n_791),
.B(n_788),
.Y(n_2235)
);

BUFx2_ASAP7_75t_L g2236 ( 
.A(n_2017),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2073),
.B(n_1515),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2074),
.B(n_1517),
.Y(n_2238)
);

AOI21xp5_ASAP7_75t_L g2239 ( 
.A1(n_2023),
.A2(n_2012),
.B(n_2075),
.Y(n_2239)
);

HB1xp67_ASAP7_75t_L g2240 ( 
.A(n_2047),
.Y(n_2240)
);

AOI21xp5_ASAP7_75t_L g2241 ( 
.A1(n_2076),
.A2(n_794),
.B(n_793),
.Y(n_2241)
);

OAI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_2077),
.A2(n_1521),
.B1(n_1523),
.B2(n_1520),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1982),
.Y(n_2243)
);

AO32x2_ASAP7_75t_L g2244 ( 
.A1(n_2048),
.A2(n_10),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2078),
.Y(n_2245)
);

OAI21x1_ASAP7_75t_L g2246 ( 
.A1(n_2029),
.A2(n_2025),
.B(n_1973),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2080),
.B(n_1524),
.Y(n_2247)
);

AOI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2081),
.A2(n_1526),
.B1(n_1527),
.B2(n_1525),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2083),
.Y(n_2249)
);

NAND3xp33_ASAP7_75t_L g2250 ( 
.A(n_2069),
.B(n_1530),
.C(n_1529),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_R g2251 ( 
.A(n_2072),
.B(n_1531),
.Y(n_2251)
);

INVxp67_ASAP7_75t_SL g2252 ( 
.A(n_2085),
.Y(n_2252)
);

OAI21x1_ASAP7_75t_L g2253 ( 
.A1(n_2030),
.A2(n_797),
.B(n_795),
.Y(n_2253)
);

AOI21x1_ASAP7_75t_L g2254 ( 
.A1(n_1935),
.A2(n_799),
.B(n_798),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2087),
.Y(n_2255)
);

A2O1A1Ixp33_ASAP7_75t_L g2256 ( 
.A1(n_2022),
.A2(n_1534),
.B(n_1538),
.C(n_1533),
.Y(n_2256)
);

OAI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2090),
.A2(n_1554),
.B1(n_1556),
.B2(n_1541),
.Y(n_2257)
);

INVx4_ASAP7_75t_L g2258 ( 
.A(n_1984),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_2091),
.B(n_1557),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_2079),
.Y(n_2260)
);

AOI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2092),
.A2(n_803),
.B(n_800),
.Y(n_2261)
);

INVxp67_ASAP7_75t_L g2262 ( 
.A(n_2049),
.Y(n_2262)
);

OAI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_2094),
.A2(n_2098),
.B(n_2097),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_2099),
.A2(n_806),
.B(n_804),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_2101),
.B(n_1561),
.Y(n_2265)
);

OAI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_2102),
.A2(n_1563),
.B(n_812),
.Y(n_2266)
);

INVx5_ASAP7_75t_L g2267 ( 
.A(n_2015),
.Y(n_2267)
);

AOI21xp5_ASAP7_75t_L g2268 ( 
.A1(n_2104),
.A2(n_813),
.B(n_808),
.Y(n_2268)
);

AO31x2_ASAP7_75t_L g2269 ( 
.A1(n_2037),
.A2(n_1056),
.A3(n_1057),
.B(n_1055),
.Y(n_2269)
);

AO22x2_ASAP7_75t_L g2270 ( 
.A1(n_2050),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.Y(n_2270)
);

OAI21x1_ASAP7_75t_L g2271 ( 
.A1(n_2032),
.A2(n_817),
.B(n_816),
.Y(n_2271)
);

NOR2xp67_ASAP7_75t_L g2272 ( 
.A(n_2107),
.B(n_818),
.Y(n_2272)
);

OA22x2_ASAP7_75t_L g2273 ( 
.A1(n_2053),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2273)
);

OR2x6_ASAP7_75t_L g2274 ( 
.A(n_2041),
.B(n_15),
.Y(n_2274)
);

AOI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_2109),
.A2(n_820),
.B(n_819),
.Y(n_2275)
);

O2A1O1Ixp33_ASAP7_75t_SL g2276 ( 
.A1(n_2110),
.A2(n_824),
.B(n_825),
.C(n_823),
.Y(n_2276)
);

BUFx6f_ASAP7_75t_L g2277 ( 
.A(n_2035),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2154),
.Y(n_2278)
);

OAI21x1_ASAP7_75t_L g2279 ( 
.A1(n_2156),
.A2(n_2112),
.B(n_2111),
.Y(n_2279)
);

OAI21x1_ASAP7_75t_L g2280 ( 
.A1(n_2136),
.A2(n_2144),
.B(n_2187),
.Y(n_2280)
);

A2O1A1Ixp33_ASAP7_75t_L g2281 ( 
.A1(n_2161),
.A2(n_2027),
.B(n_2026),
.C(n_2019),
.Y(n_2281)
);

OAI21x1_ASAP7_75t_L g2282 ( 
.A1(n_2190),
.A2(n_2211),
.B(n_2195),
.Y(n_2282)
);

OAI222xp33_ASAP7_75t_L g2283 ( 
.A1(n_2273),
.A2(n_2054),
.B1(n_2055),
.B2(n_2058),
.C1(n_2045),
.C2(n_2113),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2143),
.Y(n_2284)
);

OAI21x1_ASAP7_75t_L g2285 ( 
.A1(n_2224),
.A2(n_2115),
.B(n_2114),
.Y(n_2285)
);

OR2x2_ASAP7_75t_L g2286 ( 
.A(n_2124),
.B(n_2117),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2150),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2151),
.Y(n_2288)
);

OA21x2_ASAP7_75t_L g2289 ( 
.A1(n_2194),
.A2(n_2119),
.B(n_2118),
.Y(n_2289)
);

OAI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2162),
.A2(n_2122),
.B(n_2120),
.Y(n_2290)
);

OAI21x1_ASAP7_75t_L g2291 ( 
.A1(n_2232),
.A2(n_2004),
.B(n_2001),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2142),
.Y(n_2292)
);

AOI22xp33_ASAP7_75t_L g2293 ( 
.A1(n_2182),
.A2(n_2051),
.B1(n_2084),
.B2(n_2082),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2164),
.Y(n_2294)
);

OAI21x1_ASAP7_75t_L g2295 ( 
.A1(n_2181),
.A2(n_2007),
.B(n_2006),
.Y(n_2295)
);

AND2x6_ASAP7_75t_L g2296 ( 
.A(n_2206),
.B(n_2008),
.Y(n_2296)
);

A2O1A1Ixp33_ASAP7_75t_L g2297 ( 
.A1(n_2266),
.A2(n_2057),
.B(n_2016),
.C(n_2096),
.Y(n_2297)
);

INVx4_ASAP7_75t_L g2298 ( 
.A(n_2179),
.Y(n_2298)
);

NOR2x1_ASAP7_75t_R g2299 ( 
.A(n_2152),
.B(n_2040),
.Y(n_2299)
);

OAI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2214),
.A2(n_2106),
.B1(n_2121),
.B2(n_2103),
.Y(n_2300)
);

OAI21x1_ASAP7_75t_L g2301 ( 
.A1(n_2177),
.A2(n_830),
.B(n_826),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2203),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_2202),
.Y(n_2303)
);

OAI22xp33_ASAP7_75t_L g2304 ( 
.A1(n_2158),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_2304)
);

AOI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_2259),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2149),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2184),
.B(n_20),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2131),
.Y(n_2308)
);

AOI22xp33_ASAP7_75t_L g2309 ( 
.A1(n_2130),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_2309)
);

AOI22xp33_ASAP7_75t_SL g2310 ( 
.A1(n_2175),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2179),
.Y(n_2311)
);

OR2x2_ASAP7_75t_L g2312 ( 
.A(n_2186),
.B(n_26),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2125),
.Y(n_2313)
);

O2A1O1Ixp33_ASAP7_75t_L g2314 ( 
.A1(n_2127),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2210),
.Y(n_2315)
);

AOI221xp5_ASAP7_75t_L g2316 ( 
.A1(n_2137),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.C(n_30),
.Y(n_2316)
);

AO21x1_ASAP7_75t_L g2317 ( 
.A1(n_2171),
.A2(n_31),
.B(n_30),
.Y(n_2317)
);

OAI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2239),
.A2(n_832),
.B(n_831),
.Y(n_2318)
);

O2A1O1Ixp33_ASAP7_75t_L g2319 ( 
.A1(n_2126),
.A2(n_32),
.B(n_29),
.C(n_31),
.Y(n_2319)
);

AOI22xp33_ASAP7_75t_L g2320 ( 
.A1(n_2230),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_2320)
);

AO31x2_ASAP7_75t_L g2321 ( 
.A1(n_2159),
.A2(n_835),
.A3(n_836),
.B(n_833),
.Y(n_2321)
);

OAI21x1_ASAP7_75t_L g2322 ( 
.A1(n_2234),
.A2(n_839),
.B(n_838),
.Y(n_2322)
);

BUFx3_ASAP7_75t_L g2323 ( 
.A(n_2188),
.Y(n_2323)
);

AO21x2_ASAP7_75t_L g2324 ( 
.A1(n_2218),
.A2(n_841),
.B(n_840),
.Y(n_2324)
);

OAI21x1_ASAP7_75t_L g2325 ( 
.A1(n_2253),
.A2(n_2271),
.B(n_2198),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2204),
.Y(n_2326)
);

AO21x2_ASAP7_75t_L g2327 ( 
.A1(n_2173),
.A2(n_844),
.B(n_842),
.Y(n_2327)
);

INVx3_ASAP7_75t_SL g2328 ( 
.A(n_2191),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2249),
.Y(n_2329)
);

INVxp67_ASAP7_75t_L g2330 ( 
.A(n_2145),
.Y(n_2330)
);

O2A1O1Ixp5_ASAP7_75t_L g2331 ( 
.A1(n_2170),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_2331)
);

BUFx2_ASAP7_75t_R g2332 ( 
.A(n_2163),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2243),
.Y(n_2333)
);

BUFx10_ASAP7_75t_L g2334 ( 
.A(n_2140),
.Y(n_2334)
);

OAI21x1_ASAP7_75t_L g2335 ( 
.A1(n_2254),
.A2(n_846),
.B(n_845),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2133),
.Y(n_2336)
);

OAI21x1_ASAP7_75t_L g2337 ( 
.A1(n_2134),
.A2(n_848),
.B(n_847),
.Y(n_2337)
);

AO31x2_ASAP7_75t_L g2338 ( 
.A1(n_2174),
.A2(n_2155),
.A3(n_2169),
.B(n_2147),
.Y(n_2338)
);

CKINVDCx8_ASAP7_75t_R g2339 ( 
.A(n_2191),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2139),
.Y(n_2340)
);

CKINVDCx20_ASAP7_75t_R g2341 ( 
.A(n_2146),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2128),
.B(n_36),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_L g2343 ( 
.A(n_2193),
.B(n_36),
.Y(n_2343)
);

AND2x6_ASAP7_75t_L g2344 ( 
.A(n_2245),
.B(n_852),
.Y(n_2344)
);

AOI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2252),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2345)
);

INVx4_ASAP7_75t_L g2346 ( 
.A(n_2188),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2255),
.Y(n_2347)
);

INVx4_ASAP7_75t_L g2348 ( 
.A(n_2267),
.Y(n_2348)
);

AOI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_2148),
.A2(n_855),
.B(n_853),
.Y(n_2349)
);

AOI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2199),
.A2(n_858),
.B(n_856),
.Y(n_2350)
);

AO31x2_ASAP7_75t_L g2351 ( 
.A1(n_2256),
.A2(n_860),
.A3(n_862),
.B(n_859),
.Y(n_2351)
);

OAI21x1_ASAP7_75t_L g2352 ( 
.A1(n_2246),
.A2(n_865),
.B(n_863),
.Y(n_2352)
);

AOI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_2221),
.A2(n_868),
.B(n_866),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2217),
.Y(n_2354)
);

OAI21x1_ASAP7_75t_L g2355 ( 
.A1(n_2178),
.A2(n_871),
.B(n_870),
.Y(n_2355)
);

AO21x2_ASAP7_75t_L g2356 ( 
.A1(n_2263),
.A2(n_873),
.B(n_872),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_2172),
.B(n_876),
.Y(n_2357)
);

AOI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2129),
.A2(n_2153),
.B(n_2141),
.Y(n_2358)
);

OAI211xp5_ASAP7_75t_L g2359 ( 
.A1(n_2248),
.A2(n_40),
.B(n_37),
.C(n_39),
.Y(n_2359)
);

INVx1_ASAP7_75t_SL g2360 ( 
.A(n_2220),
.Y(n_2360)
);

OAI21x1_ASAP7_75t_L g2361 ( 
.A1(n_2215),
.A2(n_879),
.B(n_878),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2219),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2225),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_2233),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2180),
.B(n_41),
.Y(n_2365)
);

AND2x4_ASAP7_75t_L g2366 ( 
.A(n_2233),
.B(n_880),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2189),
.B(n_41),
.Y(n_2367)
);

OA21x2_ASAP7_75t_L g2368 ( 
.A1(n_2135),
.A2(n_883),
.B(n_882),
.Y(n_2368)
);

HB1xp67_ASAP7_75t_L g2369 ( 
.A(n_2240),
.Y(n_2369)
);

OAI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2227),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2157),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2231),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2165),
.B(n_42),
.Y(n_2373)
);

OA21x2_ASAP7_75t_L g2374 ( 
.A1(n_2183),
.A2(n_885),
.B(n_884),
.Y(n_2374)
);

AOI222xp33_ASAP7_75t_L g2375 ( 
.A1(n_2132),
.A2(n_46),
.B1(n_48),
.B2(n_44),
.C1(n_45),
.C2(n_47),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2244),
.Y(n_2376)
);

NAND2x1p5_ASAP7_75t_L g2377 ( 
.A(n_2267),
.B(n_889),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2160),
.B(n_45),
.Y(n_2378)
);

OAI21x1_ASAP7_75t_L g2379 ( 
.A1(n_2209),
.A2(n_887),
.B(n_886),
.Y(n_2379)
);

OAI21x1_ASAP7_75t_SL g2380 ( 
.A1(n_2241),
.A2(n_893),
.B(n_888),
.Y(n_2380)
);

OAI22xp5_ASAP7_75t_L g2381 ( 
.A1(n_2166),
.A2(n_49),
.B1(n_46),
.B2(n_48),
.Y(n_2381)
);

NAND2x1p5_ASAP7_75t_L g2382 ( 
.A(n_2258),
.B(n_904),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2229),
.Y(n_2383)
);

OAI21x1_ASAP7_75t_L g2384 ( 
.A1(n_2223),
.A2(n_899),
.B(n_896),
.Y(n_2384)
);

AOI21x1_ASAP7_75t_L g2385 ( 
.A1(n_2201),
.A2(n_901),
.B(n_900),
.Y(n_2385)
);

OAI21x1_ASAP7_75t_L g2386 ( 
.A1(n_2261),
.A2(n_903),
.B(n_902),
.Y(n_2386)
);

AO21x2_ASAP7_75t_L g2387 ( 
.A1(n_2176),
.A2(n_908),
.B(n_905),
.Y(n_2387)
);

CKINVDCx8_ASAP7_75t_R g2388 ( 
.A(n_2277),
.Y(n_2388)
);

AO31x2_ASAP7_75t_L g2389 ( 
.A1(n_2264),
.A2(n_910),
.A3(n_911),
.B(n_909),
.Y(n_2389)
);

OAI21x1_ASAP7_75t_L g2390 ( 
.A1(n_2268),
.A2(n_917),
.B(n_913),
.Y(n_2390)
);

OAI22xp33_ASAP7_75t_L g2391 ( 
.A1(n_2274),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_2391)
);

AOI21x1_ASAP7_75t_L g2392 ( 
.A1(n_2192),
.A2(n_920),
.B(n_919),
.Y(n_2392)
);

AOI221xp5_ASAP7_75t_L g2393 ( 
.A1(n_2242),
.A2(n_54),
.B1(n_50),
.B2(n_52),
.C(n_55),
.Y(n_2393)
);

OAI21x1_ASAP7_75t_L g2394 ( 
.A1(n_2275),
.A2(n_922),
.B(n_921),
.Y(n_2394)
);

AOI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_2167),
.A2(n_925),
.B(n_924),
.Y(n_2395)
);

INVxp67_ASAP7_75t_L g2396 ( 
.A(n_2277),
.Y(n_2396)
);

OAI21x1_ASAP7_75t_L g2397 ( 
.A1(n_2138),
.A2(n_927),
.B(n_926),
.Y(n_2397)
);

OAI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2262),
.A2(n_55),
.B1(n_52),
.B2(n_54),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2237),
.B(n_56),
.Y(n_2399)
);

INVxp67_ASAP7_75t_L g2400 ( 
.A(n_2213),
.Y(n_2400)
);

BUFx3_ASAP7_75t_L g2401 ( 
.A(n_2260),
.Y(n_2401)
);

OAI22xp33_ASAP7_75t_L g2402 ( 
.A1(n_2274),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2402)
);

AOI221xp5_ASAP7_75t_L g2403 ( 
.A1(n_2257),
.A2(n_61),
.B1(n_58),
.B2(n_59),
.C(n_62),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_2236),
.Y(n_2404)
);

OAI21x1_ASAP7_75t_L g2405 ( 
.A1(n_2265),
.A2(n_933),
.B(n_928),
.Y(n_2405)
);

O2A1O1Ixp33_ASAP7_75t_SL g2406 ( 
.A1(n_2200),
.A2(n_935),
.B(n_938),
.C(n_934),
.Y(n_2406)
);

OAI22xp5_ASAP7_75t_L g2407 ( 
.A1(n_2197),
.A2(n_2238),
.B1(n_2272),
.B2(n_2216),
.Y(n_2407)
);

OAI21x1_ASAP7_75t_L g2408 ( 
.A1(n_2196),
.A2(n_2212),
.B(n_2208),
.Y(n_2408)
);

INVx2_ASAP7_75t_SL g2409 ( 
.A(n_2205),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2229),
.Y(n_2410)
);

AND2x4_ASAP7_75t_L g2411 ( 
.A(n_2247),
.B(n_940),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2244),
.Y(n_2412)
);

AOI21xp5_ASAP7_75t_L g2413 ( 
.A1(n_2276),
.A2(n_942),
.B(n_941),
.Y(n_2413)
);

OAI21x1_ASAP7_75t_L g2414 ( 
.A1(n_2222),
.A2(n_944),
.B(n_943),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_2251),
.Y(n_2415)
);

AOI21xp5_ASAP7_75t_L g2416 ( 
.A1(n_2228),
.A2(n_946),
.B(n_945),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2235),
.Y(n_2417)
);

INVx1_ASAP7_75t_SL g2418 ( 
.A(n_2270),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2168),
.B(n_947),
.Y(n_2419)
);

HB1xp67_ASAP7_75t_L g2420 ( 
.A(n_2235),
.Y(n_2420)
);

OAI21x1_ASAP7_75t_L g2421 ( 
.A1(n_2226),
.A2(n_952),
.B(n_951),
.Y(n_2421)
);

BUFx6f_ASAP7_75t_L g2422 ( 
.A(n_2185),
.Y(n_2422)
);

OAI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2270),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2207),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2185),
.Y(n_2425)
);

OA21x2_ASAP7_75t_L g2426 ( 
.A1(n_2250),
.A2(n_2207),
.B(n_2269),
.Y(n_2426)
);

AOI22x1_ASAP7_75t_L g2427 ( 
.A1(n_2269),
.A2(n_955),
.B1(n_956),
.B2(n_953),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2154),
.Y(n_2428)
);

OAI21x1_ASAP7_75t_L g2429 ( 
.A1(n_2156),
.A2(n_960),
.B(n_959),
.Y(n_2429)
);

BUFx3_ASAP7_75t_L g2430 ( 
.A(n_2152),
.Y(n_2430)
);

AND2x4_ASAP7_75t_L g2431 ( 
.A(n_2191),
.B(n_961),
.Y(n_2431)
);

OAI21x1_ASAP7_75t_L g2432 ( 
.A1(n_2156),
.A2(n_964),
.B(n_962),
.Y(n_2432)
);

BUFx10_ASAP7_75t_L g2433 ( 
.A(n_2140),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2161),
.B(n_63),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2154),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2278),
.Y(n_2436)
);

INVx3_ASAP7_75t_L g2437 ( 
.A(n_2388),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2294),
.Y(n_2438)
);

OAI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_2358),
.A2(n_64),
.B(n_65),
.Y(n_2439)
);

INVx4_ASAP7_75t_L g2440 ( 
.A(n_2328),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2428),
.Y(n_2441)
);

OAI21x1_ASAP7_75t_L g2442 ( 
.A1(n_2280),
.A2(n_966),
.B(n_965),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2333),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2435),
.Y(n_2444)
);

OA21x2_ASAP7_75t_L g2445 ( 
.A1(n_2424),
.A2(n_969),
.B(n_967),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2365),
.B(n_64),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2292),
.Y(n_2447)
);

AO21x2_ASAP7_75t_L g2448 ( 
.A1(n_2417),
.A2(n_975),
.B(n_973),
.Y(n_2448)
);

CKINVDCx16_ASAP7_75t_R g2449 ( 
.A(n_2341),
.Y(n_2449)
);

AO31x2_ASAP7_75t_L g2450 ( 
.A1(n_2383),
.A2(n_977),
.A3(n_978),
.B(n_976),
.Y(n_2450)
);

AOI21x1_ASAP7_75t_L g2451 ( 
.A1(n_2306),
.A2(n_980),
.B(n_979),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2347),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2326),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2329),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2302),
.Y(n_2455)
);

AO21x2_ASAP7_75t_L g2456 ( 
.A1(n_2410),
.A2(n_986),
.B(n_985),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2372),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2343),
.B(n_67),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2362),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2315),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2363),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2354),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_2339),
.Y(n_2463)
);

INVx2_ASAP7_75t_SL g2464 ( 
.A(n_2364),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2287),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2284),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2288),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2313),
.Y(n_2468)
);

HB1xp67_ASAP7_75t_L g2469 ( 
.A(n_2330),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2434),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_L g2471 ( 
.A(n_2286),
.B(n_987),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2422),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2422),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2336),
.Y(n_2474)
);

AND2x4_ASAP7_75t_L g2475 ( 
.A(n_2311),
.B(n_988),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2400),
.B(n_67),
.Y(n_2476)
);

INVxp67_ASAP7_75t_L g2477 ( 
.A(n_2369),
.Y(n_2477)
);

NOR2x1_ASAP7_75t_L g2478 ( 
.A(n_2348),
.B(n_989),
.Y(n_2478)
);

BUFx3_ASAP7_75t_L g2479 ( 
.A(n_2364),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2308),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2371),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2425),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2317),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2367),
.B(n_68),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2342),
.Y(n_2485)
);

BUFx8_ASAP7_75t_SL g2486 ( 
.A(n_2415),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2378),
.B(n_69),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2352),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2373),
.B(n_70),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2340),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2296),
.B(n_70),
.Y(n_2491)
);

HB1xp67_ASAP7_75t_L g2492 ( 
.A(n_2404),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2279),
.Y(n_2493)
);

HB1xp67_ASAP7_75t_L g2494 ( 
.A(n_2404),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2289),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_2323),
.B(n_990),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2296),
.B(n_71),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2296),
.B(n_72),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2331),
.Y(n_2499)
);

HB1xp67_ASAP7_75t_L g2500 ( 
.A(n_2396),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2376),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_L g2502 ( 
.A1(n_2375),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_2502)
);

BUFx2_ASAP7_75t_L g2503 ( 
.A(n_2418),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2412),
.Y(n_2504)
);

BUFx3_ASAP7_75t_L g2505 ( 
.A(n_2298),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2385),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2307),
.Y(n_2507)
);

HB1xp67_ASAP7_75t_L g2508 ( 
.A(n_2360),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2411),
.B(n_74),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2312),
.Y(n_2510)
);

INVx2_ASAP7_75t_SL g2511 ( 
.A(n_2334),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2399),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2335),
.Y(n_2513)
);

OAI21x1_ASAP7_75t_L g2514 ( 
.A1(n_2325),
.A2(n_992),
.B(n_991),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2295),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2291),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2366),
.B(n_75),
.Y(n_2517)
);

HB1xp67_ASAP7_75t_L g2518 ( 
.A(n_2346),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2405),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2392),
.Y(n_2520)
);

HB1xp67_ASAP7_75t_L g2521 ( 
.A(n_2357),
.Y(n_2521)
);

BUFx3_ASAP7_75t_L g2522 ( 
.A(n_2401),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_2433),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2285),
.Y(n_2524)
);

BUFx12f_ASAP7_75t_L g2525 ( 
.A(n_2409),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2381),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2386),
.Y(n_2527)
);

INVx3_ASAP7_75t_L g2528 ( 
.A(n_2430),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2390),
.Y(n_2529)
);

NAND2x1p5_ASAP7_75t_L g2530 ( 
.A(n_2431),
.B(n_993),
.Y(n_2530)
);

BUFx3_ASAP7_75t_L g2531 ( 
.A(n_2303),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2394),
.Y(n_2532)
);

NOR2xp33_ASAP7_75t_L g2533 ( 
.A(n_2283),
.B(n_2290),
.Y(n_2533)
);

AND2x6_ASAP7_75t_L g2534 ( 
.A(n_2419),
.B(n_995),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2389),
.Y(n_2535)
);

AOI22xp33_ASAP7_75t_L g2536 ( 
.A1(n_2320),
.A2(n_2393),
.B1(n_2403),
.B2(n_2316),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2379),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2384),
.Y(n_2538)
);

INVx4_ASAP7_75t_L g2539 ( 
.A(n_2344),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2468),
.Y(n_2540)
);

XOR2xp5_ASAP7_75t_L g2541 ( 
.A(n_2449),
.B(n_2332),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_R g2542 ( 
.A(n_2437),
.B(n_2344),
.Y(n_2542)
);

BUFx5_ASAP7_75t_L g2543 ( 
.A(n_2519),
.Y(n_2543)
);

AND2x4_ASAP7_75t_L g2544 ( 
.A(n_2522),
.B(n_2281),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2492),
.B(n_2344),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_R g2546 ( 
.A(n_2463),
.B(n_2293),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2470),
.B(n_2309),
.Y(n_2547)
);

INVxp67_ASAP7_75t_L g2548 ( 
.A(n_2469),
.Y(n_2548)
);

INVx3_ASAP7_75t_L g2549 ( 
.A(n_2505),
.Y(n_2549)
);

OR2x6_ASAP7_75t_L g2550 ( 
.A(n_2539),
.B(n_2377),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_R g2551 ( 
.A(n_2479),
.B(n_2305),
.Y(n_2551)
);

BUFx3_ASAP7_75t_L g2552 ( 
.A(n_2525),
.Y(n_2552)
);

NAND2xp33_ASAP7_75t_R g2553 ( 
.A(n_2528),
.B(n_2426),
.Y(n_2553)
);

NAND2xp33_ASAP7_75t_R g2554 ( 
.A(n_2523),
.B(n_2374),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2485),
.B(n_2423),
.Y(n_2555)
);

OR2x6_ASAP7_75t_L g2556 ( 
.A(n_2530),
.B(n_2382),
.Y(n_2556)
);

AND2x4_ASAP7_75t_L g2557 ( 
.A(n_2494),
.B(n_2397),
.Y(n_2557)
);

NAND2xp33_ASAP7_75t_R g2558 ( 
.A(n_2533),
.B(n_2368),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_R g2559 ( 
.A(n_2464),
.B(n_2299),
.Y(n_2559)
);

NOR2xp33_ASAP7_75t_R g2560 ( 
.A(n_2531),
.B(n_2420),
.Y(n_2560)
);

INVxp67_ASAP7_75t_L g2561 ( 
.A(n_2508),
.Y(n_2561)
);

XNOR2xp5_ASAP7_75t_L g2562 ( 
.A(n_2509),
.B(n_2300),
.Y(n_2562)
);

NAND2xp33_ASAP7_75t_R g2563 ( 
.A(n_2496),
.B(n_2318),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_R g2564 ( 
.A(n_2440),
.B(n_996),
.Y(n_2564)
);

INVxp67_ASAP7_75t_L g2565 ( 
.A(n_2500),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2507),
.B(n_2345),
.Y(n_2566)
);

XNOR2xp5_ASAP7_75t_L g2567 ( 
.A(n_2521),
.B(n_2391),
.Y(n_2567)
);

CKINVDCx5p33_ASAP7_75t_R g2568 ( 
.A(n_2486),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2438),
.Y(n_2569)
);

NAND2xp33_ASAP7_75t_R g2570 ( 
.A(n_2496),
.B(n_2408),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2443),
.Y(n_2571)
);

BUFx3_ASAP7_75t_L g2572 ( 
.A(n_2511),
.Y(n_2572)
);

BUFx3_ASAP7_75t_L g2573 ( 
.A(n_2518),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2455),
.Y(n_2574)
);

AND2x4_ASAP7_75t_L g2575 ( 
.A(n_2477),
.B(n_2297),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_R g2576 ( 
.A(n_2510),
.B(n_997),
.Y(n_2576)
);

NAND2xp33_ASAP7_75t_R g2577 ( 
.A(n_2471),
.B(n_2414),
.Y(n_2577)
);

NAND2xp33_ASAP7_75t_R g2578 ( 
.A(n_2458),
.B(n_2421),
.Y(n_2578)
);

NOR2xp33_ASAP7_75t_R g2579 ( 
.A(n_2534),
.B(n_1000),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_R g2580 ( 
.A(n_2534),
.B(n_1001),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2512),
.B(n_2407),
.Y(n_2581)
);

AND2x4_ASAP7_75t_L g2582 ( 
.A(n_2475),
.B(n_2351),
.Y(n_2582)
);

BUFx12f_ASAP7_75t_L g2583 ( 
.A(n_2534),
.Y(n_2583)
);

BUFx10_ASAP7_75t_L g2584 ( 
.A(n_2475),
.Y(n_2584)
);

NAND2xp33_ASAP7_75t_SL g2585 ( 
.A(n_2502),
.B(n_2398),
.Y(n_2585)
);

XNOR2xp5_ASAP7_75t_L g2586 ( 
.A(n_2517),
.B(n_2402),
.Y(n_2586)
);

NAND2xp33_ASAP7_75t_R g2587 ( 
.A(n_2491),
.B(n_2350),
.Y(n_2587)
);

NAND2xp33_ASAP7_75t_R g2588 ( 
.A(n_2497),
.B(n_2353),
.Y(n_2588)
);

AND2x2_ASAP7_75t_SL g2589 ( 
.A(n_2536),
.B(n_2319),
.Y(n_2589)
);

NAND2xp33_ASAP7_75t_R g2590 ( 
.A(n_2498),
.B(n_2395),
.Y(n_2590)
);

AND2x4_ASAP7_75t_L g2591 ( 
.A(n_2436),
.B(n_2351),
.Y(n_2591)
);

NAND2xp33_ASAP7_75t_R g2592 ( 
.A(n_2476),
.B(n_2349),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2452),
.Y(n_2593)
);

XNOR2xp5_ASAP7_75t_L g2594 ( 
.A(n_2446),
.B(n_2310),
.Y(n_2594)
);

NAND3xp33_ASAP7_75t_SL g2595 ( 
.A(n_2439),
.B(n_2314),
.C(n_2359),
.Y(n_2595)
);

AND2x4_ASAP7_75t_L g2596 ( 
.A(n_2441),
.B(n_2356),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2526),
.B(n_2304),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2453),
.Y(n_2598)
);

NAND2xp33_ASAP7_75t_R g2599 ( 
.A(n_2503),
.B(n_2416),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2548),
.B(n_2503),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2569),
.Y(n_2601)
);

OR2x2_ASAP7_75t_L g2602 ( 
.A(n_2571),
.B(n_2501),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2593),
.B(n_2598),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2575),
.B(n_2472),
.Y(n_2604)
);

HB1xp67_ASAP7_75t_L g2605 ( 
.A(n_2540),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2574),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2544),
.B(n_2473),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2591),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2543),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2561),
.B(n_2484),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2565),
.B(n_2487),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2581),
.B(n_2459),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2543),
.Y(n_2613)
);

AOI22xp33_ASAP7_75t_L g2614 ( 
.A1(n_2589),
.A2(n_2370),
.B1(n_2489),
.B2(n_2324),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2543),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2543),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2566),
.B(n_2461),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2582),
.B(n_2504),
.Y(n_2618)
);

BUFx3_ASAP7_75t_L g2619 ( 
.A(n_2549),
.Y(n_2619)
);

AOI22xp33_ASAP7_75t_L g2620 ( 
.A1(n_2585),
.A2(n_2483),
.B1(n_2478),
.B2(n_2490),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2596),
.Y(n_2621)
);

OR2x2_ASAP7_75t_L g2622 ( 
.A(n_2555),
.B(n_2482),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2573),
.B(n_2447),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2562),
.B(n_2457),
.Y(n_2624)
);

OAI21xp5_ASAP7_75t_L g2625 ( 
.A1(n_2595),
.A2(n_2413),
.B(n_2499),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2557),
.B(n_2481),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2545),
.B(n_2462),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2560),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2584),
.Y(n_2629)
);

OR2x2_ASAP7_75t_L g2630 ( 
.A(n_2547),
.B(n_2474),
.Y(n_2630)
);

OR2x2_ASAP7_75t_L g2631 ( 
.A(n_2597),
.B(n_2535),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2567),
.B(n_2465),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2572),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2546),
.B(n_2466),
.Y(n_2634)
);

AND2x4_ASAP7_75t_L g2635 ( 
.A(n_2552),
.B(n_2495),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2550),
.Y(n_2636)
);

HB1xp67_ASAP7_75t_L g2637 ( 
.A(n_2553),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2550),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_2579),
.B(n_2480),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2556),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2594),
.B(n_2444),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2576),
.B(n_2467),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2586),
.B(n_2454),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2583),
.Y(n_2644)
);

HB1xp67_ASAP7_75t_L g2645 ( 
.A(n_2570),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2556),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2554),
.Y(n_2647)
);

OR2x2_ASAP7_75t_L g2648 ( 
.A(n_2541),
.B(n_2524),
.Y(n_2648)
);

OR2x2_ASAP7_75t_L g2649 ( 
.A(n_2578),
.B(n_2515),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2542),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2558),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2599),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2580),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2551),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2590),
.Y(n_2655)
);

AOI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_2564),
.A2(n_2427),
.B1(n_2380),
.B2(n_2448),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2577),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2587),
.Y(n_2658)
);

AOI22xp33_ASAP7_75t_L g2659 ( 
.A1(n_2559),
.A2(n_2456),
.B1(n_2387),
.B2(n_2527),
.Y(n_2659)
);

OAI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2563),
.A2(n_2460),
.B1(n_2506),
.B2(n_2445),
.Y(n_2660)
);

HB1xp67_ASAP7_75t_L g2661 ( 
.A(n_2605),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_SL g2662 ( 
.A(n_2655),
.B(n_2568),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2657),
.B(n_2651),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2601),
.Y(n_2664)
);

AND2x4_ASAP7_75t_L g2665 ( 
.A(n_2618),
.B(n_2516),
.Y(n_2665)
);

AND2x4_ASAP7_75t_SL g2666 ( 
.A(n_2642),
.B(n_2532),
.Y(n_2666)
);

OR2x2_ASAP7_75t_L g2667 ( 
.A(n_2657),
.B(n_2493),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2602),
.Y(n_2668)
);

BUFx2_ASAP7_75t_L g2669 ( 
.A(n_2647),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2603),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2606),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2631),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2622),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2658),
.B(n_2645),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2623),
.B(n_2520),
.Y(n_2675)
);

OAI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2614),
.A2(n_2445),
.B1(n_2537),
.B2(n_2529),
.Y(n_2676)
);

AOI222xp33_ASAP7_75t_L g2677 ( 
.A1(n_2625),
.A2(n_2592),
.B1(n_2588),
.B2(n_104),
.C1(n_85),
.C2(n_112),
.Y(n_2677)
);

NAND3xp33_ASAP7_75t_L g2678 ( 
.A(n_2620),
.B(n_2406),
.C(n_2538),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2652),
.B(n_2321),
.Y(n_2679)
);

AO21x2_ASAP7_75t_L g2680 ( 
.A1(n_2615),
.A2(n_2451),
.B(n_2488),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2600),
.B(n_2321),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2612),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2648),
.B(n_2450),
.Y(n_2683)
);

AND2x2_ASAP7_75t_SL g2684 ( 
.A(n_2637),
.B(n_2513),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2621),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2616),
.Y(n_2686)
);

INVxp67_ASAP7_75t_SL g2687 ( 
.A(n_2649),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2617),
.Y(n_2688)
);

INVx1_ASAP7_75t_SL g2689 ( 
.A(n_2619),
.Y(n_2689)
);

NAND2x1_ASAP7_75t_L g2690 ( 
.A(n_2609),
.B(n_2450),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2608),
.Y(n_2691)
);

INVxp67_ASAP7_75t_SL g2692 ( 
.A(n_2613),
.Y(n_2692)
);

NOR2xp33_ASAP7_75t_L g2693 ( 
.A(n_2654),
.B(n_2650),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2630),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2628),
.B(n_2514),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2611),
.B(n_2442),
.Y(n_2696)
);

OAI33xp33_ASAP7_75t_L g2697 ( 
.A1(n_2632),
.A2(n_78),
.A3(n_81),
.B1(n_76),
.B2(n_77),
.B3(n_79),
.Y(n_2697)
);

INVx2_ASAP7_75t_SL g2698 ( 
.A(n_2633),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2610),
.B(n_2327),
.Y(n_2699)
);

AOI22xp33_ASAP7_75t_L g2700 ( 
.A1(n_2654),
.A2(n_2337),
.B1(n_2301),
.B2(n_2429),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_2653),
.A2(n_2432),
.B1(n_2361),
.B2(n_2355),
.Y(n_2701)
);

OR2x2_ASAP7_75t_L g2702 ( 
.A(n_2640),
.B(n_2338),
.Y(n_2702)
);

NAND4xp25_ASAP7_75t_L g2703 ( 
.A(n_2641),
.B(n_79),
.C(n_76),
.D(n_77),
.Y(n_2703)
);

BUFx6f_ASAP7_75t_L g2704 ( 
.A(n_2629),
.Y(n_2704)
);

HB1xp67_ASAP7_75t_L g2705 ( 
.A(n_2638),
.Y(n_2705)
);

OAI31xp33_ASAP7_75t_L g2706 ( 
.A1(n_2639),
.A2(n_84),
.A3(n_82),
.B(n_83),
.Y(n_2706)
);

INVx3_ASAP7_75t_L g2707 ( 
.A(n_2635),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2626),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2638),
.Y(n_2709)
);

INVx3_ASAP7_75t_L g2710 ( 
.A(n_2635),
.Y(n_2710)
);

OAI33xp33_ASAP7_75t_L g2711 ( 
.A1(n_2660),
.A2(n_84),
.A3(n_87),
.B1(n_82),
.B2(n_83),
.B3(n_86),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2626),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2624),
.B(n_2451),
.Y(n_2713)
);

NAND4xp25_ASAP7_75t_SL g2714 ( 
.A(n_2653),
.B(n_90),
.C(n_86),
.D(n_88),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2636),
.Y(n_2715)
);

AOI22xp33_ASAP7_75t_L g2716 ( 
.A1(n_2646),
.A2(n_2322),
.B1(n_2282),
.B2(n_93),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2627),
.Y(n_2717)
);

INVx4_ASAP7_75t_L g2718 ( 
.A(n_2634),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2604),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2607),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2643),
.B(n_2389),
.Y(n_2721)
);

INVx2_ASAP7_75t_SL g2722 ( 
.A(n_2644),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2659),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2656),
.B(n_2338),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2601),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2601),
.Y(n_2726)
);

BUFx2_ASAP7_75t_L g2727 ( 
.A(n_2640),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2655),
.B(n_91),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2605),
.Y(n_2729)
);

INVx2_ASAP7_75t_SL g2730 ( 
.A(n_2619),
.Y(n_2730)
);

CKINVDCx16_ASAP7_75t_R g2731 ( 
.A(n_2619),
.Y(n_2731)
);

OAI33xp33_ASAP7_75t_L g2732 ( 
.A1(n_2617),
.A2(n_94),
.A3(n_97),
.B1(n_91),
.B2(n_92),
.B3(n_95),
.Y(n_2732)
);

INVx2_ASAP7_75t_SL g2733 ( 
.A(n_2619),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2655),
.B(n_92),
.Y(n_2734)
);

NAND2x1_ASAP7_75t_L g2735 ( 
.A(n_2655),
.B(n_94),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2601),
.Y(n_2736)
);

OR2x2_ASAP7_75t_L g2737 ( 
.A(n_2651),
.B(n_97),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2657),
.B(n_98),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_2619),
.Y(n_2739)
);

NOR2xp33_ASAP7_75t_L g2740 ( 
.A(n_2654),
.B(n_99),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2655),
.B(n_99),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2601),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2669),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2682),
.B(n_100),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2661),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2664),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2674),
.B(n_100),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2688),
.B(n_2663),
.Y(n_2748)
);

HB1xp67_ASAP7_75t_L g2749 ( 
.A(n_2669),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2694),
.B(n_2672),
.Y(n_2750)
);

OR2x2_ASAP7_75t_L g2751 ( 
.A(n_2687),
.B(n_102),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2727),
.B(n_103),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2729),
.Y(n_2753)
);

INVx2_ASAP7_75t_SL g2754 ( 
.A(n_2731),
.Y(n_2754)
);

AND2x4_ASAP7_75t_L g2755 ( 
.A(n_2707),
.B(n_105),
.Y(n_2755)
);

BUFx2_ASAP7_75t_L g2756 ( 
.A(n_2710),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2718),
.B(n_105),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2673),
.B(n_106),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_2677),
.B(n_107),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_L g2760 ( 
.A(n_2662),
.B(n_107),
.Y(n_2760)
);

HB1xp67_ASAP7_75t_L g2761 ( 
.A(n_2667),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2725),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2726),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2668),
.B(n_108),
.Y(n_2764)
);

HB1xp67_ASAP7_75t_L g2765 ( 
.A(n_2705),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2675),
.B(n_108),
.Y(n_2766)
);

HB1xp67_ASAP7_75t_L g2767 ( 
.A(n_2709),
.Y(n_2767)
);

OR2x2_ASAP7_75t_L g2768 ( 
.A(n_2702),
.B(n_109),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2720),
.B(n_109),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2736),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2670),
.B(n_110),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2719),
.B(n_110),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2715),
.B(n_2717),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2686),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2713),
.B(n_111),
.Y(n_2775)
);

NOR2xp33_ASAP7_75t_L g2776 ( 
.A(n_2704),
.B(n_111),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2723),
.B(n_113),
.Y(n_2777)
);

OR2x2_ASAP7_75t_L g2778 ( 
.A(n_2692),
.B(n_113),
.Y(n_2778)
);

INVxp33_ASAP7_75t_L g2779 ( 
.A(n_2693),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2671),
.B(n_114),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2708),
.B(n_115),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2742),
.Y(n_2782)
);

AND2x4_ASAP7_75t_L g2783 ( 
.A(n_2712),
.B(n_117),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2691),
.B(n_118),
.Y(n_2784)
);

INVxp67_ASAP7_75t_L g2785 ( 
.A(n_2728),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2685),
.B(n_118),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2683),
.B(n_119),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2681),
.Y(n_2788)
);

HB1xp67_ASAP7_75t_L g2789 ( 
.A(n_2699),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2684),
.B(n_120),
.Y(n_2790)
);

OR2x2_ASAP7_75t_L g2791 ( 
.A(n_2721),
.B(n_120),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2679),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2696),
.B(n_121),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2698),
.B(n_121),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2665),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2695),
.B(n_122),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_L g2797 ( 
.A(n_2704),
.B(n_2722),
.Y(n_2797)
);

INVx2_ASAP7_75t_SL g2798 ( 
.A(n_2739),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2738),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2724),
.B(n_123),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2666),
.Y(n_2801)
);

AND2x4_ASAP7_75t_L g2802 ( 
.A(n_2730),
.B(n_124),
.Y(n_2802)
);

INVx2_ASAP7_75t_SL g2803 ( 
.A(n_2733),
.Y(n_2803)
);

AND2x2_ASAP7_75t_L g2804 ( 
.A(n_2689),
.B(n_2737),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2734),
.B(n_124),
.Y(n_2805)
);

HB1xp67_ASAP7_75t_L g2806 ( 
.A(n_2690),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2741),
.B(n_125),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2680),
.Y(n_2808)
);

INVxp67_ASAP7_75t_L g2809 ( 
.A(n_2740),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2735),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2676),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2703),
.B(n_2678),
.Y(n_2812)
);

OR2x2_ASAP7_75t_L g2813 ( 
.A(n_2716),
.B(n_125),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2701),
.Y(n_2814)
);

OR2x6_ASAP7_75t_L g2815 ( 
.A(n_2714),
.B(n_2711),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2700),
.B(n_126),
.Y(n_2816)
);

OAI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2697),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2732),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2706),
.B(n_128),
.Y(n_2819)
);

NAND2x1_ASAP7_75t_L g2820 ( 
.A(n_2669),
.B(n_129),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2669),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2674),
.B(n_129),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2661),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_L g2824 ( 
.A1(n_2677),
.A2(n_1005),
.B(n_1004),
.Y(n_2824)
);

AOI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2677),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2661),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2661),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2669),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2661),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2661),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2674),
.B(n_130),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2674),
.B(n_133),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2661),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2674),
.B(n_134),
.Y(n_2834)
);

OR2x2_ASAP7_75t_L g2835 ( 
.A(n_2687),
.B(n_134),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2682),
.B(n_135),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2661),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2674),
.B(n_135),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2682),
.B(n_136),
.Y(n_2839)
);

AND2x2_ASAP7_75t_L g2840 ( 
.A(n_2674),
.B(n_136),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2674),
.B(n_138),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2669),
.Y(n_2842)
);

NAND2x1p5_ASAP7_75t_L g2843 ( 
.A(n_2684),
.B(n_1006),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2674),
.B(n_138),
.Y(n_2844)
);

OR2x2_ASAP7_75t_L g2845 ( 
.A(n_2687),
.B(n_139),
.Y(n_2845)
);

INVxp67_ASAP7_75t_L g2846 ( 
.A(n_2705),
.Y(n_2846)
);

NAND2x1p5_ASAP7_75t_L g2847 ( 
.A(n_2684),
.B(n_1007),
.Y(n_2847)
);

NOR2xp33_ASAP7_75t_L g2848 ( 
.A(n_2718),
.B(n_139),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2669),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2674),
.B(n_140),
.Y(n_2850)
);

OAI21xp5_ASAP7_75t_L g2851 ( 
.A1(n_2677),
.A2(n_140),
.B(n_141),
.Y(n_2851)
);

AND2x2_ASAP7_75t_L g2852 ( 
.A(n_2674),
.B(n_141),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2674),
.B(n_142),
.Y(n_2853)
);

INVx3_ASAP7_75t_L g2854 ( 
.A(n_2704),
.Y(n_2854)
);

AND3x1_ASAP7_75t_L g2855 ( 
.A(n_2706),
.B(n_142),
.C(n_143),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_SL g2856 ( 
.A(n_2731),
.B(n_144),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2661),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2674),
.B(n_144),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2661),
.Y(n_2859)
);

AND2x4_ASAP7_75t_L g2860 ( 
.A(n_2754),
.B(n_145),
.Y(n_2860)
);

NAND2xp33_ASAP7_75t_SL g2861 ( 
.A(n_2820),
.B(n_145),
.Y(n_2861)
);

AO221x2_ASAP7_75t_L g2862 ( 
.A1(n_2851),
.A2(n_149),
.B1(n_151),
.B2(n_148),
.C(n_150),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2788),
.B(n_146),
.Y(n_2863)
);

NAND2xp33_ASAP7_75t_SL g2864 ( 
.A(n_2856),
.B(n_146),
.Y(n_2864)
);

CKINVDCx5p33_ASAP7_75t_R g2865 ( 
.A(n_2798),
.Y(n_2865)
);

AO221x2_ASAP7_75t_L g2866 ( 
.A1(n_2812),
.A2(n_151),
.B1(n_153),
.B2(n_149),
.C(n_152),
.Y(n_2866)
);

NAND2xp33_ASAP7_75t_SL g2867 ( 
.A(n_2790),
.B(n_148),
.Y(n_2867)
);

NAND2xp33_ASAP7_75t_SL g2868 ( 
.A(n_2779),
.B(n_152),
.Y(n_2868)
);

AOI22xp5_ASAP7_75t_L g2869 ( 
.A1(n_2759),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2869)
);

INVxp67_ASAP7_75t_L g2870 ( 
.A(n_2768),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2792),
.B(n_2745),
.Y(n_2871)
);

OAI22xp33_ASAP7_75t_L g2872 ( 
.A1(n_2824),
.A2(n_157),
.B1(n_154),
.B2(n_155),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2789),
.B(n_157),
.Y(n_2873)
);

NAND2xp33_ASAP7_75t_R g2874 ( 
.A(n_2810),
.B(n_158),
.Y(n_2874)
);

OAI221xp5_ASAP7_75t_L g2875 ( 
.A1(n_2825),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.C(n_162),
.Y(n_2875)
);

OR2x2_ASAP7_75t_L g2876 ( 
.A(n_2761),
.B(n_159),
.Y(n_2876)
);

BUFx2_ASAP7_75t_L g2877 ( 
.A(n_2749),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2814),
.B(n_160),
.Y(n_2878)
);

AO221x2_ASAP7_75t_L g2879 ( 
.A1(n_2817),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.C(n_164),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2823),
.B(n_163),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2743),
.Y(n_2881)
);

BUFx12f_ASAP7_75t_L g2882 ( 
.A(n_2805),
.Y(n_2882)
);

BUFx2_ASAP7_75t_L g2883 ( 
.A(n_2765),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_L g2884 ( 
.A(n_2785),
.B(n_164),
.Y(n_2884)
);

NOR2xp33_ASAP7_75t_L g2885 ( 
.A(n_2809),
.B(n_165),
.Y(n_2885)
);

AO221x2_ASAP7_75t_L g2886 ( 
.A1(n_2799),
.A2(n_167),
.B1(n_169),
.B2(n_166),
.C(n_168),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2826),
.B(n_165),
.Y(n_2887)
);

NOR2x1_ASAP7_75t_L g2888 ( 
.A(n_2751),
.B(n_166),
.Y(n_2888)
);

CKINVDCx5p33_ASAP7_75t_R g2889 ( 
.A(n_2803),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2821),
.Y(n_2890)
);

AND2x4_ASAP7_75t_L g2891 ( 
.A(n_2827),
.B(n_167),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2756),
.B(n_168),
.Y(n_2892)
);

A2O1A1Ixp33_ASAP7_75t_L g2893 ( 
.A1(n_2818),
.A2(n_177),
.B(n_185),
.C(n_169),
.Y(n_2893)
);

HB1xp67_ASAP7_75t_L g2894 ( 
.A(n_2767),
.Y(n_2894)
);

AO221x2_ASAP7_75t_L g2895 ( 
.A1(n_2777),
.A2(n_172),
.B1(n_174),
.B2(n_171),
.C(n_173),
.Y(n_2895)
);

CKINVDCx5p33_ASAP7_75t_R g2896 ( 
.A(n_2854),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2829),
.B(n_170),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2830),
.B(n_171),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2746),
.Y(n_2899)
);

AO221x2_ASAP7_75t_L g2900 ( 
.A1(n_2800),
.A2(n_175),
.B1(n_172),
.B2(n_173),
.C(n_176),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2833),
.B(n_175),
.Y(n_2901)
);

OAI22xp33_ASAP7_75t_L g2902 ( 
.A1(n_2815),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_2902)
);

AO221x2_ASAP7_75t_L g2903 ( 
.A1(n_2775),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.C(n_181),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2837),
.B(n_179),
.Y(n_2904)
);

NAND2xp33_ASAP7_75t_R g2905 ( 
.A(n_2802),
.B(n_180),
.Y(n_2905)
);

AO221x2_ASAP7_75t_L g2906 ( 
.A1(n_2794),
.A2(n_184),
.B1(n_186),
.B2(n_183),
.C(n_185),
.Y(n_2906)
);

AO221x2_ASAP7_75t_L g2907 ( 
.A1(n_2758),
.A2(n_186),
.B1(n_188),
.B2(n_184),
.C(n_187),
.Y(n_2907)
);

CKINVDCx16_ASAP7_75t_R g2908 ( 
.A(n_2804),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2857),
.B(n_182),
.Y(n_2909)
);

NOR2x1_ASAP7_75t_L g2910 ( 
.A(n_2835),
.B(n_2845),
.Y(n_2910)
);

AOI22xp5_ASAP7_75t_L g2911 ( 
.A1(n_2855),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_L g2912 ( 
.A(n_2791),
.B(n_189),
.Y(n_2912)
);

CKINVDCx5p33_ASAP7_75t_R g2913 ( 
.A(n_2802),
.Y(n_2913)
);

OAI221xp5_ASAP7_75t_L g2914 ( 
.A1(n_2815),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.C(n_193),
.Y(n_2914)
);

AND2x4_ASAP7_75t_L g2915 ( 
.A(n_2859),
.B(n_191),
.Y(n_2915)
);

OAI22xp5_ASAP7_75t_SL g2916 ( 
.A1(n_2757),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2748),
.B(n_195),
.Y(n_2917)
);

NOR2xp33_ASAP7_75t_SL g2918 ( 
.A(n_2843),
.B(n_197),
.Y(n_2918)
);

AOI22xp5_ASAP7_75t_L g2919 ( 
.A1(n_2819),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_2919)
);

AO221x2_ASAP7_75t_L g2920 ( 
.A1(n_2764),
.A2(n_201),
.B1(n_203),
.B2(n_200),
.C(n_202),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_R g2921 ( 
.A(n_2848),
.B(n_199),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2753),
.B(n_200),
.Y(n_2922)
);

AO221x2_ASAP7_75t_L g2923 ( 
.A1(n_2793),
.A2(n_205),
.B1(n_207),
.B2(n_203),
.C(n_206),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2774),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2828),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2750),
.B(n_202),
.Y(n_2926)
);

AOI22xp5_ASAP7_75t_SL g2927 ( 
.A1(n_2752),
.A2(n_211),
.B1(n_212),
.B2(n_208),
.Y(n_2927)
);

OAI22xp5_ASAP7_75t_SL g2928 ( 
.A1(n_2760),
.A2(n_212),
.B1(n_207),
.B2(n_211),
.Y(n_2928)
);

INVx1_ASAP7_75t_SL g2929 ( 
.A(n_2778),
.Y(n_2929)
);

NOR2x1_ASAP7_75t_L g2930 ( 
.A(n_2797),
.B(n_2744),
.Y(n_2930)
);

NAND2xp33_ASAP7_75t_SL g2931 ( 
.A(n_2747),
.B(n_213),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2846),
.B(n_213),
.Y(n_2932)
);

BUFx3_ASAP7_75t_L g2933 ( 
.A(n_2755),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2773),
.B(n_214),
.Y(n_2934)
);

NOR2x1_ASAP7_75t_L g2935 ( 
.A(n_2836),
.B(n_214),
.Y(n_2935)
);

AOI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_2811),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_2936)
);

OAI221xp5_ASAP7_75t_L g2937 ( 
.A1(n_2813),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.C(n_220),
.Y(n_2937)
);

INVxp67_ASAP7_75t_SL g2938 ( 
.A(n_2806),
.Y(n_2938)
);

OR2x2_ASAP7_75t_L g2939 ( 
.A(n_2842),
.B(n_219),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2762),
.B(n_220),
.Y(n_2940)
);

NOR2xp33_ASAP7_75t_L g2941 ( 
.A(n_2807),
.B(n_221),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2763),
.B(n_221),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2770),
.B(n_222),
.Y(n_2943)
);

INVxp33_ASAP7_75t_SL g2944 ( 
.A(n_2776),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2782),
.B(n_2849),
.Y(n_2945)
);

OR2x2_ASAP7_75t_L g2946 ( 
.A(n_2795),
.B(n_223),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2796),
.B(n_224),
.Y(n_2947)
);

NAND2x1_ASAP7_75t_L g2948 ( 
.A(n_2808),
.B(n_224),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2787),
.B(n_225),
.Y(n_2949)
);

CKINVDCx5p33_ASAP7_75t_R g2950 ( 
.A(n_2781),
.Y(n_2950)
);

OAI221xp5_ASAP7_75t_L g2951 ( 
.A1(n_2766),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.C(n_229),
.Y(n_2951)
);

CKINVDCx5p33_ASAP7_75t_R g2952 ( 
.A(n_2822),
.Y(n_2952)
);

CKINVDCx5p33_ASAP7_75t_R g2953 ( 
.A(n_2831),
.Y(n_2953)
);

OAI22xp33_ASAP7_75t_L g2954 ( 
.A1(n_2847),
.A2(n_231),
.B1(n_228),
.B2(n_230),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2771),
.B(n_230),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2839),
.B(n_232),
.Y(n_2956)
);

NAND2xp33_ASAP7_75t_SL g2957 ( 
.A(n_2832),
.B(n_232),
.Y(n_2957)
);

INVx3_ASAP7_75t_L g2958 ( 
.A(n_2801),
.Y(n_2958)
);

CKINVDCx20_ASAP7_75t_R g2959 ( 
.A(n_2834),
.Y(n_2959)
);

CKINVDCx5p33_ASAP7_75t_R g2960 ( 
.A(n_2838),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2784),
.B(n_233),
.Y(n_2961)
);

NAND2xp33_ASAP7_75t_R g2962 ( 
.A(n_2840),
.B(n_2841),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2786),
.B(n_233),
.Y(n_2963)
);

NAND2xp33_ASAP7_75t_SL g2964 ( 
.A(n_2844),
.B(n_234),
.Y(n_2964)
);

OR2x2_ASAP7_75t_L g2965 ( 
.A(n_2780),
.B(n_234),
.Y(n_2965)
);

AND2x4_ASAP7_75t_L g2966 ( 
.A(n_2769),
.B(n_235),
.Y(n_2966)
);

AO221x2_ASAP7_75t_L g2967 ( 
.A1(n_2850),
.A2(n_238),
.B1(n_241),
.B2(n_237),
.C(n_240),
.Y(n_2967)
);

INVx4_ASAP7_75t_L g2968 ( 
.A(n_2783),
.Y(n_2968)
);

OAI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2816),
.A2(n_240),
.B1(n_236),
.B2(n_238),
.Y(n_2969)
);

INVx2_ASAP7_75t_SL g2970 ( 
.A(n_2852),
.Y(n_2970)
);

NAND2xp33_ASAP7_75t_SL g2971 ( 
.A(n_2853),
.B(n_236),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2772),
.B(n_241),
.Y(n_2972)
);

A2O1A1Ixp33_ASAP7_75t_L g2973 ( 
.A1(n_2858),
.A2(n_252),
.B(n_260),
.C(n_242),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2788),
.B(n_242),
.Y(n_2974)
);

AND2x4_ASAP7_75t_L g2975 ( 
.A(n_2754),
.B(n_243),
.Y(n_2975)
);

AO221x2_ASAP7_75t_L g2976 ( 
.A1(n_2851),
.A2(n_247),
.B1(n_249),
.B2(n_246),
.C(n_248),
.Y(n_2976)
);

NOR4xp25_ASAP7_75t_SL g2977 ( 
.A(n_2790),
.B(n_247),
.C(n_243),
.D(n_246),
.Y(n_2977)
);

AO221x2_ASAP7_75t_L g2978 ( 
.A1(n_2851),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.C(n_253),
.Y(n_2978)
);

NOR2xp67_ASAP7_75t_L g2979 ( 
.A(n_2754),
.B(n_250),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2788),
.B(n_253),
.Y(n_2980)
);

AO221x2_ASAP7_75t_L g2981 ( 
.A1(n_2851),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.C(n_257),
.Y(n_2981)
);

AND2x2_ASAP7_75t_L g2982 ( 
.A(n_2789),
.B(n_254),
.Y(n_2982)
);

AO221x2_ASAP7_75t_L g2983 ( 
.A1(n_2851),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.C(n_259),
.Y(n_2983)
);

CKINVDCx5p33_ASAP7_75t_R g2984 ( 
.A(n_2798),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2788),
.B(n_258),
.Y(n_2985)
);

AND2x2_ASAP7_75t_L g2986 ( 
.A(n_2789),
.B(n_260),
.Y(n_2986)
);

AO221x2_ASAP7_75t_L g2987 ( 
.A1(n_2851),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.C(n_265),
.Y(n_2987)
);

AOI22xp5_ASAP7_75t_L g2988 ( 
.A1(n_2759),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_2988)
);

AND2x2_ASAP7_75t_L g2989 ( 
.A(n_2789),
.B(n_265),
.Y(n_2989)
);

OAI22xp33_ASAP7_75t_L g2990 ( 
.A1(n_2851),
.A2(n_269),
.B1(n_266),
.B2(n_268),
.Y(n_2990)
);

OR2x2_ASAP7_75t_L g2991 ( 
.A(n_2761),
.B(n_266),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2788),
.B(n_268),
.Y(n_2992)
);

AO221x2_ASAP7_75t_L g2993 ( 
.A1(n_2851),
.A2(n_274),
.B1(n_276),
.B2(n_272),
.C(n_275),
.Y(n_2993)
);

AO221x2_ASAP7_75t_L g2994 ( 
.A1(n_2851),
.A2(n_274),
.B1(n_276),
.B2(n_272),
.C(n_275),
.Y(n_2994)
);

OAI221xp5_ASAP7_75t_L g2995 ( 
.A1(n_2851),
.A2(n_278),
.B1(n_271),
.B2(n_277),
.C(n_279),
.Y(n_2995)
);

AND2x4_ASAP7_75t_SL g2996 ( 
.A(n_2754),
.B(n_271),
.Y(n_2996)
);

NOR2xp67_ASAP7_75t_L g2997 ( 
.A(n_2754),
.B(n_277),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2788),
.B(n_278),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2788),
.B(n_279),
.Y(n_2999)
);

OAI221xp5_ASAP7_75t_L g3000 ( 
.A1(n_2851),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.C(n_283),
.Y(n_3000)
);

OAI22xp33_ASAP7_75t_L g3001 ( 
.A1(n_2851),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_3001)
);

INVx3_ASAP7_75t_L g3002 ( 
.A(n_2854),
.Y(n_3002)
);

OR2x2_ASAP7_75t_L g3003 ( 
.A(n_2761),
.B(n_283),
.Y(n_3003)
);

NOR4xp25_ASAP7_75t_SL g3004 ( 
.A(n_2790),
.B(n_286),
.C(n_284),
.D(n_285),
.Y(n_3004)
);

OAI221xp5_ASAP7_75t_L g3005 ( 
.A1(n_2851),
.A2(n_287),
.B1(n_284),
.B2(n_286),
.C(n_289),
.Y(n_3005)
);

NOR2xp33_ASAP7_75t_L g3006 ( 
.A(n_2785),
.B(n_287),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2881),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2899),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2908),
.B(n_290),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2930),
.B(n_290),
.Y(n_3010)
);

BUFx3_ASAP7_75t_L g3011 ( 
.A(n_2865),
.Y(n_3011)
);

NOR2x1_ASAP7_75t_L g3012 ( 
.A(n_2979),
.B(n_291),
.Y(n_3012)
);

INVxp67_ASAP7_75t_L g3013 ( 
.A(n_2905),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2929),
.B(n_292),
.Y(n_3014)
);

INVx1_ASAP7_75t_SL g3015 ( 
.A(n_2889),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2883),
.B(n_292),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2871),
.Y(n_3017)
);

AND2x2_ASAP7_75t_L g3018 ( 
.A(n_3002),
.B(n_2958),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_SL g3019 ( 
.A(n_2997),
.B(n_293),
.Y(n_3019)
);

INVx1_ASAP7_75t_SL g3020 ( 
.A(n_2996),
.Y(n_3020)
);

INVx1_ASAP7_75t_SL g3021 ( 
.A(n_2984),
.Y(n_3021)
);

HB1xp67_ASAP7_75t_L g3022 ( 
.A(n_2894),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2890),
.Y(n_3023)
);

BUFx2_ASAP7_75t_L g3024 ( 
.A(n_2877),
.Y(n_3024)
);

NOR2xp33_ASAP7_75t_L g3025 ( 
.A(n_2944),
.B(n_294),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2925),
.Y(n_3026)
);

AOI22xp33_ASAP7_75t_L g3027 ( 
.A1(n_2879),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2910),
.B(n_297),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2924),
.Y(n_3029)
);

BUFx2_ASAP7_75t_L g3030 ( 
.A(n_2938),
.Y(n_3030)
);

HB1xp67_ASAP7_75t_L g3031 ( 
.A(n_2945),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2940),
.Y(n_3032)
);

OR2x2_ASAP7_75t_L g3033 ( 
.A(n_2939),
.B(n_298),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2970),
.B(n_298),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2942),
.Y(n_3035)
);

OAI22xp5_ASAP7_75t_L g3036 ( 
.A1(n_2911),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2968),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2863),
.B(n_299),
.Y(n_3038)
);

BUFx3_ASAP7_75t_L g3039 ( 
.A(n_2933),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_2873),
.B(n_2982),
.Y(n_3040)
);

OR2x2_ASAP7_75t_L g3041 ( 
.A(n_2876),
.B(n_300),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2974),
.B(n_302),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2943),
.Y(n_3043)
);

HB1xp67_ASAP7_75t_L g3044 ( 
.A(n_2991),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2946),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2986),
.B(n_303),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_3003),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2989),
.B(n_303),
.Y(n_3048)
);

INVx1_ASAP7_75t_SL g3049 ( 
.A(n_2921),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2892),
.B(n_304),
.Y(n_3050)
);

NOR2xp33_ASAP7_75t_L g3051 ( 
.A(n_2965),
.B(n_2947),
.Y(n_3051)
);

AND2x4_ASAP7_75t_SL g3052 ( 
.A(n_2860),
.B(n_305),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2956),
.B(n_305),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2980),
.Y(n_3054)
);

OAI22xp5_ASAP7_75t_L g3055 ( 
.A1(n_2995),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2985),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2992),
.Y(n_3057)
);

HB1xp67_ASAP7_75t_L g3058 ( 
.A(n_2948),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2998),
.B(n_2999),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2922),
.Y(n_3060)
);

OAI21x1_ASAP7_75t_L g3061 ( 
.A1(n_2880),
.A2(n_306),
.B(n_307),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2932),
.Y(n_3062)
);

CKINVDCx16_ASAP7_75t_R g3063 ( 
.A(n_2874),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2917),
.B(n_308),
.Y(n_3064)
);

AOI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_2879),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2887),
.B(n_311),
.Y(n_3066)
);

OR2x2_ASAP7_75t_L g3067 ( 
.A(n_2897),
.B(n_312),
.Y(n_3067)
);

AOI22xp33_ASAP7_75t_SL g3068 ( 
.A1(n_2978),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_3068)
);

INVx4_ASAP7_75t_L g3069 ( 
.A(n_2975),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2891),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2896),
.B(n_313),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2898),
.B(n_314),
.Y(n_3072)
);

INVx1_ASAP7_75t_SL g3073 ( 
.A(n_2913),
.Y(n_3073)
);

AO21x2_ASAP7_75t_L g3074 ( 
.A1(n_2901),
.A2(n_315),
.B(n_316),
.Y(n_3074)
);

BUFx2_ASAP7_75t_L g3075 ( 
.A(n_2882),
.Y(n_3075)
);

HB1xp67_ASAP7_75t_L g3076 ( 
.A(n_2888),
.Y(n_3076)
);

AND2x2_ASAP7_75t_L g3077 ( 
.A(n_2915),
.B(n_315),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2904),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2909),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2934),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2926),
.Y(n_3081)
);

NOR2xp33_ASAP7_75t_L g3082 ( 
.A(n_2912),
.B(n_316),
.Y(n_3082)
);

OAI22xp5_ASAP7_75t_L g3083 ( 
.A1(n_3000),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_3083)
);

HB1xp67_ASAP7_75t_L g3084 ( 
.A(n_2962),
.Y(n_3084)
);

OAI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_3005),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_3085)
);

INVx2_ASAP7_75t_SL g3086 ( 
.A(n_2966),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2961),
.Y(n_3087)
);

AOI22xp33_ASAP7_75t_L g3088 ( 
.A1(n_2978),
.A2(n_2983),
.B1(n_2987),
.B2(n_2981),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2952),
.B(n_320),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2950),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2963),
.Y(n_3091)
);

CKINVDCx16_ASAP7_75t_R g3092 ( 
.A(n_2868),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2935),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_L g3094 ( 
.A(n_3006),
.B(n_320),
.Y(n_3094)
);

BUFx6f_ASAP7_75t_L g3095 ( 
.A(n_2955),
.Y(n_3095)
);

INVx3_ASAP7_75t_L g3096 ( 
.A(n_2953),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2959),
.Y(n_3097)
);

NAND2x1_ASAP7_75t_SL g3098 ( 
.A(n_2884),
.B(n_2885),
.Y(n_3098)
);

AND2x4_ASAP7_75t_L g3099 ( 
.A(n_2960),
.B(n_321),
.Y(n_3099)
);

AND2x2_ASAP7_75t_L g3100 ( 
.A(n_2949),
.B(n_321),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2900),
.B(n_322),
.Y(n_3101)
);

INVx1_ASAP7_75t_SL g3102 ( 
.A(n_2931),
.Y(n_3102)
);

INVxp67_ASAP7_75t_L g3103 ( 
.A(n_2957),
.Y(n_3103)
);

AOI22xp5_ASAP7_75t_L g3104 ( 
.A1(n_2981),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_3104)
);

INVx1_ASAP7_75t_SL g3105 ( 
.A(n_2964),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2900),
.B(n_2903),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_2972),
.B(n_323),
.Y(n_3107)
);

AND2x2_ASAP7_75t_L g3108 ( 
.A(n_2941),
.B(n_326),
.Y(n_3108)
);

AOI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_2983),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_3109)
);

NOR2xp33_ASAP7_75t_L g3110 ( 
.A(n_2914),
.B(n_2951),
.Y(n_3110)
);

OAI22xp5_ASAP7_75t_L g3111 ( 
.A1(n_2919),
.A2(n_3001),
.B1(n_2990),
.B2(n_2988),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2903),
.B(n_327),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_2927),
.B(n_2967),
.Y(n_3113)
);

NOR2xp33_ASAP7_75t_L g3114 ( 
.A(n_2902),
.B(n_328),
.Y(n_3114)
);

AOI22xp5_ASAP7_75t_L g3115 ( 
.A1(n_2987),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_3115)
);

INVx6_ASAP7_75t_L g3116 ( 
.A(n_2971),
.Y(n_3116)
);

INVx4_ASAP7_75t_L g3117 ( 
.A(n_2886),
.Y(n_3117)
);

INVx3_ASAP7_75t_L g3118 ( 
.A(n_2895),
.Y(n_3118)
);

AND2x2_ASAP7_75t_L g3119 ( 
.A(n_2878),
.B(n_330),
.Y(n_3119)
);

INVx1_ASAP7_75t_SL g3120 ( 
.A(n_2861),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2907),
.Y(n_3121)
);

AOI22xp33_ASAP7_75t_L g3122 ( 
.A1(n_2862),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2906),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2920),
.Y(n_3124)
);

NOR2x1_ASAP7_75t_L g3125 ( 
.A(n_2969),
.B(n_332),
.Y(n_3125)
);

AOI22xp33_ASAP7_75t_L g3126 ( 
.A1(n_2976),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_3126)
);

AND2x2_ASAP7_75t_L g3127 ( 
.A(n_2923),
.B(n_334),
.Y(n_3127)
);

CKINVDCx16_ASAP7_75t_R g3128 ( 
.A(n_2864),
.Y(n_3128)
);

AND2x2_ASAP7_75t_L g3129 ( 
.A(n_2918),
.B(n_335),
.Y(n_3129)
);

OR2x2_ASAP7_75t_L g3130 ( 
.A(n_2993),
.B(n_336),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_2866),
.B(n_336),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2936),
.Y(n_3132)
);

INVx4_ASAP7_75t_L g3133 ( 
.A(n_2867),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_2994),
.B(n_337),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_2973),
.B(n_337),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2937),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2893),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2916),
.Y(n_3138)
);

HB1xp67_ASAP7_75t_L g3139 ( 
.A(n_2928),
.Y(n_3139)
);

AND2x4_ASAP7_75t_L g3140 ( 
.A(n_2869),
.B(n_338),
.Y(n_3140)
);

INVxp67_ASAP7_75t_L g3141 ( 
.A(n_2872),
.Y(n_3141)
);

OAI221xp5_ASAP7_75t_L g3142 ( 
.A1(n_2875),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.C(n_341),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2977),
.Y(n_3143)
);

OR2x2_ASAP7_75t_L g3144 ( 
.A(n_2954),
.B(n_340),
.Y(n_3144)
);

INVx2_ASAP7_75t_SL g3145 ( 
.A(n_3004),
.Y(n_3145)
);

AND2x4_ASAP7_75t_L g3146 ( 
.A(n_2870),
.B(n_341),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2881),
.Y(n_3147)
);

AND2x2_ASAP7_75t_L g3148 ( 
.A(n_2908),
.B(n_343),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_2908),
.B(n_344),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_2908),
.B(n_344),
.Y(n_3150)
);

INVxp67_ASAP7_75t_L g3151 ( 
.A(n_2905),
.Y(n_3151)
);

OR2x2_ASAP7_75t_L g3152 ( 
.A(n_2908),
.B(n_346),
.Y(n_3152)
);

OAI22xp5_ASAP7_75t_L g3153 ( 
.A1(n_2908),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2899),
.Y(n_3154)
);

INVx2_ASAP7_75t_SL g3155 ( 
.A(n_2889),
.Y(n_3155)
);

OR2x2_ASAP7_75t_L g3156 ( 
.A(n_2908),
.B(n_348),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2870),
.B(n_349),
.Y(n_3157)
);

OR2x2_ASAP7_75t_L g3158 ( 
.A(n_2908),
.B(n_349),
.Y(n_3158)
);

AND2x4_ASAP7_75t_L g3159 ( 
.A(n_2938),
.B(n_351),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_2908),
.B(n_350),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2899),
.Y(n_3161)
);

INVxp67_ASAP7_75t_L g3162 ( 
.A(n_2905),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2870),
.B(n_351),
.Y(n_3163)
);

INVx1_ASAP7_75t_SL g3164 ( 
.A(n_2908),
.Y(n_3164)
);

OR2x2_ASAP7_75t_L g3165 ( 
.A(n_2908),
.B(n_352),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2899),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2881),
.Y(n_3167)
);

INVx2_ASAP7_75t_SL g3168 ( 
.A(n_2889),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2870),
.B(n_352),
.Y(n_3169)
);

NAND2xp33_ASAP7_75t_SL g3170 ( 
.A(n_2874),
.B(n_353),
.Y(n_3170)
);

AND3x2_ASAP7_75t_L g3171 ( 
.A(n_2892),
.B(n_353),
.C(n_354),
.Y(n_3171)
);

HB1xp67_ASAP7_75t_L g3172 ( 
.A(n_2883),
.Y(n_3172)
);

AOI22xp33_ASAP7_75t_L g3173 ( 
.A1(n_2879),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_3173)
);

INVx1_ASAP7_75t_SL g3174 ( 
.A(n_2908),
.Y(n_3174)
);

NOR2x1_ASAP7_75t_L g3175 ( 
.A(n_2979),
.B(n_357),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2881),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2899),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2881),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2870),
.B(n_358),
.Y(n_3179)
);

INVx1_ASAP7_75t_SL g3180 ( 
.A(n_2908),
.Y(n_3180)
);

BUFx2_ASAP7_75t_L g3181 ( 
.A(n_2908),
.Y(n_3181)
);

INVxp67_ASAP7_75t_L g3182 ( 
.A(n_2905),
.Y(n_3182)
);

OR2x2_ASAP7_75t_L g3183 ( 
.A(n_2908),
.B(n_358),
.Y(n_3183)
);

INVx1_ASAP7_75t_SL g3184 ( 
.A(n_2908),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2899),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_2908),
.B(n_359),
.Y(n_3186)
);

AOI222xp33_ASAP7_75t_L g3187 ( 
.A1(n_2995),
.A2(n_362),
.B1(n_364),
.B2(n_360),
.C1(n_361),
.C2(n_363),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_2881),
.Y(n_3188)
);

HB1xp67_ASAP7_75t_L g3189 ( 
.A(n_2883),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2881),
.Y(n_3190)
);

BUFx3_ASAP7_75t_L g3191 ( 
.A(n_2865),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2881),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_2944),
.B(n_360),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2899),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2870),
.B(n_363),
.Y(n_3195)
);

AND2x4_ASAP7_75t_L g3196 ( 
.A(n_2870),
.B(n_365),
.Y(n_3196)
);

OAI22xp5_ASAP7_75t_L g3197 ( 
.A1(n_2908),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2870),
.B(n_367),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2870),
.B(n_368),
.Y(n_3199)
);

OR2x2_ASAP7_75t_L g3200 ( 
.A(n_2908),
.B(n_369),
.Y(n_3200)
);

HB1xp67_ASAP7_75t_L g3201 ( 
.A(n_2883),
.Y(n_3201)
);

OR2x2_ASAP7_75t_L g3202 ( 
.A(n_2908),
.B(n_369),
.Y(n_3202)
);

OR2x2_ASAP7_75t_L g3203 ( 
.A(n_2908),
.B(n_370),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2899),
.Y(n_3204)
);

INVx1_ASAP7_75t_SL g3205 ( 
.A(n_2908),
.Y(n_3205)
);

BUFx3_ASAP7_75t_L g3206 ( 
.A(n_2865),
.Y(n_3206)
);

OAI22xp5_ASAP7_75t_L g3207 ( 
.A1(n_2908),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2899),
.Y(n_3208)
);

INVx3_ASAP7_75t_L g3209 ( 
.A(n_2968),
.Y(n_3209)
);

OR2x2_ASAP7_75t_L g3210 ( 
.A(n_2908),
.B(n_371),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2881),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3008),
.Y(n_3212)
);

AOI22xp5_ASAP7_75t_L g3213 ( 
.A1(n_3110),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_3213)
);

OR2x2_ASAP7_75t_L g3214 ( 
.A(n_3084),
.B(n_374),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3154),
.Y(n_3215)
);

AND2x2_ASAP7_75t_L g3216 ( 
.A(n_3181),
.B(n_375),
.Y(n_3216)
);

NAND2xp33_ASAP7_75t_L g3217 ( 
.A(n_3076),
.B(n_376),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_3161),
.Y(n_3218)
);

AOI322xp5_ASAP7_75t_L g3219 ( 
.A1(n_3088),
.A2(n_381),
.A3(n_380),
.B1(n_378),
.B2(n_376),
.C1(n_377),
.C2(n_379),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3166),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3177),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_3093),
.B(n_3132),
.Y(n_3222)
);

INVxp67_ASAP7_75t_L g3223 ( 
.A(n_3058),
.Y(n_3223)
);

INVx1_ASAP7_75t_SL g3224 ( 
.A(n_3170),
.Y(n_3224)
);

AOI22xp5_ASAP7_75t_L g3225 ( 
.A1(n_3092),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_3225)
);

AND2x4_ASAP7_75t_L g3226 ( 
.A(n_3164),
.B(n_3174),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_3045),
.B(n_380),
.Y(n_3227)
);

A2O1A1Ixp33_ASAP7_75t_SL g3228 ( 
.A1(n_3114),
.A2(n_383),
.B(n_381),
.C(n_382),
.Y(n_3228)
);

OR2x2_ASAP7_75t_L g3229 ( 
.A(n_3172),
.B(n_384),
.Y(n_3229)
);

OAI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_3063),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_3230)
);

AND2x2_ASAP7_75t_L g3231 ( 
.A(n_3180),
.B(n_386),
.Y(n_3231)
);

INVx1_ASAP7_75t_SL g3232 ( 
.A(n_3049),
.Y(n_3232)
);

AOI21xp33_ASAP7_75t_SL g3233 ( 
.A1(n_3128),
.A2(n_387),
.B(n_388),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3044),
.B(n_389),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3185),
.Y(n_3235)
);

OAI21xp33_ASAP7_75t_L g3236 ( 
.A1(n_3068),
.A2(n_390),
.B(n_391),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3194),
.Y(n_3237)
);

AOI21xp33_ASAP7_75t_L g3238 ( 
.A1(n_3111),
.A2(n_391),
.B(n_392),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_3184),
.B(n_392),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3204),
.Y(n_3240)
);

OAI33xp33_ASAP7_75t_L g3241 ( 
.A1(n_3106),
.A2(n_3101),
.A3(n_3112),
.B1(n_3137),
.B2(n_3121),
.B3(n_3124),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3205),
.B(n_393),
.Y(n_3242)
);

INVx2_ASAP7_75t_L g3243 ( 
.A(n_3209),
.Y(n_3243)
);

NOR3xp33_ASAP7_75t_L g3244 ( 
.A(n_3055),
.B(n_393),
.C(n_394),
.Y(n_3244)
);

INVxp33_ASAP7_75t_L g3245 ( 
.A(n_3098),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3208),
.Y(n_3246)
);

OAI22xp5_ASAP7_75t_L g3247 ( 
.A1(n_3117),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3013),
.A2(n_395),
.B(n_396),
.Y(n_3248)
);

NOR3xp33_ASAP7_75t_L g3249 ( 
.A(n_3083),
.B(n_399),
.C(n_400),
.Y(n_3249)
);

O2A1O1Ixp33_ASAP7_75t_L g3250 ( 
.A1(n_3139),
.A2(n_403),
.B(n_401),
.C(n_402),
.Y(n_3250)
);

OAI221xp5_ASAP7_75t_L g3251 ( 
.A1(n_3151),
.A2(n_405),
.B1(n_401),
.B2(n_404),
.C(n_406),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3087),
.B(n_404),
.Y(n_3252)
);

OAI22xp5_ASAP7_75t_L g3253 ( 
.A1(n_3118),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_3075),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3091),
.B(n_408),
.Y(n_3255)
);

NOR2x1_ASAP7_75t_L g3256 ( 
.A(n_3152),
.B(n_409),
.Y(n_3256)
);

OAI22xp33_ASAP7_75t_L g3257 ( 
.A1(n_3104),
.A2(n_3115),
.B1(n_3133),
.B2(n_3162),
.Y(n_3257)
);

NOR2xp33_ASAP7_75t_L g3258 ( 
.A(n_3182),
.B(n_409),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3022),
.Y(n_3259)
);

OAI21xp33_ASAP7_75t_L g3260 ( 
.A1(n_3109),
.A2(n_410),
.B(n_411),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3029),
.Y(n_3261)
);

AOI222xp33_ASAP7_75t_L g3262 ( 
.A1(n_3141),
.A2(n_412),
.B1(n_414),
.B2(n_410),
.C1(n_411),
.C2(n_413),
.Y(n_3262)
);

OAI332xp33_ASAP7_75t_L g3263 ( 
.A1(n_3130),
.A2(n_419),
.A3(n_418),
.B1(n_416),
.B2(n_420),
.B3(n_412),
.C1(n_415),
.C2(n_417),
.Y(n_3263)
);

OR2x2_ASAP7_75t_L g3264 ( 
.A(n_3189),
.B(n_415),
.Y(n_3264)
);

BUFx3_ASAP7_75t_L g3265 ( 
.A(n_3011),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3136),
.B(n_418),
.Y(n_3266)
);

OR2x2_ASAP7_75t_L g3267 ( 
.A(n_3201),
.B(n_419),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_3018),
.B(n_420),
.Y(n_3268)
);

OAI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_3027),
.A2(n_3173),
.B1(n_3065),
.B2(n_3126),
.Y(n_3269)
);

AOI22xp5_ASAP7_75t_L g3270 ( 
.A1(n_3113),
.A2(n_424),
.B1(n_421),
.B2(n_422),
.Y(n_3270)
);

OAI22xp33_ASAP7_75t_SL g3271 ( 
.A1(n_3116),
.A2(n_424),
.B1(n_421),
.B2(n_422),
.Y(n_3271)
);

AND2x2_ASAP7_75t_L g3272 ( 
.A(n_3024),
.B(n_425),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3047),
.Y(n_3273)
);

OAI322xp33_ASAP7_75t_L g3274 ( 
.A1(n_3123),
.A2(n_431),
.A3(n_430),
.B1(n_427),
.B2(n_425),
.C1(n_426),
.C2(n_428),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3030),
.Y(n_3275)
);

OAI32xp33_ASAP7_75t_L g3276 ( 
.A1(n_3120),
.A2(n_432),
.A3(n_426),
.B1(n_428),
.B2(n_433),
.Y(n_3276)
);

INVx1_ASAP7_75t_SL g3277 ( 
.A(n_3021),
.Y(n_3277)
);

OAI21xp5_ASAP7_75t_SL g3278 ( 
.A1(n_3187),
.A2(n_432),
.B(n_433),
.Y(n_3278)
);

AND2x2_ASAP7_75t_L g3279 ( 
.A(n_3037),
.B(n_434),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_3081),
.B(n_434),
.Y(n_3280)
);

INVxp67_ASAP7_75t_L g3281 ( 
.A(n_3156),
.Y(n_3281)
);

OR2x2_ASAP7_75t_L g3282 ( 
.A(n_3031),
.B(n_435),
.Y(n_3282)
);

INVxp67_ASAP7_75t_L g3283 ( 
.A(n_3158),
.Y(n_3283)
);

OAI222xp33_ASAP7_75t_L g3284 ( 
.A1(n_3125),
.A2(n_438),
.B1(n_440),
.B2(n_436),
.C1(n_437),
.C2(n_439),
.Y(n_3284)
);

OAI22xp33_ASAP7_75t_L g3285 ( 
.A1(n_3019),
.A2(n_438),
.B1(n_436),
.B2(n_437),
.Y(n_3285)
);

OAI21xp33_ASAP7_75t_L g3286 ( 
.A1(n_3122),
.A2(n_439),
.B(n_440),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3039),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_SL g3288 ( 
.A(n_3012),
.B(n_441),
.Y(n_3288)
);

O2A1O1Ixp33_ASAP7_75t_L g3289 ( 
.A1(n_3138),
.A2(n_444),
.B(n_441),
.C(n_443),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3116),
.Y(n_3290)
);

AOI22xp33_ASAP7_75t_L g3291 ( 
.A1(n_3085),
.A2(n_447),
.B1(n_445),
.B2(n_446),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3032),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3054),
.B(n_445),
.Y(n_3293)
);

HB1xp67_ASAP7_75t_L g3294 ( 
.A(n_3159),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3035),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_3056),
.B(n_3057),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3069),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3142),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3080),
.B(n_3028),
.Y(n_3299)
);

AOI22xp5_ASAP7_75t_L g3300 ( 
.A1(n_3131),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_3062),
.B(n_449),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3078),
.B(n_452),
.Y(n_3302)
);

AOI211xp5_ASAP7_75t_L g3303 ( 
.A1(n_3036),
.A2(n_454),
.B(n_452),
.C(n_453),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3079),
.B(n_454),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_3102),
.A2(n_455),
.B(n_456),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3043),
.Y(n_3306)
);

AOI322xp5_ASAP7_75t_L g3307 ( 
.A1(n_3134),
.A2(n_461),
.A3(n_460),
.B1(n_458),
.B2(n_456),
.C1(n_457),
.C2(n_459),
.Y(n_3307)
);

OAI32xp33_ASAP7_75t_L g3308 ( 
.A1(n_3105),
.A2(n_461),
.A3(n_457),
.B1(n_459),
.B2(n_462),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3159),
.B(n_462),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3060),
.Y(n_3310)
);

INVxp67_ASAP7_75t_SL g3311 ( 
.A(n_3103),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3010),
.B(n_463),
.Y(n_3312)
);

AOI221xp5_ASAP7_75t_L g3313 ( 
.A1(n_3153),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.C(n_466),
.Y(n_3313)
);

OAI22xp5_ASAP7_75t_SL g3314 ( 
.A1(n_3175),
.A2(n_466),
.B1(n_464),
.B2(n_465),
.Y(n_3314)
);

OAI31xp33_ASAP7_75t_L g3315 ( 
.A1(n_3197),
.A2(n_469),
.A3(n_467),
.B(n_468),
.Y(n_3315)
);

AOI222xp33_ASAP7_75t_L g3316 ( 
.A1(n_3127),
.A2(n_470),
.B1(n_472),
.B2(n_467),
.C1(n_469),
.C2(n_471),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_SL g3317 ( 
.A(n_3155),
.B(n_470),
.Y(n_3317)
);

AOI31xp33_ASAP7_75t_L g3318 ( 
.A1(n_3145),
.A2(n_3183),
.A3(n_3200),
.B(n_3165),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3017),
.Y(n_3319)
);

INVxp67_ASAP7_75t_L g3320 ( 
.A(n_3202),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3097),
.B(n_472),
.Y(n_3321)
);

AOI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3207),
.A2(n_477),
.B1(n_474),
.B2(n_475),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3095),
.B(n_474),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3007),
.Y(n_3324)
);

OR2x2_ASAP7_75t_L g3325 ( 
.A(n_3023),
.B(n_477),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3026),
.Y(n_3326)
);

INVxp67_ASAP7_75t_SL g3327 ( 
.A(n_3203),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3147),
.Y(n_3328)
);

AND2x4_ASAP7_75t_L g3329 ( 
.A(n_3168),
.B(n_478),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3095),
.B(n_3040),
.Y(n_3330)
);

INVxp67_ASAP7_75t_L g3331 ( 
.A(n_3210),
.Y(n_3331)
);

AOI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_3140),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_3332)
);

NOR2xp67_ASAP7_75t_L g3333 ( 
.A(n_3096),
.B(n_479),
.Y(n_3333)
);

AOI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_3143),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3167),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_3070),
.B(n_481),
.Y(n_3336)
);

AOI21xp33_ASAP7_75t_L g3337 ( 
.A1(n_3082),
.A2(n_482),
.B(n_484),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3135),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.Y(n_3338)
);

AOI22xp33_ASAP7_75t_L g3339 ( 
.A1(n_3094),
.A2(n_488),
.B1(n_485),
.B2(n_487),
.Y(n_3339)
);

OR2x2_ASAP7_75t_L g3340 ( 
.A(n_3176),
.B(n_3178),
.Y(n_3340)
);

AOI22xp33_ASAP7_75t_SL g3341 ( 
.A1(n_3009),
.A2(n_490),
.B1(n_487),
.B2(n_489),
.Y(n_3341)
);

AOI22xp33_ASAP7_75t_SL g3342 ( 
.A1(n_3148),
.A2(n_491),
.B1(n_489),
.B2(n_490),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_3149),
.B(n_491),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_3015),
.B(n_492),
.Y(n_3344)
);

OAI21xp5_ASAP7_75t_L g3345 ( 
.A1(n_3129),
.A2(n_493),
.B(n_494),
.Y(n_3345)
);

XNOR2xp5_ASAP7_75t_L g3346 ( 
.A(n_3150),
.B(n_493),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3160),
.B(n_494),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3074),
.B(n_495),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3188),
.Y(n_3349)
);

OAI22xp33_ASAP7_75t_L g3350 ( 
.A1(n_3144),
.A2(n_497),
.B1(n_495),
.B2(n_496),
.Y(n_3350)
);

AOI22xp5_ASAP7_75t_L g3351 ( 
.A1(n_3186),
.A2(n_500),
.B1(n_496),
.B2(n_498),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3190),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3192),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3211),
.Y(n_3354)
);

INVx1_ASAP7_75t_SL g3355 ( 
.A(n_3191),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_3086),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_3051),
.B(n_498),
.Y(n_3357)
);

OAI222xp33_ASAP7_75t_L g3358 ( 
.A1(n_3157),
.A2(n_504),
.B1(n_506),
.B2(n_502),
.C1(n_503),
.C2(n_505),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_SL g3359 ( 
.A(n_3206),
.B(n_502),
.Y(n_3359)
);

OR2x2_ASAP7_75t_L g3360 ( 
.A(n_3327),
.B(n_3059),
.Y(n_3360)
);

INVxp67_ASAP7_75t_L g3361 ( 
.A(n_3294),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_3226),
.B(n_3073),
.Y(n_3362)
);

NAND2xp33_ASAP7_75t_L g3363 ( 
.A(n_3224),
.B(n_3020),
.Y(n_3363)
);

OR2x2_ASAP7_75t_L g3364 ( 
.A(n_3275),
.B(n_3199),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3261),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3226),
.B(n_3090),
.Y(n_3366)
);

NOR2xp33_ASAP7_75t_L g3367 ( 
.A(n_3241),
.B(n_3067),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3290),
.B(n_3107),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3311),
.B(n_3171),
.Y(n_3369)
);

INVx1_ASAP7_75t_SL g3370 ( 
.A(n_3277),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3265),
.Y(n_3371)
);

NOR2x1_ASAP7_75t_L g3372 ( 
.A(n_3333),
.B(n_3016),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3257),
.B(n_3119),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3254),
.B(n_3100),
.Y(n_3374)
);

AND2x4_ASAP7_75t_L g3375 ( 
.A(n_3287),
.B(n_3146),
.Y(n_3375)
);

OR2x2_ASAP7_75t_L g3376 ( 
.A(n_3281),
.B(n_3163),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3212),
.Y(n_3377)
);

OR2x2_ASAP7_75t_L g3378 ( 
.A(n_3283),
.B(n_3198),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3215),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_L g3380 ( 
.A(n_3232),
.B(n_3025),
.Y(n_3380)
);

AND2x2_ASAP7_75t_L g3381 ( 
.A(n_3330),
.B(n_3034),
.Y(n_3381)
);

OR2x2_ASAP7_75t_L g3382 ( 
.A(n_3320),
.B(n_3169),
.Y(n_3382)
);

HB1xp67_ASAP7_75t_L g3383 ( 
.A(n_3331),
.Y(n_3383)
);

AND2x2_ASAP7_75t_L g3384 ( 
.A(n_3297),
.B(n_3196),
.Y(n_3384)
);

INVxp67_ASAP7_75t_L g3385 ( 
.A(n_3288),
.Y(n_3385)
);

OAI22xp5_ASAP7_75t_L g3386 ( 
.A1(n_3245),
.A2(n_3195),
.B1(n_3179),
.B2(n_3193),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3318),
.B(n_3053),
.Y(n_3387)
);

OAI31xp33_ASAP7_75t_SL g3388 ( 
.A1(n_3269),
.A2(n_3061),
.A3(n_3108),
.B(n_3089),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3223),
.B(n_3050),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_L g3390 ( 
.A(n_3355),
.B(n_3038),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3356),
.B(n_3046),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3218),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3220),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3259),
.B(n_3048),
.Y(n_3394)
);

NAND2xp33_ASAP7_75t_L g3395 ( 
.A(n_3256),
.B(n_3071),
.Y(n_3395)
);

HB1xp67_ASAP7_75t_L g3396 ( 
.A(n_3214),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3216),
.B(n_3042),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3243),
.B(n_3099),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3221),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_3231),
.B(n_3077),
.Y(n_3400)
);

NOR2xp33_ASAP7_75t_L g3401 ( 
.A(n_3299),
.B(n_3066),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3235),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3237),
.Y(n_3403)
);

AND2x2_ASAP7_75t_L g3404 ( 
.A(n_3239),
.B(n_3052),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_3325),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3240),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3334),
.B(n_3072),
.Y(n_3407)
);

INVxp67_ASAP7_75t_SL g3408 ( 
.A(n_3217),
.Y(n_3408)
);

INVxp67_ASAP7_75t_L g3409 ( 
.A(n_3258),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3271),
.B(n_3064),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3242),
.B(n_3033),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3280),
.B(n_3014),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3233),
.B(n_3041),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3246),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3324),
.Y(n_3415)
);

AND2x4_ASAP7_75t_L g3416 ( 
.A(n_3329),
.B(n_503),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3225),
.B(n_3301),
.Y(n_3417)
);

AO22x2_ASAP7_75t_L g3418 ( 
.A1(n_3222),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3326),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3305),
.B(n_507),
.Y(n_3420)
);

OR2x2_ASAP7_75t_L g3421 ( 
.A(n_3340),
.B(n_507),
.Y(n_3421)
);

NOR2xp67_ASAP7_75t_L g3422 ( 
.A(n_3282),
.B(n_508),
.Y(n_3422)
);

AOI22xp33_ASAP7_75t_R g3423 ( 
.A1(n_3263),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.Y(n_3423)
);

AND2x4_ASAP7_75t_L g3424 ( 
.A(n_3273),
.B(n_511),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3272),
.B(n_512),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3328),
.Y(n_3426)
);

OR2x2_ASAP7_75t_L g3427 ( 
.A(n_3296),
.B(n_513),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3335),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3270),
.B(n_513),
.Y(n_3429)
);

INVx2_ASAP7_75t_SL g3430 ( 
.A(n_3329),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_3227),
.B(n_514),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3268),
.B(n_514),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3349),
.Y(n_3433)
);

AOI22xp5_ASAP7_75t_L g3434 ( 
.A1(n_3278),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_3279),
.B(n_516),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3343),
.B(n_518),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3300),
.B(n_518),
.Y(n_3437)
);

NOR2xp33_ASAP7_75t_L g3438 ( 
.A(n_3252),
.B(n_519),
.Y(n_3438)
);

AND2x2_ASAP7_75t_L g3439 ( 
.A(n_3347),
.B(n_520),
.Y(n_3439)
);

NOR2xp33_ASAP7_75t_L g3440 ( 
.A(n_3255),
.B(n_520),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3292),
.B(n_521),
.Y(n_3441)
);

NOR2xp33_ASAP7_75t_L g3442 ( 
.A(n_3293),
.B(n_521),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3352),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_SL g3444 ( 
.A(n_3285),
.B(n_522),
.Y(n_3444)
);

INVx1_ASAP7_75t_SL g3445 ( 
.A(n_3229),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3295),
.B(n_522),
.Y(n_3446)
);

NAND2xp33_ASAP7_75t_L g3447 ( 
.A(n_3236),
.B(n_523),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3336),
.B(n_524),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3306),
.B(n_524),
.Y(n_3449)
);

NAND2x1_ASAP7_75t_L g3450 ( 
.A(n_3354),
.B(n_525),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3353),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_SL g3452 ( 
.A(n_3341),
.B(n_525),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3310),
.B(n_526),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3319),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3234),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3321),
.B(n_526),
.Y(n_3456)
);

HB1xp67_ASAP7_75t_L g3457 ( 
.A(n_3264),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3267),
.Y(n_3458)
);

CKINVDCx5p33_ASAP7_75t_R g3459 ( 
.A(n_3370),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3383),
.Y(n_3460)
);

BUFx2_ASAP7_75t_L g3461 ( 
.A(n_3372),
.Y(n_3461)
);

INVx1_ASAP7_75t_SL g3462 ( 
.A(n_3404),
.Y(n_3462)
);

HB1xp67_ASAP7_75t_L g3463 ( 
.A(n_3430),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3396),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3366),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_3398),
.B(n_3344),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3361),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_3375),
.Y(n_3468)
);

INVx2_ASAP7_75t_L g3469 ( 
.A(n_3371),
.Y(n_3469)
);

INVx1_ASAP7_75t_SL g3470 ( 
.A(n_3362),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3457),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3421),
.Y(n_3472)
);

BUFx2_ASAP7_75t_L g3473 ( 
.A(n_3385),
.Y(n_3473)
);

BUFx4f_ASAP7_75t_SL g3474 ( 
.A(n_3416),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3405),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3411),
.B(n_3248),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3458),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3377),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3379),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3392),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3393),
.Y(n_3481)
);

CKINVDCx5p33_ASAP7_75t_R g3482 ( 
.A(n_3380),
.Y(n_3482)
);

BUFx2_ASAP7_75t_L g3483 ( 
.A(n_3408),
.Y(n_3483)
);

INVxp67_ASAP7_75t_L g3484 ( 
.A(n_3395),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3399),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3402),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3403),
.Y(n_3487)
);

INVx5_ASAP7_75t_L g3488 ( 
.A(n_3424),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3406),
.Y(n_3489)
);

INVxp33_ASAP7_75t_SL g3490 ( 
.A(n_3369),
.Y(n_3490)
);

INVxp33_ASAP7_75t_SL g3491 ( 
.A(n_3390),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3414),
.Y(n_3492)
);

INVxp33_ASAP7_75t_L g3493 ( 
.A(n_3400),
.Y(n_3493)
);

NOR2xp33_ASAP7_75t_R g3494 ( 
.A(n_3363),
.B(n_3346),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3365),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3415),
.Y(n_3496)
);

NOR2xp33_ASAP7_75t_L g3497 ( 
.A(n_3413),
.B(n_3302),
.Y(n_3497)
);

INVxp67_ASAP7_75t_L g3498 ( 
.A(n_3422),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3419),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3426),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3367),
.B(n_3230),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3428),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3433),
.Y(n_3503)
);

NOR2xp33_ASAP7_75t_L g3504 ( 
.A(n_3409),
.B(n_3410),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3443),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3451),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3384),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3424),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3381),
.B(n_3304),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3454),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3360),
.Y(n_3511)
);

HB1xp67_ASAP7_75t_L g3512 ( 
.A(n_3445),
.Y(n_3512)
);

HB1xp67_ASAP7_75t_L g3513 ( 
.A(n_3450),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3394),
.Y(n_3514)
);

BUFx2_ASAP7_75t_L g3515 ( 
.A(n_3374),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_L g3516 ( 
.A(n_3387),
.B(n_3266),
.Y(n_3516)
);

BUFx6f_ASAP7_75t_L g3517 ( 
.A(n_3435),
.Y(n_3517)
);

NAND2x1_ASAP7_75t_SL g3518 ( 
.A(n_3368),
.B(n_3351),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3388),
.B(n_3348),
.Y(n_3519)
);

INVx1_ASAP7_75t_SL g3520 ( 
.A(n_3436),
.Y(n_3520)
);

HB1xp67_ASAP7_75t_L g3521 ( 
.A(n_3389),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3441),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3446),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3449),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_3391),
.Y(n_3525)
);

NOR2xp33_ASAP7_75t_L g3526 ( 
.A(n_3397),
.B(n_3357),
.Y(n_3526)
);

BUFx6f_ASAP7_75t_SL g3527 ( 
.A(n_3455),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3364),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3453),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3376),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3378),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3448),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3382),
.Y(n_3533)
);

INVxp33_ASAP7_75t_SL g3534 ( 
.A(n_3386),
.Y(n_3534)
);

NOR2xp33_ASAP7_75t_L g3535 ( 
.A(n_3417),
.B(n_3312),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3418),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3418),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3427),
.Y(n_3538)
);

INVx1_ASAP7_75t_SL g3539 ( 
.A(n_3439),
.Y(n_3539)
);

INVxp33_ASAP7_75t_SL g3540 ( 
.A(n_3434),
.Y(n_3540)
);

INVx2_ASAP7_75t_L g3541 ( 
.A(n_3432),
.Y(n_3541)
);

XNOR2x2_ASAP7_75t_L g3542 ( 
.A(n_3452),
.B(n_3247),
.Y(n_3542)
);

INVx1_ASAP7_75t_SL g3543 ( 
.A(n_3456),
.Y(n_3543)
);

NOR2xp33_ASAP7_75t_L g3544 ( 
.A(n_3373),
.B(n_3309),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3412),
.Y(n_3545)
);

HB1xp67_ASAP7_75t_L g3546 ( 
.A(n_3425),
.Y(n_3546)
);

HB1xp67_ASAP7_75t_L g3547 ( 
.A(n_3444),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3431),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3420),
.Y(n_3549)
);

INVx5_ASAP7_75t_SL g3550 ( 
.A(n_3423),
.Y(n_3550)
);

INVx3_ASAP7_75t_L g3551 ( 
.A(n_3407),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3437),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3438),
.Y(n_3553)
);

INVx2_ASAP7_75t_SL g3554 ( 
.A(n_3429),
.Y(n_3554)
);

INVx8_ASAP7_75t_L g3555 ( 
.A(n_3440),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3442),
.Y(n_3556)
);

NOR2xp33_ASAP7_75t_L g3557 ( 
.A(n_3401),
.B(n_3317),
.Y(n_3557)
);

INVx2_ASAP7_75t_SL g3558 ( 
.A(n_3447),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3370),
.B(n_3307),
.Y(n_3559)
);

NOR2x1_ASAP7_75t_L g3560 ( 
.A(n_3372),
.B(n_3284),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3383),
.Y(n_3561)
);

NAND2x1_ASAP7_75t_SL g3562 ( 
.A(n_3372),
.B(n_3338),
.Y(n_3562)
);

NOR2x1_ASAP7_75t_L g3563 ( 
.A(n_3560),
.B(n_3250),
.Y(n_3563)
);

NAND3xp33_ASAP7_75t_SL g3564 ( 
.A(n_3494),
.B(n_3303),
.C(n_3316),
.Y(n_3564)
);

NOR2x1_ASAP7_75t_L g3565 ( 
.A(n_3461),
.B(n_3358),
.Y(n_3565)
);

NOR4xp25_ASAP7_75t_L g3566 ( 
.A(n_3501),
.B(n_3289),
.C(n_3238),
.D(n_3274),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3550),
.B(n_3262),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3512),
.Y(n_3568)
);

AOI221xp5_ASAP7_75t_L g3569 ( 
.A1(n_3536),
.A2(n_3253),
.B1(n_3350),
.B2(n_3314),
.C(n_3337),
.Y(n_3569)
);

NOR2xp33_ASAP7_75t_L g3570 ( 
.A(n_3491),
.B(n_3323),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3550),
.B(n_3342),
.Y(n_3571)
);

NOR3x1_ASAP7_75t_L g3572 ( 
.A(n_3473),
.B(n_3251),
.C(n_3345),
.Y(n_3572)
);

AOI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_3540),
.A2(n_3244),
.B1(n_3249),
.B2(n_3260),
.Y(n_3573)
);

NAND3xp33_ASAP7_75t_SL g3574 ( 
.A(n_3470),
.B(n_3219),
.C(n_3315),
.Y(n_3574)
);

NOR3xp33_ASAP7_75t_SL g3575 ( 
.A(n_3482),
.B(n_3308),
.C(n_3276),
.Y(n_3575)
);

NOR3x1_ASAP7_75t_SL g3576 ( 
.A(n_3463),
.B(n_3213),
.C(n_3359),
.Y(n_3576)
);

NAND3x2_ASAP7_75t_L g3577 ( 
.A(n_3483),
.B(n_3228),
.C(n_3286),
.Y(n_3577)
);

OAI322xp33_ASAP7_75t_L g3578 ( 
.A1(n_3537),
.A2(n_3322),
.A3(n_3313),
.B1(n_3298),
.B2(n_3339),
.C1(n_3332),
.C2(n_3291),
.Y(n_3578)
);

AOI211xp5_ASAP7_75t_L g3579 ( 
.A1(n_3519),
.A2(n_530),
.B(n_528),
.C(n_529),
.Y(n_3579)
);

OAI211xp5_ASAP7_75t_L g3580 ( 
.A1(n_3518),
.A2(n_3562),
.B(n_3484),
.C(n_3547),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3459),
.B(n_3498),
.Y(n_3581)
);

AOI22xp5_ASAP7_75t_L g3582 ( 
.A1(n_3534),
.A2(n_530),
.B1(n_528),
.B2(n_529),
.Y(n_3582)
);

NOR2xp33_ASAP7_75t_SL g3583 ( 
.A(n_3474),
.B(n_3490),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3488),
.B(n_531),
.Y(n_3584)
);

NOR2x1_ASAP7_75t_L g3585 ( 
.A(n_3460),
.B(n_531),
.Y(n_3585)
);

OAI21xp33_ASAP7_75t_SL g3586 ( 
.A1(n_3513),
.A2(n_532),
.B(n_533),
.Y(n_3586)
);

NAND2x1_ASAP7_75t_SL g3587 ( 
.A(n_3466),
.B(n_532),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3561),
.Y(n_3588)
);

OAI21xp5_ASAP7_75t_SL g3589 ( 
.A1(n_3557),
.A2(n_534),
.B(n_535),
.Y(n_3589)
);

NOR4xp25_ASAP7_75t_L g3590 ( 
.A(n_3559),
.B(n_3504),
.C(n_3551),
.D(n_3554),
.Y(n_3590)
);

AOI22xp5_ASAP7_75t_L g3591 ( 
.A1(n_3558),
.A2(n_3527),
.B1(n_3497),
.B2(n_3462),
.Y(n_3591)
);

NAND4xp75_ASAP7_75t_L g3592 ( 
.A(n_3464),
.B(n_536),
.C(n_534),
.D(n_535),
.Y(n_3592)
);

NOR2x1p5_ASAP7_75t_L g3593 ( 
.A(n_3465),
.B(n_536),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3471),
.Y(n_3594)
);

NAND4xp25_ASAP7_75t_SL g3595 ( 
.A(n_3542),
.B(n_539),
.C(n_537),
.D(n_538),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_SL g3596 ( 
.A(n_3488),
.B(n_537),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3488),
.B(n_539),
.Y(n_3597)
);

OAI221xp5_ASAP7_75t_L g3598 ( 
.A1(n_3516),
.A2(n_3544),
.B1(n_3535),
.B2(n_3552),
.C(n_3476),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_SL g3599 ( 
.A(n_3517),
.B(n_540),
.Y(n_3599)
);

AOI21xp33_ASAP7_75t_L g3600 ( 
.A1(n_3493),
.A2(n_3543),
.B(n_3539),
.Y(n_3600)
);

NOR2xp33_ASAP7_75t_L g3601 ( 
.A(n_3517),
.B(n_540),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3515),
.B(n_541),
.Y(n_3602)
);

NOR2x1_ASAP7_75t_L g3603 ( 
.A(n_3467),
.B(n_3469),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_3555),
.A2(n_542),
.B(n_543),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3472),
.Y(n_3605)
);

NOR2xp33_ASAP7_75t_L g3606 ( 
.A(n_3520),
.B(n_542),
.Y(n_3606)
);

NAND5xp2_ASAP7_75t_L g3607 ( 
.A(n_3511),
.B(n_545),
.C(n_543),
.D(n_544),
.E(n_546),
.Y(n_3607)
);

OR3x1_ASAP7_75t_L g3608 ( 
.A(n_3508),
.B(n_544),
.C(n_545),
.Y(n_3608)
);

OAI21xp5_ASAP7_75t_SL g3609 ( 
.A1(n_3530),
.A2(n_546),
.B(n_547),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_SL g3610 ( 
.A(n_3468),
.B(n_547),
.Y(n_3610)
);

NAND2xp33_ASAP7_75t_L g3611 ( 
.A(n_3555),
.B(n_548),
.Y(n_3611)
);

NOR4xp25_ASAP7_75t_L g3612 ( 
.A(n_3549),
.B(n_550),
.C(n_548),
.D(n_549),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3507),
.B(n_549),
.Y(n_3613)
);

NOR2xp67_ASAP7_75t_L g3614 ( 
.A(n_3528),
.B(n_3531),
.Y(n_3614)
);

OAI21xp33_ASAP7_75t_SL g3615 ( 
.A1(n_3533),
.A2(n_550),
.B(n_551),
.Y(n_3615)
);

INVxp67_ASAP7_75t_L g3616 ( 
.A(n_3521),
.Y(n_3616)
);

NOR2x1_ASAP7_75t_L g3617 ( 
.A(n_3553),
.B(n_552),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3541),
.B(n_553),
.Y(n_3618)
);

NOR3xp33_ASAP7_75t_L g3619 ( 
.A(n_3538),
.B(n_3523),
.C(n_3522),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3532),
.B(n_554),
.Y(n_3620)
);

NOR3xp33_ASAP7_75t_SL g3621 ( 
.A(n_3475),
.B(n_554),
.C(n_555),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3477),
.Y(n_3622)
);

AND4x1_ASAP7_75t_L g3623 ( 
.A(n_3526),
.B(n_557),
.C(n_555),
.D(n_556),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3546),
.Y(n_3624)
);

OAI21x1_ASAP7_75t_L g3625 ( 
.A1(n_3478),
.A2(n_556),
.B(n_557),
.Y(n_3625)
);

NAND3xp33_ASAP7_75t_L g3626 ( 
.A(n_3514),
.B(n_558),
.C(n_559),
.Y(n_3626)
);

O2A1O1Ixp5_ASAP7_75t_L g3627 ( 
.A1(n_3525),
.A2(n_560),
.B(n_558),
.C(n_559),
.Y(n_3627)
);

NOR2xp67_ASAP7_75t_L g3628 ( 
.A(n_3556),
.B(n_560),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_SL g3629 ( 
.A(n_3509),
.B(n_561),
.Y(n_3629)
);

OAI221xp5_ASAP7_75t_L g3630 ( 
.A1(n_3548),
.A2(n_568),
.B1(n_564),
.B2(n_567),
.C(n_570),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_3545),
.A2(n_567),
.B(n_568),
.Y(n_3631)
);

NAND3xp33_ASAP7_75t_L g3632 ( 
.A(n_3524),
.B(n_571),
.C(n_572),
.Y(n_3632)
);

AOI21x1_ASAP7_75t_L g3633 ( 
.A1(n_3596),
.A2(n_3496),
.B(n_3495),
.Y(n_3633)
);

AOI221xp5_ASAP7_75t_L g3634 ( 
.A1(n_3590),
.A2(n_3481),
.B1(n_3485),
.B2(n_3480),
.C(n_3479),
.Y(n_3634)
);

NAND3x1_ASAP7_75t_SL g3635 ( 
.A(n_3563),
.B(n_3529),
.C(n_3500),
.Y(n_3635)
);

O2A1O1Ixp33_ASAP7_75t_L g3636 ( 
.A1(n_3580),
.A2(n_3487),
.B(n_3489),
.C(n_3486),
.Y(n_3636)
);

AOI211xp5_ASAP7_75t_L g3637 ( 
.A1(n_3595),
.A2(n_3499),
.B(n_3503),
.C(n_3502),
.Y(n_3637)
);

OAI221xp5_ASAP7_75t_SL g3638 ( 
.A1(n_3566),
.A2(n_3510),
.B1(n_3492),
.B2(n_3506),
.C(n_3505),
.Y(n_3638)
);

OAI211xp5_ASAP7_75t_SL g3639 ( 
.A1(n_3565),
.A2(n_573),
.B(n_571),
.C(n_572),
.Y(n_3639)
);

AOI211xp5_ASAP7_75t_SL g3640 ( 
.A1(n_3600),
.A2(n_576),
.B(n_574),
.C(n_575),
.Y(n_3640)
);

AOI221xp5_ASAP7_75t_L g3641 ( 
.A1(n_3567),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.C(n_577),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3587),
.Y(n_3642)
);

O2A1O1Ixp33_ASAP7_75t_L g3643 ( 
.A1(n_3571),
.A2(n_581),
.B(n_578),
.C(n_580),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3568),
.Y(n_3644)
);

AOI22xp5_ASAP7_75t_L g3645 ( 
.A1(n_3574),
.A2(n_583),
.B1(n_578),
.B2(n_582),
.Y(n_3645)
);

AND2x4_ASAP7_75t_L g3646 ( 
.A(n_3614),
.B(n_582),
.Y(n_3646)
);

HB1xp67_ASAP7_75t_L g3647 ( 
.A(n_3628),
.Y(n_3647)
);

AOI211xp5_ASAP7_75t_L g3648 ( 
.A1(n_3564),
.A2(n_585),
.B(n_583),
.C(n_584),
.Y(n_3648)
);

NAND4xp75_ASAP7_75t_L g3649 ( 
.A(n_3603),
.B(n_589),
.C(n_587),
.D(n_588),
.Y(n_3649)
);

OAI321xp33_ASAP7_75t_L g3650 ( 
.A1(n_3576),
.A2(n_590),
.A3(n_592),
.B1(n_588),
.B2(n_589),
.C(n_591),
.Y(n_3650)
);

AOI21xp5_ASAP7_75t_L g3651 ( 
.A1(n_3583),
.A2(n_593),
.B(n_595),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3612),
.B(n_593),
.Y(n_3652)
);

AOI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3569),
.A2(n_597),
.B1(n_595),
.B2(n_596),
.Y(n_3653)
);

OAI211xp5_ASAP7_75t_L g3654 ( 
.A1(n_3577),
.A2(n_600),
.B(n_598),
.C(n_599),
.Y(n_3654)
);

NAND3xp33_ASAP7_75t_L g3655 ( 
.A(n_3591),
.B(n_600),
.C(n_601),
.Y(n_3655)
);

OAI221xp5_ASAP7_75t_L g3656 ( 
.A1(n_3573),
.A2(n_603),
.B1(n_601),
.B2(n_602),
.C(n_605),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3570),
.B(n_602),
.Y(n_3657)
);

OAI221xp5_ASAP7_75t_L g3658 ( 
.A1(n_3598),
.A2(n_3575),
.B1(n_3581),
.B2(n_3579),
.C(n_3616),
.Y(n_3658)
);

AOI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3608),
.A2(n_607),
.B1(n_605),
.B2(n_606),
.Y(n_3659)
);

OAI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3582),
.A2(n_610),
.B1(n_608),
.B2(n_609),
.Y(n_3660)
);

AOI211xp5_ASAP7_75t_SL g3661 ( 
.A1(n_3594),
.A2(n_610),
.B(n_608),
.C(n_609),
.Y(n_3661)
);

AOI211xp5_ASAP7_75t_L g3662 ( 
.A1(n_3578),
.A2(n_613),
.B(n_611),
.C(n_612),
.Y(n_3662)
);

HB1xp67_ASAP7_75t_L g3663 ( 
.A(n_3585),
.Y(n_3663)
);

AOI221xp5_ASAP7_75t_L g3664 ( 
.A1(n_3588),
.A2(n_614),
.B1(n_611),
.B2(n_612),
.C(n_615),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3584),
.Y(n_3665)
);

INVx1_ASAP7_75t_SL g3666 ( 
.A(n_3611),
.Y(n_3666)
);

OAI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3586),
.A2(n_614),
.B(n_615),
.Y(n_3667)
);

AOI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_3597),
.A2(n_616),
.B(n_617),
.Y(n_3668)
);

AOI211xp5_ASAP7_75t_L g3669 ( 
.A1(n_3589),
.A2(n_619),
.B(n_617),
.C(n_618),
.Y(n_3669)
);

OAI321xp33_ASAP7_75t_L g3670 ( 
.A1(n_3624),
.A2(n_619),
.A3(n_620),
.B1(n_621),
.B2(n_622),
.C(n_623),
.Y(n_3670)
);

NOR2x1_ASAP7_75t_SL g3671 ( 
.A(n_3599),
.B(n_620),
.Y(n_3671)
);

INVx1_ASAP7_75t_SL g3672 ( 
.A(n_3617),
.Y(n_3672)
);

OAI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_3627),
.A2(n_621),
.B(n_622),
.Y(n_3673)
);

NOR4xp25_ASAP7_75t_L g3674 ( 
.A(n_3605),
.B(n_3622),
.C(n_3609),
.D(n_3615),
.Y(n_3674)
);

HB1xp67_ASAP7_75t_L g3675 ( 
.A(n_3593),
.Y(n_3675)
);

OAI211xp5_ASAP7_75t_SL g3676 ( 
.A1(n_3619),
.A2(n_625),
.B(n_623),
.C(n_624),
.Y(n_3676)
);

AOI22xp5_ASAP7_75t_L g3677 ( 
.A1(n_3606),
.A2(n_626),
.B1(n_624),
.B2(n_625),
.Y(n_3677)
);

OAI22xp5_ASAP7_75t_L g3678 ( 
.A1(n_3621),
.A2(n_628),
.B1(n_626),
.B2(n_627),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3604),
.B(n_627),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3618),
.Y(n_3680)
);

AO22x2_ASAP7_75t_L g3681 ( 
.A1(n_3602),
.A2(n_633),
.B1(n_629),
.B2(n_631),
.Y(n_3681)
);

OAI22xp5_ASAP7_75t_L g3682 ( 
.A1(n_3626),
.A2(n_635),
.B1(n_633),
.B2(n_634),
.Y(n_3682)
);

AOI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_3631),
.A2(n_634),
.B(n_635),
.Y(n_3683)
);

NOR2xp33_ASAP7_75t_L g3684 ( 
.A(n_3629),
.B(n_636),
.Y(n_3684)
);

OAI21xp5_ASAP7_75t_SL g3685 ( 
.A1(n_3632),
.A2(n_3623),
.B(n_3613),
.Y(n_3685)
);

OAI21xp5_ASAP7_75t_SL g3686 ( 
.A1(n_3601),
.A2(n_636),
.B(n_637),
.Y(n_3686)
);

INVx2_ASAP7_75t_SL g3687 ( 
.A(n_3625),
.Y(n_3687)
);

AO22x2_ASAP7_75t_L g3688 ( 
.A1(n_3592),
.A2(n_639),
.B1(n_637),
.B2(n_638),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3620),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3647),
.Y(n_3690)
);

AOI22xp5_ASAP7_75t_L g3691 ( 
.A1(n_3639),
.A2(n_3610),
.B1(n_3630),
.B2(n_3572),
.Y(n_3691)
);

OR2x2_ASAP7_75t_L g3692 ( 
.A(n_3672),
.B(n_3607),
.Y(n_3692)
);

AOI22xp5_ASAP7_75t_L g3693 ( 
.A1(n_3653),
.A2(n_641),
.B1(n_638),
.B2(n_640),
.Y(n_3693)
);

NAND4xp25_ASAP7_75t_L g3694 ( 
.A(n_3658),
.B(n_642),
.C(n_640),
.D(n_641),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3663),
.Y(n_3695)
);

NOR2x1_ASAP7_75t_L g3696 ( 
.A(n_3649),
.B(n_3646),
.Y(n_3696)
);

NOR2x1p5_ASAP7_75t_L g3697 ( 
.A(n_3642),
.B(n_3655),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3675),
.Y(n_3698)
);

NOR2xp67_ASAP7_75t_L g3699 ( 
.A(n_3650),
.B(n_642),
.Y(n_3699)
);

XOR2x1_ASAP7_75t_L g3700 ( 
.A(n_3646),
.B(n_643),
.Y(n_3700)
);

OAI211xp5_ASAP7_75t_L g3701 ( 
.A1(n_3662),
.A2(n_3674),
.B(n_3645),
.C(n_3634),
.Y(n_3701)
);

AND2x4_ASAP7_75t_L g3702 ( 
.A(n_3687),
.B(n_643),
.Y(n_3702)
);

INVxp33_ASAP7_75t_L g3703 ( 
.A(n_3671),
.Y(n_3703)
);

XOR2xp5_ASAP7_75t_L g3704 ( 
.A(n_3659),
.B(n_644),
.Y(n_3704)
);

NAND4xp75_ASAP7_75t_L g3705 ( 
.A(n_3644),
.B(n_646),
.C(n_644),
.D(n_645),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3680),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3657),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3666),
.B(n_645),
.Y(n_3708)
);

AOI22xp5_ASAP7_75t_L g3709 ( 
.A1(n_3654),
.A2(n_648),
.B1(n_646),
.B2(n_647),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_3667),
.B(n_3665),
.Y(n_3710)
);

AND2x2_ASAP7_75t_L g3711 ( 
.A(n_3689),
.B(n_649),
.Y(n_3711)
);

AOI22xp5_ASAP7_75t_L g3712 ( 
.A1(n_3685),
.A2(n_652),
.B1(n_649),
.B2(n_650),
.Y(n_3712)
);

NOR2x1_ASAP7_75t_L g3713 ( 
.A(n_3686),
.B(n_652),
.Y(n_3713)
);

OR2x2_ASAP7_75t_L g3714 ( 
.A(n_3673),
.B(n_653),
.Y(n_3714)
);

NOR2x1_ASAP7_75t_L g3715 ( 
.A(n_3652),
.B(n_653),
.Y(n_3715)
);

AOI22xp5_ASAP7_75t_L g3716 ( 
.A1(n_3648),
.A2(n_657),
.B1(n_654),
.B2(n_655),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3633),
.Y(n_3717)
);

NAND5xp2_ASAP7_75t_L g3718 ( 
.A(n_3636),
.B(n_657),
.C(n_654),
.D(n_655),
.E(n_658),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3681),
.Y(n_3719)
);

NOR2x1p5_ASAP7_75t_L g3720 ( 
.A(n_3679),
.B(n_659),
.Y(n_3720)
);

INVx1_ASAP7_75t_SL g3721 ( 
.A(n_3688),
.Y(n_3721)
);

NAND2xp33_ASAP7_75t_SL g3722 ( 
.A(n_3703),
.B(n_3678),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_R g3723 ( 
.A(n_3690),
.B(n_3684),
.Y(n_3723)
);

NOR2xp33_ASAP7_75t_SL g3724 ( 
.A(n_3696),
.B(n_3638),
.Y(n_3724)
);

NAND2xp33_ASAP7_75t_SL g3725 ( 
.A(n_3692),
.B(n_3682),
.Y(n_3725)
);

NAND3xp33_ASAP7_75t_L g3726 ( 
.A(n_3701),
.B(n_3637),
.C(n_3640),
.Y(n_3726)
);

NAND2xp33_ASAP7_75t_SL g3727 ( 
.A(n_3717),
.B(n_3635),
.Y(n_3727)
);

NOR2xp33_ASAP7_75t_R g3728 ( 
.A(n_3698),
.B(n_3661),
.Y(n_3728)
);

NAND3xp33_ASAP7_75t_SL g3729 ( 
.A(n_3721),
.B(n_3643),
.C(n_3669),
.Y(n_3729)
);

NOR2xp33_ASAP7_75t_R g3730 ( 
.A(n_3695),
.B(n_3688),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3700),
.B(n_3651),
.Y(n_3731)
);

NOR2xp33_ASAP7_75t_R g3732 ( 
.A(n_3719),
.B(n_3707),
.Y(n_3732)
);

NAND2xp33_ASAP7_75t_L g3733 ( 
.A(n_3713),
.B(n_3681),
.Y(n_3733)
);

XNOR2x1_ASAP7_75t_L g3734 ( 
.A(n_3697),
.B(n_3660),
.Y(n_3734)
);

NOR2xp33_ASAP7_75t_R g3735 ( 
.A(n_3706),
.B(n_3670),
.Y(n_3735)
);

NOR2xp33_ASAP7_75t_R g3736 ( 
.A(n_3710),
.B(n_3668),
.Y(n_3736)
);

NOR2xp33_ASAP7_75t_R g3737 ( 
.A(n_3708),
.B(n_3676),
.Y(n_3737)
);

XNOR2x1_ASAP7_75t_L g3738 ( 
.A(n_3734),
.B(n_3715),
.Y(n_3738)
);

NAND4xp75_ASAP7_75t_L g3739 ( 
.A(n_3731),
.B(n_3699),
.C(n_3641),
.D(n_3711),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3733),
.Y(n_3740)
);

INVxp33_ASAP7_75t_L g3741 ( 
.A(n_3728),
.Y(n_3741)
);

AOI22xp5_ASAP7_75t_L g3742 ( 
.A1(n_3724),
.A2(n_3691),
.B1(n_3694),
.B2(n_3704),
.Y(n_3742)
);

AOI321xp33_ASAP7_75t_L g3743 ( 
.A1(n_3726),
.A2(n_3714),
.A3(n_3656),
.B1(n_3702),
.B2(n_3683),
.C(n_3716),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3740),
.Y(n_3744)
);

NAND2x1p5_ASAP7_75t_L g3745 ( 
.A(n_3738),
.B(n_3702),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3739),
.Y(n_3746)
);

NOR2xp67_ASAP7_75t_L g3747 ( 
.A(n_3744),
.B(n_3718),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3745),
.Y(n_3748)
);

OAI21x1_ASAP7_75t_L g3749 ( 
.A1(n_3746),
.A2(n_3720),
.B(n_3742),
.Y(n_3749)
);

AOI31xp33_ASAP7_75t_L g3750 ( 
.A1(n_3748),
.A2(n_3741),
.A3(n_3727),
.B(n_3722),
.Y(n_3750)
);

AOI31xp33_ASAP7_75t_L g3751 ( 
.A1(n_3747),
.A2(n_3725),
.A3(n_3729),
.B(n_3712),
.Y(n_3751)
);

AOI31xp33_ASAP7_75t_L g3752 ( 
.A1(n_3749),
.A2(n_3709),
.A3(n_3732),
.B(n_3730),
.Y(n_3752)
);

NAND5xp2_ASAP7_75t_L g3753 ( 
.A(n_3751),
.B(n_3743),
.C(n_3723),
.D(n_3735),
.E(n_3736),
.Y(n_3753)
);

OA22x2_ASAP7_75t_L g3754 ( 
.A1(n_3752),
.A2(n_3693),
.B1(n_3677),
.B2(n_3737),
.Y(n_3754)
);

XNOR2xp5_ASAP7_75t_L g3755 ( 
.A(n_3750),
.B(n_3705),
.Y(n_3755)
);

OAI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3754),
.A2(n_3664),
.B1(n_3753),
.B2(n_3755),
.Y(n_3756)
);

AOI221xp5_ASAP7_75t_L g3757 ( 
.A1(n_3753),
.A2(n_662),
.B1(n_660),
.B2(n_661),
.C(n_663),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3756),
.Y(n_3758)
);

AOI221xp5_ASAP7_75t_L g3759 ( 
.A1(n_3758),
.A2(n_3757),
.B1(n_664),
.B2(n_660),
.C(n_662),
.Y(n_3759)
);

AOI211xp5_ASAP7_75t_L g3760 ( 
.A1(n_3759),
.A2(n_667),
.B(n_665),
.C(n_666),
.Y(n_3760)
);


endmodule