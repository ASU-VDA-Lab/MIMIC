module fake_netlist_1_10200_n_21 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_21;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
CKINVDCx20_ASAP7_75t_R g8 ( .A(n_6), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_3), .B(n_2), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
INVx3_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
AOI22xp33_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_12), .B1(n_11), .B2(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
NOR2x1_ASAP7_75t_L g18 ( .A(n_17), .B(n_9), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_19), .B(n_1), .Y(n_20) );
XNOR2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_5), .Y(n_21) );
endmodule