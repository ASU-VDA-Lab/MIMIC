module fake_jpeg_13223_n_62 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

MAJIxp5_ASAP7_75t_L g11 ( 
.A(n_8),
.B(n_2),
.C(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

AND2x2_ASAP7_75t_SL g16 ( 
.A(n_6),
.B(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_12),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_17),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_15),
.Y(n_31)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_22),
.B(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_17),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_25),
.B1(n_10),
.B2(n_12),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_11),
.A2(n_18),
.B(n_1),
.C(n_3),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_24),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_14),
.B(n_18),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_33),
.B(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_15),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_9),
.B1(n_10),
.B2(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_22),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_19),
.B1(n_21),
.B2(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_42),
.Y(n_46)
);

AND2x4_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_21),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_43),
.B(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_8),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_30),
.B1(n_19),
.B2(n_41),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_47),
.B1(n_0),
.B2(n_4),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_27),
.C(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_49),
.A2(n_50),
.B1(n_46),
.B2(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_55),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_46),
.C(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_54),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_4),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_6),
.C(n_3),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_57),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_57),
.B(n_60),
.Y(n_62)
);


endmodule