module fake_jpeg_26257_n_67 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_67);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_67;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_38;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;
wire n_66;

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.Y(n_45)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_1),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_35),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_37),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_49),
.B(n_53),
.Y(n_55)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_51),
.B1(n_29),
.B2(n_7),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_32),
.Y(n_53)
);

OAI22x1_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_56),
.B1(n_57),
.B2(n_52),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_5),
.B(n_8),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_9),
.B(n_10),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_48),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_58),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_59),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

AOI321xp33_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_12),
.A3(n_13),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_65),
.A2(n_50),
.B1(n_25),
.B2(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_22),
.Y(n_67)
);


endmodule