module real_jpeg_29602_n_16 (n_338, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_338;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_0),
.A2(n_22),
.B1(n_23),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_0),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_0),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_46),
.Y(n_290)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_1),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_1),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_1),
.A2(n_135),
.B(n_149),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_2),
.A2(n_44),
.B1(n_57),
.B2(n_58),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_44),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_3),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_3),
.B(n_29),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_3),
.A2(n_29),
.B(n_161),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_118),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_3),
.A2(n_11),
.B(n_57),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_3),
.B(n_75),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_3),
.A2(n_97),
.B1(n_98),
.B2(n_212),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_115),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_115),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_115),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_8),
.A2(n_35),
.B1(n_51),
.B2(n_52),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_8),
.A2(n_35),
.B1(n_57),
.B2(n_58),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_24),
.B1(n_51),
.B2(n_52),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_9),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_9),
.A2(n_24),
.B1(n_57),
.B2(n_58),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_10),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_113),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_113),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_113),
.Y(n_204)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_12),
.A2(n_22),
.B1(n_23),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_12),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_120),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_12),
.A2(n_51),
.B1(n_52),
.B2(n_120),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_120),
.Y(n_212)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_14),
.A2(n_51),
.B1(n_52),
.B2(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_15),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_82),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_80),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_36),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_19),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_20),
.A2(n_42),
.B(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_21),
.A2(n_31),
.B(n_79),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_25),
.B(n_26),
.C(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_26),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_22),
.B(n_118),
.CON(n_117),
.SN(n_117)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_25),
.A2(n_31),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_26),
.B(n_29),
.Y(n_132)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_28),
.A2(n_29),
.B1(n_65),
.B2(n_66),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_28),
.A2(n_32),
.B1(n_117),
.B2(n_132),
.Y(n_131)
);

AOI32xp33_ASAP7_75t_L g160 ( 
.A1(n_28),
.A2(n_51),
.A3(n_64),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_30),
.A2(n_43),
.B(n_47),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_31),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_34),
.B(n_47),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_72),
.C(n_77),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_38),
.A2(n_39),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_48),
.C(n_61),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_40),
.A2(n_41),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_42),
.A2(n_47),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_42),
.A2(n_47),
.B1(n_126),
.B2(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_47),
.B(n_118),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_48),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_48),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_48),
.A2(n_61),
.B1(n_305),
.B2(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_56),
.B(n_59),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_49),
.A2(n_59),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_49),
.A2(n_56),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_49),
.A2(n_169),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_49),
.A2(n_56),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_49),
.A2(n_56),
.B1(n_168),
.B2(n_187),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_49),
.A2(n_56),
.B1(n_92),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_49),
.A2(n_108),
.B(n_245),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g162 ( 
.A(n_52),
.B(n_65),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_52),
.A2(n_55),
.B(n_118),
.C(n_189),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_56),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_56),
.B(n_118),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_58),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_60),
.B(n_109),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_61),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_62),
.A2(n_74),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_63),
.A2(n_70),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_63),
.A2(n_70),
.B1(n_112),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_63),
.A2(n_70),
.B1(n_145),
.B2(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_63),
.B(n_69),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_63),
.A2(n_70),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_68),
.A2(n_75),
.B(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_74),
.A2(n_76),
.B(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_74),
.A2(n_255),
.B(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_77),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_330),
.B(n_336),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_300),
.A3(n_322),
.B1(n_328),
.B2(n_329),
.C(n_338),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_281),
.B(n_299),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_259),
.B(n_280),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_150),
.B(n_235),
.C(n_258),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_137),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_88),
.B(n_137),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_121),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_105),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_90),
.B(n_105),
.C(n_121),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_91),
.B(n_96),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_93),
.B(n_179),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B(n_100),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_97),
.A2(n_99),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_97),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_97),
.A2(n_136),
.B1(n_204),
.B2(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_97),
.A2(n_136),
.B(n_276),
.Y(n_275)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_98),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_98),
.B(n_118),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_101),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_116),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_130),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_123),
.B(n_128),
.C(n_130),
.Y(n_256)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_133),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_143),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_138),
.A2(n_139),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_147),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_144),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_174),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_149),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_234),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_227),
.B(n_233),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_180),
.B(n_226),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_170),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_154),
.B(n_170),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_163),
.C(n_166),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_155),
.A2(n_156),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_160),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_158),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_159),
.A2(n_199),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_171),
.B(n_177),
.C(n_178),
.Y(n_228)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_220),
.B(n_225),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_200),
.B(n_219),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_183),
.B(n_190),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_208),
.B(n_218),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_202),
.B(n_206),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_213),
.B(n_217),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_228),
.B(n_229),
.Y(n_233)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_236),
.B(n_237),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_256),
.B2(n_257),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_247),
.C(n_257),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_250),
.C(n_254),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_261),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_279),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_272),
.B2(n_273),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_273),
.C(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_268),
.C(n_270),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_278),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_275),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_277),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_275),
.A2(n_293),
.B(n_296),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_283),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_297),
.B2(n_298),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_292),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_292),
.C(n_298),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B(n_291),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_290),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_302),
.C(n_312),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_291),
.A2(n_302),
.B1(n_303),
.B2(n_327),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_291),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_314),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_314),
.Y(n_329)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_307),
.C(n_309),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_309),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_311),
.B1(n_316),
.B2(n_320),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_320),
.C(n_321),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_313),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_321),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);


endmodule