module real_jpeg_4115_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_0),
.B(n_43),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_0),
.A2(n_42),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_0),
.B(n_135),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_0),
.B(n_270),
.C(n_273),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_0),
.A2(n_140),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_0),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_0),
.B(n_225),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_0),
.A2(n_46),
.B1(n_313),
.B2(n_321),
.Y(n_320)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_2),
.A2(n_56),
.B1(n_188),
.B2(n_191),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_3),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_3),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_3),
.A2(n_106),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_106),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_4),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_5),
.A2(n_114),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_5),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_132),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_5),
.A2(n_132),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_5),
.A2(n_132),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_6),
.A2(n_140),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_6),
.A2(n_47),
.B1(n_163),
.B2(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_6),
.A2(n_36),
.B1(n_163),
.B2(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_7),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_7),
.A2(n_69),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_8),
.Y(n_179)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_12),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_12),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_12),
.A2(n_44),
.B1(n_99),
.B2(n_231),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_12),
.A2(n_48),
.B1(n_99),
.B2(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_12),
.A2(n_99),
.B1(n_202),
.B2(n_353),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_13),
.Y(n_120)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_13),
.Y(n_123)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_13),
.Y(n_134)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_13),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_13),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_14),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_14),
.A2(n_113),
.B1(n_253),
.B2(n_256),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_14),
.A2(n_113),
.B1(n_202),
.B2(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_14),
.A2(n_113),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_15),
.Y(n_148)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_15),
.Y(n_151)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_15),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_236),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_235),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_193),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_20),
.B(n_193),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_137),
.C(n_174),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_21),
.B(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_73),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_22),
.B(n_74),
.C(n_110),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_45),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_23),
.B(n_45),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.A3(n_31),
.B1(n_34),
.B2(n_41),
.Y(n_23)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_27),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_27),
.Y(n_350)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_28),
.Y(n_255)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_33),
.A2(n_101),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVxp33_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_53),
.B1(n_61),
.B2(n_65),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_46),
.A2(n_65),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_46),
.B(n_181),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_46),
.A2(n_209),
.B(n_295),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_46),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_46),
.A2(n_178),
.B1(n_301),
.B2(n_313),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_46),
.A2(n_176),
.B(n_211),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_52),
.Y(n_247)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_52),
.Y(n_325)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_54),
.A2(n_208),
.B(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_58),
.Y(n_296)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_60),
.Y(n_217)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_60),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_68),
.Y(n_213)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_70),
.Y(n_302)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_71),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_110),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_94),
.B(n_102),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_75),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_75),
.A2(n_225),
.B1(n_252),
.B2(n_349),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_85),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_76),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_76),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_76),
.A2(n_171),
.B1(n_172),
.B2(n_251),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_76)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_77),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_77),
.Y(n_277)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_79),
.Y(n_344)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_81),
.Y(n_338)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_82),
.Y(n_201)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_83),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_83),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_83),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_92),
.Y(n_85)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI32xp33_ASAP7_75t_L g333 ( 
.A1(n_100),
.A2(n_334),
.A3(n_336),
.B1(n_339),
.B2(n_343),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_101),
.Y(n_228)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_101),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_103),
.A2(n_172),
.B(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_116),
.B1(n_130),
.B2(n_135),
.Y(n_110)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_117),
.A2(n_136),
.B1(n_165),
.B2(n_169),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_117),
.A2(n_131),
.B1(n_136),
.B2(n_230),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_127),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_128),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_137),
.B(n_174),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_164),
.C(n_170),
.Y(n_137)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_138),
.B(n_164),
.CI(n_170),
.CON(n_239),
.SN(n_239)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_144),
.B(n_158),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_139),
.B(n_192),
.Y(n_367)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_146)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_142),
.Y(n_345)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_186),
.B1(n_187),
.B2(n_192),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_144),
.A2(n_365),
.B(n_366),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_145),
.A2(n_159),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_145),
.A2(n_159),
.B1(n_275),
.B2(n_278),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_145),
.A2(n_159),
.B1(n_278),
.B2(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_145),
.A2(n_159),
.B1(n_287),
.B2(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_152),
.Y(n_145)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_147),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_149),
.B1(n_153),
.B2(n_156),
.Y(n_152)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_153),
.Y(n_273)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_185),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_175),
.B(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_179),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_188),
.Y(n_353)
);

INVx5_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_192),
.B(n_276),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_220),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_205),
.B2(n_206),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_218),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_217),
.Y(n_315)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_218),
.Y(n_321)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_234),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_229),
.B2(n_233),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_259),
.B(n_376),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_257),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_238),
.B(n_257),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_239),
.B(n_374),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_239),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_240),
.B(n_241),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.C(n_250),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_242),
.A2(n_243),
.B1(n_248),
.B2(n_249),
.Y(n_360)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_250),
.B(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_371),
.B(n_375),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_355),
.B(n_370),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_329),
.B(n_354),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_297),
.B(n_328),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_282),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_264),
.B(n_282),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_274),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_274),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_276),
.B(n_340),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_SL g349 ( 
.A1(n_276),
.A2(n_339),
.B(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_294),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_293),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_293),
.C(n_294),
.Y(n_330)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_286),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_309),
.B(n_327),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_308),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_308),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_302),
.B(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_319),
.B(n_326),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_311),
.B(n_312),
.Y(n_326)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_331),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_347),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_348),
.C(n_351),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_346),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_346),
.Y(n_363)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_352),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_356),
.B(n_357),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_361),
.B2(n_362),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_364),
.C(n_368),
.Y(n_372)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_368),
.B2(n_369),
.Y(n_362)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_363),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_364),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_373),
.Y(n_375)
);


endmodule