module fake_jpeg_13929_n_564 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_564);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_564;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_57),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_8),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_16),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_64),
.B(n_83),
.Y(n_161)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_21),
.B(n_8),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_28),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_82),
.Y(n_133)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_26),
.B(n_8),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_84),
.Y(n_175)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_86),
.Y(n_166)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_23),
.B(n_9),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_89),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_26),
.A2(n_9),
.B(n_15),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_90),
.Y(n_177)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_94),
.Y(n_163)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_18),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_102),
.Y(n_151)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_28),
.B(n_7),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_31),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_60),
.A2(n_37),
.B1(n_18),
.B2(n_47),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_111),
.A2(n_119),
.B(n_148),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_37),
.B1(n_29),
.B2(n_49),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_117),
.A2(n_124),
.B1(n_150),
.B2(n_152),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_47),
.B1(n_29),
.B2(n_20),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_65),
.A2(n_93),
.B1(n_106),
.B2(n_108),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_62),
.A2(n_29),
.B1(n_47),
.B2(n_49),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_138),
.B(n_27),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_142),
.B(n_155),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_69),
.A2(n_49),
.B1(n_50),
.B2(n_17),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_76),
.A2(n_17),
.B1(n_34),
.B2(n_50),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_74),
.A2(n_17),
.B1(n_34),
.B2(n_50),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_59),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_54),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_157),
.B(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_55),
.A2(n_53),
.B1(n_38),
.B2(n_41),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_174),
.B1(n_36),
.B2(n_33),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_54),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_78),
.B(n_40),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_169),
.B(n_38),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_57),
.A2(n_53),
.B1(n_42),
.B2(n_41),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_74),
.Y(n_201)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_180),
.Y(n_287)
);

AO22x1_ASAP7_75t_SL g182 ( 
.A1(n_117),
.A2(n_43),
.B1(n_48),
.B2(n_27),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_182),
.B(n_195),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_183),
.B(n_184),
.Y(n_254)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_185),
.Y(n_258)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_187),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_188),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_189),
.B(n_211),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_161),
.C(n_118),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_190),
.B(n_216),
.C(n_11),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_113),
.A2(n_34),
.B1(n_52),
.B2(n_95),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_192),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_193),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_120),
.B(n_42),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_121),
.Y(n_196)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_196),
.Y(n_303)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_197),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_198),
.A2(n_212),
.B1(n_213),
.B2(n_234),
.Y(n_260)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_200),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_201),
.Y(n_259)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_202),
.Y(n_295)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_203),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_SL g281 ( 
.A(n_204),
.B(n_220),
.Y(n_281)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_205),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_126),
.B(n_52),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_206),
.B(n_219),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_133),
.B(n_33),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_207),
.B(n_209),
.Y(n_257)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_208),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_39),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_177),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_164),
.A2(n_71),
.B1(n_66),
.B2(n_70),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_174),
.A2(n_92),
.B1(n_72),
.B2(n_58),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_144),
.Y(n_215)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_131),
.B(n_102),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_136),
.B(n_31),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_141),
.Y(n_221)
);

INVx11_ASAP7_75t_L g301 ( 
.A(n_221),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_132),
.B(n_40),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_237),
.Y(n_266)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_156),
.A2(n_98),
.B1(n_97),
.B2(n_96),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_225),
.A2(n_240),
.B1(n_0),
.B2(n_2),
.Y(n_270)
);

BUFx2_ASAP7_75t_SL g226 ( 
.A(n_129),
.Y(n_226)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_152),
.A2(n_150),
.B(n_111),
.C(n_119),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_227),
.B(n_232),
.Y(n_284)
);

INVx3_ASAP7_75t_SL g228 ( 
.A(n_116),
.Y(n_228)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_112),
.Y(n_229)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_116),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g233 ( 
.A1(n_160),
.A2(n_36),
.B(n_48),
.Y(n_233)
);

AOI32xp33_ASAP7_75t_L g285 ( 
.A1(n_233),
.A2(n_0),
.A3(n_4),
.B1(n_5),
.B2(n_219),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_148),
.A2(n_48),
.B1(n_43),
.B2(n_27),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_115),
.Y(n_235)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_235),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_163),
.B(n_39),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_139),
.B(n_102),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_135),
.A2(n_43),
.B1(n_22),
.B2(n_10),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_239),
.A2(n_141),
.B1(n_166),
.B2(n_125),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_110),
.A2(n_22),
.B1(n_7),
.B2(n_11),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_145),
.B(n_6),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_6),
.Y(n_278)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_145),
.Y(n_242)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_110),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_153),
.B1(n_146),
.B2(n_140),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_149),
.A2(n_123),
.B1(n_128),
.B2(n_175),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_245),
.A2(n_173),
.B1(n_146),
.B2(n_140),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_166),
.B1(n_149),
.B2(n_153),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_250),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_173),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_253),
.B(n_281),
.C(n_284),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_255),
.A2(n_264),
.B1(n_270),
.B2(n_228),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_274),
.B(n_280),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_186),
.A2(n_0),
.B(n_3),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_275),
.A2(n_269),
.B(n_246),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_212),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_277),
.A2(n_285),
.B1(n_291),
.B2(n_225),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_278),
.B(n_238),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_186),
.A2(n_12),
.B1(n_16),
.B2(n_5),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_279),
.A2(n_256),
.B1(n_272),
.B2(n_263),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_204),
.B(n_0),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_206),
.B(n_0),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_4),
.Y(n_309)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_215),
.Y(n_290)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_213),
.A2(n_181),
.B1(n_182),
.B2(n_220),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_196),
.Y(n_294)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_294),
.Y(n_317)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_196),
.Y(n_296)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_195),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_302),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_216),
.Y(n_302)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_306),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_309),
.B(n_310),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_216),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_312),
.B(n_350),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_257),
.B(n_210),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_313),
.B(n_323),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_261),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_314),
.B(n_330),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_316),
.A2(n_324),
.B1(n_327),
.B2(n_334),
.Y(n_355)
);

OA21x2_ASAP7_75t_L g318 ( 
.A1(n_284),
.A2(n_182),
.B(n_240),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_318),
.A2(n_326),
.B(n_333),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_253),
.B(n_243),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_331),
.C(n_349),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_271),
.B(n_208),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_320),
.B(n_325),
.Y(n_372)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_268),
.Y(n_321)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_259),
.B(n_222),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_269),
.A2(n_288),
.B1(n_270),
.B2(n_275),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_202),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_246),
.A2(n_231),
.B(n_217),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_260),
.A2(n_251),
.B1(n_274),
.B2(n_280),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g331 ( 
.A(n_266),
.B(n_218),
.C(n_214),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_260),
.A2(n_183),
.B(n_189),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_251),
.A2(n_200),
.B1(n_197),
.B2(n_187),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_335),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_301),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_337),
.B(n_339),
.Y(n_377)
);

BUFx24_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_338),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_254),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_185),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_341),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_205),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_303),
.Y(n_342)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_343),
.A2(n_351),
.B1(n_298),
.B2(n_248),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_273),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_348),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_252),
.B(n_199),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_267),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_263),
.A2(n_224),
.B1(n_235),
.B2(n_203),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_346),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_252),
.A2(n_193),
.B1(n_194),
.B2(n_192),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_347),
.A2(n_352),
.B1(n_287),
.B2(n_300),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_256),
.B(n_229),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_268),
.B(n_230),
.C(n_242),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_247),
.B(n_188),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_290),
.A2(n_247),
.B1(n_273),
.B2(n_282),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_262),
.A2(n_180),
.B1(n_221),
.B2(n_4),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_272),
.B(n_262),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_353),
.Y(n_379)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_354),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_358),
.A2(n_368),
.B1(n_376),
.B2(n_389),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_359),
.B(n_335),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_318),
.A2(n_297),
.B1(n_248),
.B2(n_304),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_312),
.B(n_267),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_327),
.Y(n_401)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_315),
.Y(n_370)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_375),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_318),
.A2(n_298),
.B1(n_300),
.B2(n_295),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_345),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_386),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_283),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_381),
.C(n_395),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_328),
.B(n_283),
.C(n_295),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_382),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_384),
.A2(n_387),
.B1(n_392),
.B2(n_396),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_340),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_324),
.A2(n_293),
.B1(n_292),
.B2(n_289),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_307),
.A2(n_258),
.B1(n_293),
.B2(n_292),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_321),
.Y(n_390)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_322),
.A2(n_289),
.B1(n_258),
.B2(n_287),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_317),
.Y(n_394)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_328),
.B(n_276),
.C(n_265),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_333),
.A2(n_276),
.B1(n_265),
.B2(n_5),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_385),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_397),
.B(n_409),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_371),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_310),
.C(n_307),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_405),
.C(n_407),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_356),
.B(n_320),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_358),
.A2(n_314),
.B1(n_339),
.B2(n_329),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_406),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_356),
.B(n_349),
.C(n_311),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_382),
.A2(n_329),
.B1(n_316),
.B2(n_308),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_410),
.A2(n_418),
.B1(n_423),
.B2(n_365),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_363),
.A2(n_326),
.B(n_308),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_412),
.A2(n_425),
.B(n_373),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_378),
.B(n_325),
.Y(n_413)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_413),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_331),
.C(n_317),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_380),
.C(n_371),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_372),
.B(n_309),
.Y(n_416)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_416),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_363),
.A2(n_342),
.B1(n_332),
.B2(n_347),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_392),
.Y(n_419)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_419),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_355),
.A2(n_342),
.B1(n_332),
.B2(n_341),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_420),
.A2(n_427),
.B1(n_429),
.B2(n_430),
.Y(n_440)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_362),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_421),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_377),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_422),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_368),
.A2(n_334),
.B1(n_352),
.B2(n_306),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_372),
.B(n_391),
.Y(n_424)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_424),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_393),
.A2(n_338),
.B(n_354),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_391),
.B(n_305),
.Y(n_426)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_355),
.A2(n_4),
.B1(n_338),
.B2(n_388),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_395),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_360),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_388),
.A2(n_338),
.B1(n_387),
.B2(n_384),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_379),
.A2(n_376),
.B1(n_367),
.B2(n_364),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_396),
.A2(n_393),
.B1(n_364),
.B2(n_361),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_431),
.A2(n_370),
.B1(n_389),
.B2(n_390),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_361),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_432),
.B(n_438),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_444),
.C(n_445),
.Y(n_463)
);

AND2x2_ASAP7_75t_SL g472 ( 
.A(n_437),
.B(n_412),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_441),
.A2(n_454),
.B1(n_461),
.B2(n_417),
.Y(n_485)
);

XOR2x1_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_405),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_449),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_359),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_394),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_420),
.A2(n_365),
.B1(n_362),
.B2(n_375),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_447),
.A2(n_448),
.B1(n_457),
.B2(n_460),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_400),
.B(n_374),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_453),
.C(n_428),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_407),
.B(n_360),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_419),
.A2(n_357),
.B1(n_366),
.B2(n_383),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_421),
.Y(n_455)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_402),
.A2(n_357),
.B1(n_366),
.B2(n_383),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_408),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_397),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_SL g460 ( 
.A1(n_427),
.A2(n_411),
.B1(n_429),
.B2(n_402),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_404),
.A2(n_410),
.B1(n_423),
.B2(n_418),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_440),
.A2(n_425),
.B1(n_413),
.B2(n_424),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_462),
.A2(n_441),
.B1(n_461),
.B2(n_450),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_473),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_453),
.C(n_435),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_468),
.C(n_469),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g504 ( 
.A(n_467),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_414),
.C(n_409),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_416),
.C(n_426),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_443),
.C(n_449),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_470),
.B(n_476),
.C(n_486),
.Y(n_498)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_472),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_411),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_415),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_474),
.Y(n_489)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_446),
.Y(n_475)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_436),
.B(n_415),
.C(n_399),
.Y(n_476)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_478),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_446),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_482),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_437),
.A2(n_398),
.B(n_399),
.Y(n_480)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_480),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_457),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_SL g483 ( 
.A(n_438),
.B(n_398),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_483),
.B(n_451),
.Y(n_488)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_447),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_484),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_485),
.A2(n_442),
.B1(n_454),
.B2(n_439),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_434),
.B(n_417),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_488),
.B(n_507),
.Y(n_514)
);

XOR2x1_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_462),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_490),
.B(n_493),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_472),
.A2(n_474),
.B(n_456),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_493),
.A2(n_499),
.B(n_496),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_470),
.B(n_451),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_481),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_433),
.Y(n_497)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_497),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_472),
.A2(n_450),
.B(n_433),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_500),
.B(n_505),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_501),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_469),
.B(n_477),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_476),
.B(n_473),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_502),
.A2(n_471),
.B1(n_480),
.B2(n_464),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_517),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_466),
.C(n_463),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_510),
.B(n_513),
.C(n_518),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_468),
.Y(n_511)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_511),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_463),
.Y(n_512)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_512),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_465),
.C(n_481),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_520),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_498),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_516),
.A2(n_519),
.B(n_489),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_491),
.B(n_494),
.C(n_490),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_491),
.B(n_496),
.C(n_499),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_487),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_524),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_506),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_522),
.A2(n_506),
.B1(n_492),
.B2(n_502),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_525),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_517),
.A2(n_489),
.B(n_492),
.Y(n_526)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_526),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_497),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_531),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_521),
.A2(n_492),
.B1(n_503),
.B2(n_524),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_533),
.B(n_534),
.Y(n_543)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_509),
.A2(n_503),
.B(n_521),
.C(n_520),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_514),
.A2(n_523),
.B1(n_518),
.B2(n_513),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_537),
.B(n_536),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_536),
.B(n_510),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_538),
.B(n_544),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_529),
.B(n_515),
.Y(n_541)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_541),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_532),
.B(n_537),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_545),
.B(n_546),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_530),
.B(n_526),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_528),
.B(n_533),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_547),
.B(n_527),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_528),
.C(n_527),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_548),
.B(n_551),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_542),
.A2(n_541),
.B(n_539),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_550),
.A2(n_543),
.B(n_535),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_554),
.B(n_549),
.C(n_552),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_548),
.B(n_525),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_555),
.B(n_557),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_553),
.B(n_540),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_558),
.A2(n_556),
.B(n_559),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_560),
.Y(n_561)
);

BUFx24_ASAP7_75t_SL g562 ( 
.A(n_561),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_540),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_563),
.A2(n_535),
.B(n_534),
.Y(n_564)
);


endmodule