module fake_netlist_6_3983_n_1087 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1087);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1087;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1027;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_1079;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_419;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_892;
wire n_768;
wire n_471;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_544;
wire n_372;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_601;
wire n_375;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_843;
wire n_772;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_838;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_972;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_645;
wire n_331;
wire n_916;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_608;
wire n_474;
wire n_683;
wire n_620;
wire n_420;
wire n_630;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_543;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_600;
wire n_464;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_756;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_652;
wire n_553;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_511;
wire n_715;
wire n_467;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_651;
wire n_404;
wire n_439;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_339;
wire n_784;
wire n_434;
wire n_515;
wire n_983;
wire n_427;
wire n_1059;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_663;
wire n_361;
wire n_508;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_1023;
wire n_1013;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;

INVx1_ASAP7_75t_L g325 ( 
.A(n_139),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_117),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_36),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_112),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_318),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_205),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_136),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_196),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_184),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_177),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_106),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_241),
.B(n_279),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_13),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_38),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_233),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_172),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_249),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_137),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_5),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_282),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_270),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_251),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_198),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_61),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_23),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_245),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_193),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_199),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_303),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_73),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_298),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_181),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_308),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_197),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_135),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_290),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_190),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_272),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_10),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_45),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_231),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_26),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_286),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_123),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_226),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_31),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_203),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_134),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_257),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_221),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_24),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_156),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_131),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_14),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_23),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_102),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_238),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_122),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_194),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_246),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_64),
.Y(n_389)
);

BUFx10_ASAP7_75t_L g390 ( 
.A(n_55),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_185),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_206),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_208),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_218),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_43),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_263),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_109),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_248),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_108),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_213),
.Y(n_400)
);

INVx4_ASAP7_75t_R g401 ( 
.A(n_239),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_132),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_274),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_152),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_4),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_141),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_15),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_253),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_275),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_78),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_312),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_195),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_300),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_100),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_204),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_243),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_13),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_307),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_224),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_296),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_211),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_52),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_169),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_301),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_266),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_178),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_40),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_87),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_174),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_244),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_255),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_192),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_64),
.Y(n_433)
);

BUFx5_ASAP7_75t_L g434 ( 
.A(n_126),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_114),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_313),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_268),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_202),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_118),
.Y(n_439)
);

INVx4_ASAP7_75t_R g440 ( 
.A(n_142),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_242),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_273),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_201),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_158),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_235),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_210),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_82),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_93),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_138),
.B(n_154),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_45),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_207),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_219),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_2),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_293),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_124),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_46),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_71),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_157),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_168),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_176),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_220),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_55),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_175),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_121),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_280),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_46),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_71),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_311),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_217),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_191),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_285),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_28),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_247),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_256),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_324),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_97),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_360),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_350),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_453),
.B(n_0),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_453),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_350),
.Y(n_481)
);

BUFx12f_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_360),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_354),
.B(n_451),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_433),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_457),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_327),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_360),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_330),
.B(n_6),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_447),
.B(n_7),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_350),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_373),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_327),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_350),
.B(n_8),
.Y(n_494)
);

OA21x2_ASAP7_75t_L g495 ( 
.A1(n_325),
.A2(n_8),
.B(n_9),
.Y(n_495)
);

BUFx8_ASAP7_75t_SL g496 ( 
.A(n_331),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_400),
.B(n_9),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_367),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_434),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_330),
.B(n_10),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_360),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_394),
.B(n_11),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_466),
.B(n_11),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_332),
.B(n_12),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_400),
.B(n_12),
.Y(n_505)
);

CKINVDCx11_ASAP7_75t_R g506 ( 
.A(n_420),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_419),
.Y(n_507)
);

AOI22x1_ASAP7_75t_SL g508 ( 
.A1(n_338),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_367),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_419),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_326),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_340),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_351),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g514 ( 
.A(n_443),
.B(n_16),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_455),
.B(n_17),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_394),
.B(n_17),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_434),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_366),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_434),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_434),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_369),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_467),
.B(n_18),
.Y(n_524)
);

OA21x2_ASAP7_75t_L g525 ( 
.A1(n_334),
.A2(n_18),
.B(n_19),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_382),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_337),
.A2(n_19),
.B(n_20),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_356),
.Y(n_528)
);

BUFx12f_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_383),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_332),
.B(n_20),
.Y(n_531)
);

INVx6_ASAP7_75t_L g532 ( 
.A(n_437),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_333),
.B(n_21),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_434),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_458),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_335),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_389),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_395),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_452),
.B(n_22),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_405),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_343),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_411),
.B(n_25),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_343),
.B(n_27),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_417),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_411),
.B(n_28),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_339),
.B(n_29),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_463),
.B(n_362),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_362),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_368),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_349),
.B(n_30),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_352),
.A2(n_99),
.B(n_98),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_422),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_427),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_450),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_368),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_456),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_478),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_498),
.B(n_345),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_514),
.B(n_437),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_481),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_491),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_536),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_388),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_514),
.B(n_379),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_511),
.B(n_388),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_536),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_541),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_477),
.Y(n_568)
);

NOR2x1p5_ASAP7_75t_L g569 ( 
.A(n_529),
.B(n_460),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_477),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_477),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_515),
.B(n_479),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_483),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_541),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_492),
.B(n_338),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_489),
.B(n_500),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_483),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_483),
.Y(n_578)
);

INVx8_ASAP7_75t_L g579 ( 
.A(n_497),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_511),
.B(n_393),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_488),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_488),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_541),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_488),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_548),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_501),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_548),
.B(n_549),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_501),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_507),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_484),
.B(n_460),
.Y(n_591)
);

INVxp33_ASAP7_75t_L g592 ( 
.A(n_490),
.Y(n_592)
);

INVx8_ASAP7_75t_L g593 ( 
.A(n_505),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_532),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_507),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_548),
.B(n_393),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_507),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_510),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_515),
.B(n_410),
.C(n_407),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_549),
.B(n_391),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_510),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_L g602 ( 
.A(n_533),
.B(n_428),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_555),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_510),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_532),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_523),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_513),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_555),
.B(n_392),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_484),
.B(n_365),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_576),
.B(n_516),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_588),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_568),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_572),
.A2(n_486),
.B1(n_535),
.B2(n_479),
.Y(n_613)
);

NOR2x1p5_ASAP7_75t_L g614 ( 
.A(n_599),
.B(n_482),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_513),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_571),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_L g617 ( 
.A(n_579),
.B(n_539),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_L g618 ( 
.A(n_579),
.B(n_542),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_576),
.B(n_489),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_592),
.B(n_528),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_571),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_609),
.B(n_528),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_591),
.B(n_500),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_591),
.B(n_504),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_592),
.B(n_504),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_571),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_563),
.B(n_531),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_587),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_580),
.B(n_558),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_560),
.B(n_518),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_572),
.B(n_485),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_605),
.B(n_543),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_587),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_559),
.B(n_543),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_570),
.Y(n_635)
);

BUFx5_ASAP7_75t_L g636 ( 
.A(n_557),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_575),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_559),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_560),
.B(n_561),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_561),
.B(n_520),
.Y(n_640)
);

NAND2x1_ASAP7_75t_L g641 ( 
.A(n_595),
.B(n_401),
.Y(n_641)
);

AO221x1_ASAP7_75t_L g642 ( 
.A1(n_572),
.A2(n_480),
.B1(n_341),
.B2(n_347),
.C(n_344),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_572),
.B(n_602),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_573),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_579),
.B(n_593),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_577),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_581),
.Y(n_647)
);

NAND2x1_ASAP7_75t_L g648 ( 
.A(n_582),
.B(n_440),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_602),
.B(n_506),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_593),
.B(n_523),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_565),
.B(n_487),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_564),
.A2(n_495),
.B1(n_527),
.B2(n_525),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_607),
.B(n_493),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_584),
.B(n_521),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_L g655 ( 
.A(n_596),
.B(n_542),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_607),
.B(n_545),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_586),
.B(n_499),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_607),
.B(n_545),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_586),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_589),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_589),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_590),
.B(n_370),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_590),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_562),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_597),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_598),
.B(n_381),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_598),
.B(n_534),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_601),
.B(n_534),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_601),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_643),
.A2(n_517),
.B(n_502),
.C(n_546),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_644),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_610),
.A2(n_608),
.B(n_600),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_610),
.A2(n_567),
.B(n_566),
.Y(n_673)
);

OAI21xp33_ASAP7_75t_L g674 ( 
.A1(n_613),
.A2(n_524),
.B(n_503),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_623),
.B(n_574),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_624),
.B(n_583),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_652),
.A2(n_634),
.B1(n_642),
.B2(n_638),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_619),
.B(n_585),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_653),
.B(n_371),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_654),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_611),
.B(n_627),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_651),
.B(n_603),
.Y(n_682)
);

OAI21xp33_ASAP7_75t_L g683 ( 
.A1(n_625),
.A2(n_517),
.B(n_502),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_620),
.B(n_386),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_615),
.B(n_398),
.Y(n_685)
);

O2A1O1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_655),
.A2(n_550),
.B(n_546),
.C(n_494),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_654),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_650),
.A2(n_578),
.B(n_604),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_646),
.B(n_647),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_664),
.Y(n_690)
);

AOI21x1_ASAP7_75t_L g691 ( 
.A1(n_657),
.A2(n_606),
.B(n_551),
.Y(n_691)
);

AO21x1_ASAP7_75t_L g692 ( 
.A1(n_618),
.A2(n_550),
.B(n_449),
.Y(n_692)
);

AO21x1_ASAP7_75t_L g693 ( 
.A1(n_656),
.A2(n_449),
.B(n_480),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_637),
.B(n_496),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_659),
.B(n_661),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_645),
.A2(n_525),
.B(n_495),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_658),
.B(n_408),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_649),
.A2(n_617),
.B(n_632),
.C(n_630),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_661),
.B(n_358),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_657),
.A2(n_445),
.B(n_397),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_639),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_661),
.Y(n_702)
);

AOI22x1_ASAP7_75t_L g703 ( 
.A1(n_669),
.A2(n_336),
.B1(n_569),
.B2(n_509),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_662),
.A2(n_416),
.B1(n_425),
.B2(n_414),
.Y(n_704)
);

NOR2x1_ASAP7_75t_L g705 ( 
.A(n_614),
.B(n_454),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_663),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_639),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_666),
.B(n_468),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_612),
.Y(n_709)
);

BUFx4f_ASAP7_75t_L g710 ( 
.A(n_631),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_635),
.B(n_378),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_616),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_667),
.Y(n_713)
);

BUFx12f_ASAP7_75t_L g714 ( 
.A(n_631),
.Y(n_714)
);

AO21x1_ASAP7_75t_L g715 ( 
.A1(n_668),
.A2(n_384),
.B(n_380),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_668),
.A2(n_396),
.B(n_385),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_640),
.A2(n_406),
.B(n_409),
.C(n_399),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_640),
.A2(n_418),
.B(n_413),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_641),
.A2(n_424),
.B(n_426),
.C(n_421),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_R g720 ( 
.A(n_660),
.B(n_328),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_665),
.B(n_429),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_648),
.A2(n_626),
.B(n_621),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_628),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_633),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_636),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_616),
.A2(n_442),
.B(n_441),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_636),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_659),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_629),
.B(n_530),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_622),
.B(n_448),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_654),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_623),
.B(n_459),
.Y(n_732)
);

OAI21xp33_ASAP7_75t_L g733 ( 
.A1(n_613),
.A2(n_519),
.B(n_512),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_654),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_638),
.B(n_329),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_623),
.B(n_461),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_664),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_652),
.A2(n_473),
.B(n_342),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_610),
.A2(n_348),
.B(n_346),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_643),
.A2(n_355),
.B1(n_357),
.B2(n_353),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_623),
.B(n_359),
.Y(n_741)
);

AOI33xp33_ASAP7_75t_L g742 ( 
.A1(n_629),
.A2(n_522),
.A3(n_537),
.B1(n_538),
.B2(n_526),
.B3(n_472),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_613),
.A2(n_363),
.B1(n_364),
.B2(n_361),
.Y(n_743)
);

AOI21x1_ASAP7_75t_L g744 ( 
.A1(n_610),
.A2(n_544),
.B(n_540),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_610),
.A2(n_374),
.B(n_372),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_643),
.A2(n_376),
.B1(n_377),
.B2(n_375),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_623),
.B(n_387),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_613),
.A2(n_403),
.B1(n_404),
.B2(n_402),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_613),
.A2(n_476),
.B(n_462),
.C(n_552),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_708),
.B(n_508),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_672),
.A2(n_415),
.B(n_412),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_701),
.B(n_423),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_722),
.A2(n_691),
.B(n_744),
.Y(n_753)
);

OAI21x1_ASAP7_75t_L g754 ( 
.A1(n_725),
.A2(n_544),
.B(n_540),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_696),
.A2(n_556),
.B(n_554),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_684),
.B(n_679),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_670),
.A2(n_431),
.B(n_430),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_697),
.B(n_432),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_695),
.A2(n_707),
.B(n_678),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_690),
.B(n_553),
.Y(n_760)
);

OAI21x1_ASAP7_75t_SL g761 ( 
.A1(n_692),
.A2(n_103),
.B(n_101),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_737),
.B(n_104),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_681),
.B(n_435),
.Y(n_763)
);

NAND2x1p5_ASAP7_75t_L g764 ( 
.A(n_728),
.B(n_105),
.Y(n_764)
);

O2A1O1Ixp5_ASAP7_75t_L g765 ( 
.A1(n_738),
.A2(n_438),
.B(n_439),
.C(n_436),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_680),
.B(n_444),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_687),
.B(n_446),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_713),
.A2(n_734),
.B(n_731),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_702),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_671),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_673),
.A2(n_110),
.B(n_107),
.Y(n_771)
);

CKINVDCx16_ASAP7_75t_R g772 ( 
.A(n_704),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_675),
.A2(n_465),
.B(n_464),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_729),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_676),
.A2(n_470),
.B(n_469),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_727),
.A2(n_113),
.B(n_111),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_702),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_741),
.B(n_471),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_686),
.A2(n_475),
.B(n_474),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_685),
.B(n_32),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_747),
.B(n_33),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_732),
.B(n_736),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_688),
.A2(n_116),
.B(n_115),
.Y(n_783)
);

BUFx8_ASAP7_75t_L g784 ( 
.A(n_714),
.Y(n_784)
);

AND3x4_ASAP7_75t_L g785 ( 
.A(n_705),
.B(n_34),
.C(n_35),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_677),
.A2(n_120),
.B(n_119),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_683),
.B(n_35),
.Y(n_787)
);

OAI22x1_ASAP7_75t_L g788 ( 
.A1(n_743),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_730),
.B(n_37),
.Y(n_789)
);

AOI221x1_ASAP7_75t_L g790 ( 
.A1(n_733),
.A2(n_128),
.B1(n_129),
.B2(n_127),
.C(n_125),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_706),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_689),
.A2(n_133),
.B(n_130),
.Y(n_792)
);

OR2x6_ASAP7_75t_L g793 ( 
.A(n_749),
.B(n_39),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_694),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_682),
.B(n_40),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_723),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_709),
.B(n_740),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_723),
.B(n_41),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_746),
.B(n_748),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_748),
.B(n_41),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_724),
.A2(n_322),
.B(n_140),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_735),
.B(n_42),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_742),
.B(n_42),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_712),
.Y(n_804)
);

AND2x6_ASAP7_75t_L g805 ( 
.A(n_699),
.B(n_143),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_693),
.B(n_144),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_739),
.A2(n_146),
.B(n_145),
.Y(n_807)
);

OAI21x1_ASAP7_75t_SL g808 ( 
.A1(n_715),
.A2(n_148),
.B(n_147),
.Y(n_808)
);

O2A1O1Ixp5_ASAP7_75t_L g809 ( 
.A1(n_719),
.A2(n_150),
.B(n_151),
.C(n_149),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_745),
.B(n_44),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_SL g811 ( 
.A1(n_717),
.A2(n_44),
.B(n_47),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_710),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_720),
.Y(n_813)
);

AOI21xp33_ASAP7_75t_L g814 ( 
.A1(n_703),
.A2(n_47),
.B(n_48),
.Y(n_814)
);

OAI21x1_ASAP7_75t_L g815 ( 
.A1(n_711),
.A2(n_155),
.B(n_153),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_721),
.Y(n_816)
);

CKINVDCx8_ASAP7_75t_R g817 ( 
.A(n_718),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_700),
.A2(n_160),
.B(n_159),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_726),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_716),
.Y(n_820)
);

AOI21xp33_ASAP7_75t_L g821 ( 
.A1(n_730),
.A2(n_49),
.B(n_50),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_672),
.A2(n_162),
.B(n_161),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_701),
.B(n_50),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_701),
.B(n_51),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_701),
.B(n_53),
.Y(n_825)
);

NOR2xp67_ASAP7_75t_L g826 ( 
.A(n_740),
.B(n_163),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_690),
.B(n_164),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_SL g828 ( 
.A1(n_698),
.A2(n_166),
.B(n_165),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_701),
.B(n_54),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_672),
.A2(n_170),
.B(n_167),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_672),
.A2(n_173),
.B(n_171),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_701),
.B(n_54),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_L g833 ( 
.A1(n_674),
.A2(n_56),
.B(n_57),
.Y(n_833)
);

A2O1A1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_674),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_834)
);

INVx8_ASAP7_75t_L g835 ( 
.A(n_714),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_692),
.A2(n_227),
.B(n_320),
.C(n_319),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_674),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_722),
.A2(n_180),
.B(n_179),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_672),
.A2(n_183),
.B(n_182),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_672),
.A2(n_187),
.B(n_186),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_672),
.A2(n_189),
.B(n_188),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_702),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_708),
.B(n_59),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_701),
.B(n_60),
.Y(n_844)
);

AOI221x1_ASAP7_75t_L g845 ( 
.A1(n_670),
.A2(n_236),
.B1(n_317),
.B2(n_316),
.C(n_315),
.Y(n_845)
);

OAI21x1_ASAP7_75t_L g846 ( 
.A1(n_722),
.A2(n_321),
.B(n_200),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_708),
.B(n_61),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_701),
.B(n_62),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_674),
.A2(n_62),
.B(n_63),
.C(n_65),
.Y(n_849)
);

OAI21x1_ASAP7_75t_L g850 ( 
.A1(n_722),
.A2(n_212),
.B(n_209),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_769),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_774),
.B(n_63),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_768),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_799),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_854)
);

BUFx12f_ASAP7_75t_L g855 ( 
.A(n_784),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_759),
.A2(n_846),
.B(n_838),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_835),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_813),
.B(n_214),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_793),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_789),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_765),
.A2(n_240),
.B(n_306),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_850),
.A2(n_250),
.B(n_305),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_760),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_777),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_843),
.A2(n_69),
.B(n_70),
.C(n_72),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_758),
.A2(n_237),
.B1(n_304),
.B2(n_302),
.Y(n_866)
);

NAND3xp33_ASAP7_75t_L g867 ( 
.A(n_847),
.B(n_69),
.C(n_70),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_772),
.B(n_72),
.Y(n_868)
);

OAI21x1_ASAP7_75t_L g869 ( 
.A1(n_801),
.A2(n_234),
.B(n_299),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_770),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_800),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_871)
);

OA21x2_ASAP7_75t_L g872 ( 
.A1(n_845),
.A2(n_806),
.B(n_790),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_763),
.B(n_74),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_784),
.Y(n_874)
);

AO21x2_ASAP7_75t_L g875 ( 
.A1(n_761),
.A2(n_252),
.B(n_297),
.Y(n_875)
);

NOR2x1_ASAP7_75t_L g876 ( 
.A(n_812),
.B(n_215),
.Y(n_876)
);

AOI22x1_ASAP7_75t_L g877 ( 
.A1(n_779),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_877)
);

OA21x2_ASAP7_75t_L g878 ( 
.A1(n_771),
.A2(n_254),
.B(n_294),
.Y(n_878)
);

OA21x2_ASAP7_75t_L g879 ( 
.A1(n_781),
.A2(n_232),
.B(n_292),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_787),
.A2(n_230),
.B(n_291),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_780),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_881)
);

BUFx2_ASAP7_75t_R g882 ( 
.A(n_817),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_823),
.A2(n_825),
.B(n_824),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_756),
.A2(n_229),
.B1(n_289),
.B2(n_288),
.Y(n_884)
);

AO21x2_ASAP7_75t_L g885 ( 
.A1(n_807),
.A2(n_228),
.B(n_287),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_796),
.Y(n_886)
);

NOR2xp67_ASAP7_75t_SL g887 ( 
.A(n_804),
.B(n_80),
.Y(n_887)
);

OAI21x1_ASAP7_75t_L g888 ( 
.A1(n_783),
.A2(n_776),
.B(n_792),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_791),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_812),
.B(n_83),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_829),
.A2(n_225),
.B(n_284),
.Y(n_891)
);

OA21x2_ASAP7_75t_L g892 ( 
.A1(n_836),
.A2(n_223),
.B(n_283),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_815),
.A2(n_222),
.B(n_281),
.Y(n_893)
);

CKINVDCx11_ASAP7_75t_R g894 ( 
.A(n_794),
.Y(n_894)
);

BUFx2_ASAP7_75t_R g895 ( 
.A(n_797),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_832),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_750),
.B(n_83),
.Y(n_897)
);

AO21x2_ASAP7_75t_L g898 ( 
.A1(n_757),
.A2(n_258),
.B(n_278),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_822),
.A2(n_216),
.B(n_277),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_844),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_830),
.A2(n_841),
.B(n_840),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_831),
.A2(n_314),
.B(n_276),
.Y(n_902)
);

OR2x6_ASAP7_75t_L g903 ( 
.A(n_793),
.B(n_84),
.Y(n_903)
);

INVx6_ASAP7_75t_L g904 ( 
.A(n_794),
.Y(n_904)
);

INVx8_ASAP7_75t_L g905 ( 
.A(n_827),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_816),
.B(n_85),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_762),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_842),
.Y(n_908)
);

NOR2x1_ASAP7_75t_L g909 ( 
.A(n_828),
.B(n_271),
.Y(n_909)
);

OAI21x1_ASAP7_75t_L g910 ( 
.A1(n_839),
.A2(n_269),
.B(n_267),
.Y(n_910)
);

AO21x2_ASAP7_75t_L g911 ( 
.A1(n_808),
.A2(n_265),
.B(n_264),
.Y(n_911)
);

AO21x2_ASAP7_75t_L g912 ( 
.A1(n_778),
.A2(n_262),
.B(n_261),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_848),
.A2(n_260),
.B(n_259),
.Y(n_913)
);

OAI21x1_ASAP7_75t_SL g914 ( 
.A1(n_811),
.A2(n_86),
.B(n_87),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_795),
.A2(n_88),
.B(n_89),
.Y(n_915)
);

OA21x2_ASAP7_75t_L g916 ( 
.A1(n_810),
.A2(n_89),
.B(n_90),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_766),
.A2(n_91),
.B(n_92),
.Y(n_917)
);

AO21x2_ASAP7_75t_L g918 ( 
.A1(n_751),
.A2(n_94),
.B(n_95),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_764),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_818),
.A2(n_96),
.B(n_97),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_826),
.A2(n_802),
.B1(n_767),
.B2(n_752),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_798),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_803),
.Y(n_923)
);

BUFx2_ASAP7_75t_SL g924 ( 
.A(n_805),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_788),
.B(n_821),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_805),
.Y(n_926)
);

AO21x2_ASAP7_75t_L g927 ( 
.A1(n_814),
.A2(n_775),
.B(n_773),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_833),
.B(n_849),
.Y(n_928)
);

OA21x2_ASAP7_75t_L g929 ( 
.A1(n_809),
.A2(n_837),
.B(n_834),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_819),
.Y(n_930)
);

BUFx12f_ASAP7_75t_L g931 ( 
.A(n_805),
.Y(n_931)
);

NAND2x1p5_ASAP7_75t_L g932 ( 
.A(n_820),
.B(n_785),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_820),
.A2(n_753),
.B(n_754),
.Y(n_933)
);

OA21x2_ASAP7_75t_L g934 ( 
.A1(n_755),
.A2(n_696),
.B(n_786),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_799),
.A2(n_643),
.B1(n_768),
.B2(n_638),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_782),
.B(n_681),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_812),
.B(n_762),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_851),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_870),
.Y(n_939)
);

AO21x1_ASAP7_75t_L g940 ( 
.A1(n_935),
.A2(n_883),
.B(n_880),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_863),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_SL g942 ( 
.A1(n_897),
.A2(n_877),
.B1(n_925),
.B2(n_903),
.Y(n_942)
);

OAI221xp5_ASAP7_75t_SL g943 ( 
.A1(n_854),
.A2(n_881),
.B1(n_860),
.B2(n_903),
.C(n_871),
.Y(n_943)
);

AO21x1_ASAP7_75t_SL g944 ( 
.A1(n_915),
.A2(n_917),
.B(n_928),
.Y(n_944)
);

OAI22xp33_ASAP7_75t_L g945 ( 
.A1(n_936),
.A2(n_932),
.B1(n_890),
.B2(n_923),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_857),
.Y(n_946)
);

AO21x1_ASAP7_75t_SL g947 ( 
.A1(n_921),
.A2(n_913),
.B(n_891),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_859),
.Y(n_948)
);

BUFx8_ASAP7_75t_L g949 ( 
.A(n_855),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_882),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_867),
.A2(n_914),
.B1(n_853),
.B2(n_900),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_886),
.Y(n_952)
);

AO21x1_ASAP7_75t_L g953 ( 
.A1(n_861),
.A2(n_922),
.B(n_873),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_933),
.A2(n_856),
.B(n_888),
.Y(n_954)
);

AO21x1_ASAP7_75t_L g955 ( 
.A1(n_922),
.A2(n_900),
.B(n_896),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_904),
.Y(n_956)
);

BUFx8_ASAP7_75t_SL g957 ( 
.A(n_874),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_894),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_SL g959 ( 
.A1(n_890),
.A2(n_868),
.B1(n_906),
.B2(n_852),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_864),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_937),
.B(n_930),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_907),
.B(n_895),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_901),
.A2(n_869),
.B(n_862),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_899),
.A2(n_910),
.B(n_902),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_864),
.Y(n_965)
);

OR2x6_ASAP7_75t_L g966 ( 
.A(n_905),
.B(n_919),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_918),
.A2(n_885),
.B1(n_898),
.B2(n_929),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_864),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_865),
.B(n_858),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_908),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_889),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_918),
.A2(n_898),
.B1(n_929),
.B2(n_916),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_887),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_919),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_920),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_866),
.A2(n_909),
.B1(n_872),
.B2(n_884),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_926),
.B(n_927),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_876),
.Y(n_978)
);

BUFx4f_ASAP7_75t_SL g979 ( 
.A(n_931),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_879),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_924),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_893),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_912),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_911),
.B(n_875),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_934),
.B(n_892),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_878),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_939),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_941),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_941),
.B(n_934),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_971),
.Y(n_990)
);

NAND2x1p5_ASAP7_75t_L g991 ( 
.A(n_981),
.B(n_974),
.Y(n_991)
);

INVx3_ASAP7_75t_SL g992 ( 
.A(n_958),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_962),
.B(n_950),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_942),
.A2(n_944),
.B1(n_959),
.B2(n_940),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_948),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_938),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_943),
.B(n_945),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_951),
.B(n_952),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_951),
.B(n_942),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_971),
.Y(n_1000)
);

AOI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_943),
.A2(n_959),
.B1(n_969),
.B2(n_976),
.C(n_953),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_975),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_966),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_980),
.Y(n_1004)
);

INVxp67_ASAP7_75t_SL g1005 ( 
.A(n_955),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_965),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_961),
.B(n_978),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_956),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_970),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_946),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_966),
.Y(n_1011)
);

AO31x2_ASAP7_75t_L g1012 ( 
.A1(n_983),
.A2(n_985),
.A3(n_986),
.B(n_977),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_968),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_968),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_961),
.B(n_947),
.Y(n_1015)
);

BUFx12f_ASAP7_75t_L g1016 ( 
.A(n_949),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_973),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_984),
.B(n_972),
.Y(n_1018)
);

INVx8_ASAP7_75t_L g1019 ( 
.A(n_960),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_960),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_960),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_990),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_1003),
.B(n_982),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1004),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_1003),
.B(n_1011),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_1001),
.B(n_967),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1000),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1018),
.B(n_967),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_991),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1000),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_997),
.A2(n_979),
.B1(n_949),
.B2(n_957),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_987),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_995),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_999),
.A2(n_994),
.B1(n_1017),
.B2(n_1007),
.Y(n_1034)
);

INVxp67_ASAP7_75t_SL g1035 ( 
.A(n_988),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_988),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_1015),
.B(n_964),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_999),
.B(n_954),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_994),
.A2(n_963),
.B1(n_993),
.B2(n_1015),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_989),
.B(n_998),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_1024),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_1026),
.B(n_998),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_1040),
.B(n_1012),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_1026),
.B(n_991),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_1036),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_1023),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1035),
.B(n_1009),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_1025),
.B(n_1002),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1022),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1038),
.B(n_1006),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1027),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1030),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1032),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1053),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1041),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1046),
.B(n_1028),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_SL g1057 ( 
.A(n_1043),
.B(n_1029),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1041),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1042),
.A2(n_1034),
.B1(n_1031),
.B2(n_1039),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1046),
.B(n_1050),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_1045),
.B(n_1037),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1059),
.A2(n_1044),
.B(n_1034),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_1061),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1054),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_1056),
.B(n_1048),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_1055),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1058),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_SL g1068 ( 
.A1(n_1062),
.A2(n_1057),
.B(n_1005),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1064),
.Y(n_1069)
);

NAND2x1_ASAP7_75t_L g1070 ( 
.A(n_1068),
.B(n_1066),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1068),
.A2(n_1047),
.B(n_1063),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1069),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_SL g1073 ( 
.A(n_1070),
.B(n_1071),
.C(n_1033),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1072),
.Y(n_1074)
);

NOR2xp67_ASAP7_75t_L g1075 ( 
.A(n_1073),
.B(n_1016),
.Y(n_1075)
);

NAND4xp75_ASAP7_75t_L g1076 ( 
.A(n_1074),
.B(n_1049),
.C(n_1051),
.D(n_1052),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_1075),
.B(n_992),
.Y(n_1077)
);

OA22x2_ASAP7_75t_L g1078 ( 
.A1(n_1077),
.A2(n_992),
.B1(n_1076),
.B2(n_1065),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1078),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1079),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1080),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_SL g1082 ( 
.A1(n_1081),
.A2(n_1010),
.B(n_1008),
.Y(n_1082)
);

AOI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_1082),
.A2(n_1020),
.B1(n_1021),
.B2(n_1014),
.C(n_1013),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1083),
.B(n_1067),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1084),
.B(n_1060),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_1085),
.B(n_1019),
.Y(n_1086)
);

AOI21xp33_ASAP7_75t_SL g1087 ( 
.A1(n_1086),
.A2(n_1019),
.B(n_996),
.Y(n_1087)
);


endmodule