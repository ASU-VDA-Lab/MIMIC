module fake_jpeg_16394_n_273 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_21;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_33),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_22),
.B1(n_23),
.B2(n_16),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_45),
.B1(n_13),
.B2(n_14),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_23),
.B1(n_16),
.B2(n_13),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_26),
.B1(n_25),
.B2(n_14),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_26),
.B1(n_42),
.B2(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_31),
.B1(n_29),
.B2(n_35),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_64),
.B1(n_33),
.B2(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_18),
.B1(n_49),
.B2(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_68),
.Y(n_82)
);

AO22x1_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_48),
.B1(n_47),
.B2(n_44),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_40),
.B(n_32),
.C(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_80),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_63),
.B1(n_60),
.B2(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_18),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_40),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_57),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_105),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_34),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_92),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_36),
.C(n_34),
.Y(n_92)
);

OAI22x1_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_19),
.B1(n_17),
.B2(n_28),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_73),
.B1(n_48),
.B2(n_44),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_102),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_36),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_59),
.B1(n_28),
.B2(n_43),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_98),
.B1(n_85),
.B2(n_101),
.Y(n_125)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_107),
.B(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_70),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_77),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_76),
.B1(n_47),
.B2(n_44),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_121),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_87),
.B(n_76),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_125),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_74),
.A3(n_82),
.B1(n_77),
.B2(n_71),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_81),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_133),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_92),
.C(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_142),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_94),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_140),
.C(n_145),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_94),
.C(n_84),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_67),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_71),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_106),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_106),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_111),
.C(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_15),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_150),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_122),
.B(n_118),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_169),
.B(n_151),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_157),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_113),
.C(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_158),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_120),
.C(n_108),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_108),
.B1(n_72),
.B2(n_28),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_165),
.B1(n_166),
.B2(n_170),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_161),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_108),
.B1(n_72),
.B2(n_3),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_72),
.B1(n_2),
.B2(n_3),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_1),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_148),
.A2(n_67),
.B(n_30),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_172),
.A2(n_150),
.B(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_179),
.Y(n_202)
);

NOR3xp33_ASAP7_75t_SL g179 ( 
.A(n_164),
.B(n_149),
.C(n_136),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_169),
.A2(n_133),
.B1(n_146),
.B2(n_145),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_192),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_129),
.C(n_30),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_172),
.C(n_158),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_185),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_129),
.B1(n_2),
.B2(n_4),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_170),
.B1(n_166),
.B2(n_154),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_36),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_165),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_155),
.B1(n_156),
.B2(n_169),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_36),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_207),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_182),
.B1(n_188),
.B2(n_32),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_153),
.C(n_40),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_205),
.C(n_208),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_191),
.B1(n_186),
.B2(n_179),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_210),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_153),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_34),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_34),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_180),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_32),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_211)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_218),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_196),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_223),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_221),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_19),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_12),
.B1(n_11),
.B2(n_7),
.Y(n_229)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_206),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_194),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_238),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_222),
.A2(n_200),
.B(n_201),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_224),
.B(n_212),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_219),
.B(n_209),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_12),
.B1(n_11),
.B2(n_8),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_239),
.C(n_225),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_17),
.Y(n_239)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_246),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_214),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_21),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_213),
.B(n_218),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_17),
.C(n_21),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_248),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_17),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_21),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_10),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_245),
.A2(n_244),
.B(n_231),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_251),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_233),
.B1(n_234),
.B2(n_238),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_241),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_262),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_242),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_255),
.B1(n_11),
.B2(n_8),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_15),
.C(n_20),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_265),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_258),
.B(n_12),
.Y(n_267)
);

O2A1O1Ixp33_ASAP7_75t_SL g268 ( 
.A1(n_267),
.A2(n_264),
.B(n_9),
.C(n_10),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_266),
.C(n_20),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_269),
.B(n_5),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_5),
.B(n_6),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_20),
.C(n_15),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_20),
.Y(n_273)
);


endmodule