module fake_jpeg_30612_n_54 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_54);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_54;

wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_3),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_7),
.B1(n_17),
.B2(n_16),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_1),
.B(n_2),
.Y(n_35)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_24),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_35),
.B(n_37),
.Y(n_39)
);

NOR4xp25_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_19),
.C(n_2),
.D(n_3),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_23),
.C(n_29),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_24),
.B1(n_23),
.B2(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_27),
.B1(n_5),
.B2(n_4),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_5),
.B1(n_24),
.B2(n_9),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_48),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_8),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_10),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_46),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_51),
.B(n_46),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_50),
.B(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_18),
.Y(n_54)
);


endmodule