module fake_netlist_6_2291_n_1220 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1220);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1220;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_881;
wire n_1199;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1027;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_1212;
wire n_226;
wire n_828;
wire n_208;
wire n_161;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_168;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_1203;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1217;
wire n_751;
wire n_449;
wire n_749;
wire n_1208;
wire n_798;
wire n_188;
wire n_1164;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_1209;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_1214;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1204;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_1192;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_963;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_1120;
wire n_369;
wire n_894;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_814;
wire n_389;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_1139;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_1206;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_1196;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_601;
wire n_375;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_1205;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_1163;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_1219;
wire n_1216;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_1213;
wire n_638;
wire n_234;
wire n_1181;
wire n_910;
wire n_901;
wire n_1211;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_172;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_1215;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1193;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_163;
wire n_717;
wire n_1152;
wire n_330;
wire n_771;
wire n_1121;
wire n_1145;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_1195;
wire n_356;
wire n_577;
wire n_166;
wire n_936;
wire n_184;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_813;
wire n_395;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_1201;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_1218;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_1198;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1194;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_386;
wire n_201;
wire n_249;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_162;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_652;
wire n_553;
wire n_849;
wire n_1107;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1207;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_1167;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_404;
wire n_651;
wire n_271;
wire n_439;
wire n_1153;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_1210;
wire n_679;
wire n_1069;
wire n_1185;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_1175;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1200;
wire n_1059;
wire n_1197;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_165;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1154;
wire n_177;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_170;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_410;
wire n_398;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_664;
wire n_171;
wire n_949;
wire n_678;
wire n_192;
wire n_169;
wire n_1007;
wire n_649;
wire n_855;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_38),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_49),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_142),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_64),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_59),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_15),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_20),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_43),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_4),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_155),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_17),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_56),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_77),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_6),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_86),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_47),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_81),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_29),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_33),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_15),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_23),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_42),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_34),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_1),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_45),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_13),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_60),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_122),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_46),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_73),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_76),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_24),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_132),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_37),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_18),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_22),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_99),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_88),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_39),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_82),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_46),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_55),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_124),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_134),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_14),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_141),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_92),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_100),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_12),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_62),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_48),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_70),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_130),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_160),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_21),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_103),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_145),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_97),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_75),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_24),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_56),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_20),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_30),
.Y(n_244)
);

BUFx8_ASAP7_75t_SL g245 ( 
.A(n_43),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_3),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_44),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_84),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_135),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_33),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_107),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_10),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_112),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_85),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_158),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_153),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_0),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_6),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_118),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_12),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_149),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_31),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_95),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_148),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_57),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_48),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_8),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_67),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_44),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_146),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_8),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_138),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_154),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_16),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_17),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_98),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_7),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_55),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_89),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_121),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_139),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_255),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_208),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_168),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_164),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_168),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_173),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_173),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_190),
.B(n_203),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_179),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_175),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_180),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_175),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_180),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_245),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_186),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_215),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_187),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_163),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_215),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_225),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_190),
.B(n_0),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_225),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_172),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_206),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_217),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_162),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_203),
.B(n_1),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_186),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_170),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_189),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_273),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_236),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_161),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_189),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_205),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_240),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_165),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_166),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_205),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_171),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_240),
.B(n_2),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_241),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_162),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_174),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_172),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_177),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_227),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_178),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_210),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_270),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_181),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_183),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_227),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_169),
.B(n_2),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_210),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_169),
.B(n_3),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_213),
.B(n_4),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_191),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_167),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_270),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_211),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_211),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_192),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_212),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_212),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_219),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_195),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_182),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_184),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_200),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_219),
.Y(n_354)
);

INVxp33_ASAP7_75t_SL g355 ( 
.A(n_198),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_201),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_214),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_218),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_220),
.Y(n_359)
);

INVxp33_ASAP7_75t_SL g360 ( 
.A(n_230),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_221),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_242),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_243),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_174),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_252),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_185),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_185),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_188),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_209),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_216),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_223),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_188),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_317),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_293),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_293),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_295),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_295),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_286),
.B(n_194),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_301),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_328),
.B(n_276),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_224),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_309),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_299),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_336),
.B(n_281),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_309),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_285),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_327),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_299),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_291),
.B(n_270),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_304),
.B(n_270),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_327),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_302),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_364),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_302),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_364),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_303),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_303),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_305),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_366),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_306),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_339),
.B(n_176),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_367),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_310),
.B(n_204),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_305),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_284),
.B(n_276),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_306),
.B(n_276),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_287),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_289),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_285),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_290),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_316),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_301),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_367),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_294),
.A2(n_256),
.B(n_207),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_296),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_315),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_372),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_298),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_311),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_313),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_318),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_322),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_332),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_338),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_345),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_292),
.B(n_300),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_315),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_347),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_337),
.B(n_228),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_349),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_354),
.B(n_265),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_361),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_326),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_340),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_312),
.B(n_213),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_312),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_324),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_405),
.B(n_282),
.Y(n_443)
);

INVx11_ASAP7_75t_L g444 ( 
.A(n_440),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_405),
.B(n_288),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_416),
.Y(n_446)
);

OR2x6_ASAP7_75t_L g447 ( 
.A(n_442),
.B(n_441),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_435),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_435),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_373),
.Y(n_450)
);

NAND2x1p5_ASAP7_75t_L g451 ( 
.A(n_416),
.B(n_221),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_435),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_390),
.B(n_355),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_435),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_373),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_403),
.B(n_333),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_390),
.A2(n_319),
.B1(n_202),
.B2(n_283),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_413),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_376),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_379),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_442),
.A2(n_325),
.B1(n_265),
.B2(n_193),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_403),
.B(n_343),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_419),
.B(n_329),
.C(n_323),
.Y(n_463)
);

BUFx10_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_413),
.Y(n_467)
);

OAI22x1_ASAP7_75t_L g468 ( 
.A1(n_391),
.A2(n_341),
.B1(n_362),
.B2(n_359),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_373),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_376),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_435),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_376),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_442),
.A2(n_269),
.B1(n_196),
.B2(n_199),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_391),
.B(n_360),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_373),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_442),
.B(n_365),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_376),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_376),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_381),
.B(n_408),
.Y(n_479)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_373),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_426),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_376),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_442),
.B(n_323),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_376),
.Y(n_484)
);

NOR2x1p5_ASAP7_75t_L g485 ( 
.A(n_441),
.B(n_297),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_442),
.A2(n_307),
.B1(n_308),
.B2(n_314),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_411),
.B(n_329),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_381),
.A2(n_193),
.B1(n_196),
.B2(n_232),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_411),
.A2(n_267),
.B1(n_258),
.B2(n_262),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_426),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_382),
.B(n_320),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_430),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_382),
.B(n_321),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_440),
.A2(n_371),
.B1(n_370),
.B2(n_369),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_426),
.Y(n_495)
);

AND3x4_ASAP7_75t_L g496 ( 
.A(n_419),
.B(n_334),
.C(n_331),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_374),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_373),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_411),
.B(n_331),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_423),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_441),
.B(n_334),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_423),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_381),
.A2(n_250),
.B1(n_199),
.B2(n_275),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_373),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_374),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_417),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_387),
.B(n_335),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_408),
.B(n_368),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_417),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_424),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_441),
.B(n_335),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_474),
.B(n_441),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_483),
.B(n_434),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_479),
.B(n_434),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_479),
.B(n_401),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_481),
.B(n_385),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_481),
.B(n_385),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_497),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_401),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_453),
.B(n_342),
.Y(n_523)
);

BUFx5_ASAP7_75t_L g524 ( 
.A(n_464),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_464),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_473),
.A2(n_407),
.B1(n_431),
.B2(n_207),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_448),
.Y(n_527)
);

NOR3xp33_ASAP7_75t_L g528 ( 
.A(n_463),
.B(n_414),
.C(n_380),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_497),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_497),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_462),
.B(n_351),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_466),
.B(n_401),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_448),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_449),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_408),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_500),
.B(n_401),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_491),
.A2(n_414),
.B1(n_380),
.B2(n_353),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_500),
.B(n_502),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_L g539 ( 
.A(n_451),
.B(n_197),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_502),
.B(n_509),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_509),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_511),
.B(n_401),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_466),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_511),
.A2(n_512),
.B1(n_447),
.B2(n_503),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_512),
.B(n_439),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_449),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_493),
.B(n_380),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_452),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_464),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_452),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_499),
.B(n_414),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_454),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_505),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_447),
.A2(n_407),
.B1(n_431),
.B2(n_261),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_454),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_461),
.B(n_439),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_471),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_464),
.B(n_417),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_505),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_471),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_499),
.B(n_352),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_456),
.B(n_356),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_443),
.B(n_341),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_466),
.B(n_417),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_490),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_476),
.A2(n_407),
.B1(n_350),
.B2(n_357),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_505),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_446),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_451),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_447),
.A2(n_407),
.B1(n_261),
.B2(n_256),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_447),
.B(n_438),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_467),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_507),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_451),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_507),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_447),
.A2(n_444),
.B1(n_457),
.B2(n_501),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_459),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_457),
.B(n_346),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_488),
.A2(n_407),
.B1(n_226),
.B2(n_234),
.Y(n_579)
);

NOR2xp67_ASAP7_75t_L g580 ( 
.A(n_468),
.B(n_346),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_490),
.B(n_417),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_459),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_489),
.B(n_350),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_490),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_495),
.B(n_417),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_495),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_495),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_445),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_487),
.B(n_357),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_444),
.B(n_358),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_489),
.B(n_358),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_450),
.B(n_417),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_513),
.B(n_359),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_L g594 ( 
.A(n_468),
.B(n_362),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_459),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_450),
.B(n_422),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_450),
.B(n_422),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_494),
.B(n_363),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_450),
.B(n_422),
.Y(n_599)
);

NOR2xp67_ASAP7_75t_L g600 ( 
.A(n_455),
.B(n_363),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_496),
.B(n_297),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_470),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_496),
.B(n_438),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_460),
.B(n_379),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_470),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_492),
.B(n_379),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_496),
.A2(n_263),
.B1(n_226),
.B2(n_231),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_486),
.B(n_436),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_470),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_485),
.B(n_430),
.Y(n_610)
);

NOR2xp67_ASAP7_75t_L g611 ( 
.A(n_455),
.B(n_430),
.Y(n_611)
);

O2A1O1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_517),
.A2(n_427),
.B(n_429),
.C(n_425),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_516),
.B(n_420),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_547),
.B(n_427),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_588),
.B(n_429),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_572),
.B(n_458),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_519),
.B(n_420),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_573),
.B(n_485),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_572),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_576),
.A2(n_514),
.B(n_568),
.C(n_545),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_573),
.B(n_436),
.Y(n_621)
);

AO21x1_ASAP7_75t_L g622 ( 
.A1(n_539),
.A2(n_569),
.B(n_568),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_520),
.B(n_420),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_535),
.B(n_436),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_603),
.A2(n_238),
.B(n_231),
.C(n_234),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_549),
.A2(n_498),
.B(n_469),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_524),
.B(n_472),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_544),
.A2(n_263),
.B1(n_259),
.B2(n_238),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_535),
.B(n_432),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_549),
.A2(n_498),
.B(n_469),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_522),
.B(n_420),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_565),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g633 ( 
.A1(n_539),
.A2(n_416),
.B(n_472),
.Y(n_633)
);

NOR3xp33_ASAP7_75t_L g634 ( 
.A(n_523),
.B(n_433),
.C(n_432),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_541),
.B(n_420),
.Y(n_635)
);

O2A1O1Ixp5_ASAP7_75t_L g636 ( 
.A1(n_538),
.A2(n_472),
.B(n_478),
.C(n_477),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_540),
.B(n_455),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_549),
.B(n_433),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_527),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_518),
.B(n_571),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_565),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_518),
.B(n_455),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_575),
.B(n_437),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_549),
.A2(n_498),
.B(n_469),
.Y(n_644)
);

BUFx4f_ASAP7_75t_L g645 ( 
.A(n_515),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_578),
.A2(n_437),
.B(n_259),
.C(n_383),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_549),
.B(n_506),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_518),
.A2(n_475),
.B1(n_504),
.B2(n_510),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_525),
.A2(n_498),
.B(n_469),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_556),
.A2(n_484),
.B(n_482),
.C(n_478),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_571),
.B(n_475),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_575),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_525),
.A2(n_510),
.B(n_506),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_525),
.A2(n_510),
.B(n_506),
.Y(n_654)
);

O2A1O1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_551),
.A2(n_400),
.B(n_383),
.C(n_386),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_515),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_556),
.B(n_475),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_531),
.A2(n_475),
.B1(n_504),
.B2(n_510),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_537),
.B(n_266),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_565),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_565),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_608),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_610),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_558),
.A2(n_506),
.B(n_478),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_532),
.A2(n_506),
.B(n_482),
.Y(n_665)
);

NOR2x2_ASAP7_75t_L g666 ( 
.A(n_607),
.B(n_409),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_527),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_533),
.B(n_504),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_611),
.B(n_222),
.Y(n_669)
);

O2A1O1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_583),
.A2(n_404),
.B(n_402),
.C(n_415),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_574),
.A2(n_482),
.B(n_477),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_524),
.B(n_506),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_533),
.B(n_504),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_532),
.A2(n_484),
.B(n_477),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_SL g675 ( 
.A(n_610),
.B(n_229),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_532),
.A2(n_484),
.B(n_480),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_574),
.A2(n_480),
.B(n_410),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_604),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_564),
.A2(n_585),
.B(n_581),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_570),
.A2(n_480),
.B(n_374),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_591),
.A2(n_402),
.B(n_388),
.C(n_392),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_524),
.B(n_233),
.Y(n_682)
);

AO21x1_ASAP7_75t_L g683 ( 
.A1(n_569),
.A2(n_232),
.B(n_222),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_534),
.B(n_422),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_608),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_536),
.A2(n_480),
.B(n_428),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_554),
.A2(n_249),
.B1(n_251),
.B2(n_253),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_562),
.A2(n_422),
.B1(n_428),
.B2(n_268),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_534),
.A2(n_480),
.B(n_410),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_555),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_555),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_565),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_590),
.B(n_274),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_557),
.B(n_422),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_604),
.Y(n_695)
);

O2A1O1Ixp5_ASAP7_75t_L g696 ( 
.A1(n_557),
.A2(n_409),
.B(n_421),
.C(n_410),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_543),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_606),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_560),
.A2(n_480),
.B(n_412),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_524),
.B(n_235),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_542),
.A2(n_428),
.B(n_422),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_560),
.B(n_428),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_546),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_600),
.B(n_428),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_524),
.A2(n_428),
.B(n_412),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_524),
.A2(n_428),
.B(n_412),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_548),
.A2(n_421),
.B(n_409),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_656),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_662),
.B(n_561),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_632),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_693),
.A2(n_598),
.B(n_593),
.C(n_528),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_645),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_639),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_645),
.B(n_524),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_693),
.A2(n_563),
.B1(n_589),
.B2(n_601),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_624),
.B(n_543),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_662),
.B(n_586),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_667),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_619),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_679),
.A2(n_596),
.B(n_592),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_626),
.A2(n_524),
.B(n_630),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_621),
.B(n_606),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_R g723 ( 
.A(n_616),
.B(n_584),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_632),
.Y(n_724)
);

NAND2x1p5_ASAP7_75t_L g725 ( 
.A(n_632),
.B(n_586),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_644),
.A2(n_587),
.B(n_597),
.Y(n_726)
);

NOR2x1_ASAP7_75t_L g727 ( 
.A(n_678),
.B(n_580),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_634),
.B(n_640),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_685),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_685),
.B(n_526),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_690),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_SL g732 ( 
.A(n_659),
.B(n_566),
.C(n_579),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_632),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_613),
.A2(n_587),
.B(n_599),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_628),
.A2(n_550),
.B1(n_552),
.B2(n_278),
.Y(n_735)
);

O2A1O1Ixp5_ASAP7_75t_L g736 ( 
.A1(n_622),
.A2(n_605),
.B(n_602),
.C(n_609),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_634),
.A2(n_594),
.B1(n_605),
.B2(n_602),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_695),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_620),
.A2(n_582),
.B1(n_577),
.B2(n_595),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_652),
.B(n_698),
.Y(n_740)
);

AOI221xp5_ASAP7_75t_L g741 ( 
.A1(n_659),
.A2(n_277),
.B1(n_278),
.B2(n_257),
.C(n_275),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_631),
.A2(n_582),
.B(n_577),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_652),
.B(n_595),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_629),
.B(n_567),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_615),
.B(n_567),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_615),
.B(n_521),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_691),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_677),
.A2(n_529),
.B(n_521),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_703),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_663),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_614),
.A2(n_559),
.B(n_553),
.C(n_530),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_642),
.A2(n_530),
.B(n_529),
.Y(n_752)
);

AOI21x1_ASAP7_75t_L g753 ( 
.A1(n_682),
.A2(n_559),
.B(n_553),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_697),
.B(n_386),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_614),
.B(n_237),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_643),
.B(n_421),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_618),
.B(n_388),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_SL g758 ( 
.A1(n_625),
.A2(n_246),
.B(n_247),
.C(n_250),
.Y(n_758)
);

O2A1O1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_612),
.A2(n_244),
.B(n_246),
.C(n_247),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_669),
.B(n_392),
.Y(n_760)
);

BUFx4f_ASAP7_75t_L g761 ( 
.A(n_669),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_657),
.B(n_418),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_672),
.A2(n_375),
.B(n_377),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_641),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_697),
.B(n_239),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_675),
.A2(n_264),
.B1(n_279),
.B2(n_248),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_617),
.B(n_418),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_653),
.A2(n_375),
.B(n_377),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_635),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_623),
.B(n_394),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_669),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_641),
.B(n_254),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_749),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_715),
.A2(n_670),
.B(n_681),
.C(n_655),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_736),
.A2(n_650),
.B(n_696),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_736),
.A2(n_696),
.B(n_636),
.Y(n_776)
);

CKINVDCx8_ASAP7_75t_R g777 ( 
.A(n_719),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_713),
.Y(n_778)
);

OAI221xp5_ASAP7_75t_SL g779 ( 
.A1(n_741),
.A2(n_646),
.B1(n_666),
.B2(n_688),
.C(n_269),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_734),
.A2(n_636),
.B(n_674),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_721),
.A2(n_700),
.B(n_704),
.Y(n_781)
);

AOI221x1_ASAP7_75t_L g782 ( 
.A1(n_732),
.A2(n_633),
.B1(n_671),
.B2(n_689),
.C(n_699),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_726),
.A2(n_654),
.B(n_649),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_720),
.A2(n_664),
.B(n_665),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_729),
.B(n_641),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_718),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_767),
.A2(n_647),
.B(n_637),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_709),
.A2(n_687),
.B1(n_638),
.B2(n_651),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_708),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_742),
.A2(n_706),
.B(n_705),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_738),
.B(n_641),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_731),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_748),
.A2(n_676),
.B(n_701),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_711),
.A2(n_658),
.B(n_707),
.C(n_648),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_747),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_752),
.A2(n_694),
.B(n_684),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_709),
.A2(n_680),
.B(n_686),
.C(n_702),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_746),
.A2(n_692),
.B1(n_660),
.B2(n_661),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_SL g799 ( 
.A1(n_728),
.A2(n_668),
.B(n_673),
.C(n_627),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_761),
.A2(n_257),
.B1(n_244),
.B2(n_271),
.Y(n_800)
);

AO31x2_ASAP7_75t_L g801 ( 
.A1(n_739),
.A2(n_683),
.A3(n_271),
.B(n_260),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_712),
.Y(n_802)
);

INVx3_ASAP7_75t_R g803 ( 
.A(n_722),
.Y(n_803)
);

AO31x2_ASAP7_75t_L g804 ( 
.A1(n_751),
.A2(n_260),
.A3(n_400),
.B(n_404),
.Y(n_804)
);

AOI21x1_ASAP7_75t_L g805 ( 
.A1(n_753),
.A2(n_627),
.B(n_378),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_770),
.A2(n_692),
.B(n_661),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_746),
.A2(n_692),
.B1(n_661),
.B2(n_660),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_724),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_729),
.Y(n_809)
);

OAI22x1_ASAP7_75t_L g810 ( 
.A1(n_771),
.A2(n_272),
.B1(n_280),
.B2(n_394),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_750),
.B(n_660),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_757),
.B(n_660),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_762),
.A2(n_415),
.B(n_396),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_768),
.A2(n_769),
.B(n_730),
.Y(n_814)
);

O2A1O1Ixp5_ASAP7_75t_SL g815 ( 
.A1(n_755),
.A2(n_396),
.B(n_378),
.C(n_393),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_714),
.A2(n_692),
.B(n_661),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_740),
.A2(n_406),
.B(n_397),
.C(n_393),
.Y(n_817)
);

OAI21x1_ASAP7_75t_L g818 ( 
.A1(n_763),
.A2(n_397),
.B(n_393),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_737),
.A2(n_393),
.B(n_397),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_745),
.A2(n_393),
.B(n_397),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_756),
.B(n_397),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_724),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_754),
.B(n_406),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_754),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_743),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_725),
.A2(n_406),
.B(n_375),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_740),
.A2(n_377),
.B(n_7),
.C(n_9),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_802),
.Y(n_828)
);

BUFx8_ASAP7_75t_L g829 ( 
.A(n_811),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_773),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_808),
.Y(n_831)
);

CKINVDCx11_ASAP7_75t_R g832 ( 
.A(n_777),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_803),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_800),
.A2(n_761),
.B1(n_756),
.B2(n_760),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_789),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_778),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_786),
.Y(n_837)
);

INVx6_ASAP7_75t_L g838 ( 
.A(n_811),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_825),
.A2(n_760),
.B1(n_717),
.B2(n_727),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_SL g840 ( 
.A1(n_779),
.A2(n_723),
.B1(n_716),
.B2(n_743),
.Y(n_840)
);

BUFx4f_ASAP7_75t_SL g841 ( 
.A(n_808),
.Y(n_841)
);

NAND2x1p5_ASAP7_75t_L g842 ( 
.A(n_812),
.B(n_764),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_792),
.A2(n_744),
.B1(n_735),
.B2(n_765),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_809),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_810),
.A2(n_735),
.B1(n_772),
.B2(n_766),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_795),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_SL g847 ( 
.A1(n_824),
.A2(n_725),
.B1(n_724),
.B2(n_710),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_788),
.A2(n_764),
.B1(n_724),
.B2(n_710),
.Y(n_848)
);

INVx8_ASAP7_75t_L g849 ( 
.A(n_808),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_822),
.Y(n_850)
);

INVx3_ASAP7_75t_SL g851 ( 
.A(n_785),
.Y(n_851)
);

INVx6_ASAP7_75t_L g852 ( 
.A(n_785),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_L g853 ( 
.A1(n_782),
.A2(n_733),
.B1(n_197),
.B2(n_759),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_822),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_SL g855 ( 
.A1(n_798),
.A2(n_733),
.B1(n_197),
.B2(n_758),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_804),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_823),
.B(n_377),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_823),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_SL g859 ( 
.A1(n_798),
.A2(n_197),
.B1(n_9),
.B2(n_10),
.Y(n_859)
);

INVx6_ASAP7_75t_L g860 ( 
.A(n_791),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_SL g861 ( 
.A1(n_807),
.A2(n_197),
.B1(n_11),
.B2(n_13),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_821),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_804),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_814),
.B(n_377),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_SL g865 ( 
.A1(n_807),
.A2(n_197),
.B1(n_11),
.B2(n_14),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_804),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_814),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_826),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_801),
.Y(n_869)
);

OAI22xp33_ASAP7_75t_L g870 ( 
.A1(n_813),
.A2(n_5),
.B1(n_16),
.B2(n_18),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_813),
.A2(n_399),
.B1(n_398),
.B2(n_395),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_801),
.Y(n_872)
);

INVx8_ASAP7_75t_L g873 ( 
.A(n_816),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_805),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_801),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_820),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_806),
.Y(n_877)
);

BUFx4f_ASAP7_75t_SL g878 ( 
.A(n_827),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_818),
.Y(n_879)
);

BUFx2_ASAP7_75t_SL g880 ( 
.A(n_781),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_SL g881 ( 
.A1(n_787),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_819),
.Y(n_882)
);

OAI22xp33_ASAP7_75t_L g883 ( 
.A1(n_775),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_820),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_784),
.Y(n_885)
);

BUFx2_ASAP7_75t_R g886 ( 
.A(n_844),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_856),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_856),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_863),
.Y(n_889)
);

INVx3_ASAP7_75t_SL g890 ( 
.A(n_877),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_878),
.A2(n_775),
.B1(n_780),
.B2(n_796),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_872),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_866),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_869),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_875),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_874),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_874),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_885),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_885),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_867),
.B(n_776),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_885),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_830),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_885),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_879),
.B(n_793),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_864),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_836),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_837),
.Y(n_907)
);

AND2x4_ASAP7_75t_SL g908 ( 
.A(n_868),
.B(n_799),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_868),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_873),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_880),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_873),
.Y(n_912)
);

OA21x2_ASAP7_75t_L g913 ( 
.A1(n_876),
.A2(n_776),
.B(n_780),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_846),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_873),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_884),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_878),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_829),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_829),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_883),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_883),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_870),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_870),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_891),
.A2(n_845),
.B(n_881),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_889),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_900),
.B(n_862),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_902),
.Y(n_927)
);

AOI211xp5_ASAP7_75t_L g928 ( 
.A1(n_920),
.A2(n_853),
.B(n_774),
.C(n_794),
.Y(n_928)
);

INVx4_ASAP7_75t_SL g929 ( 
.A(n_890),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_920),
.A2(n_882),
.B1(n_834),
.B2(n_865),
.Y(n_930)
);

NOR2x1_ASAP7_75t_SL g931 ( 
.A(n_911),
.B(n_848),
.Y(n_931)
);

AOI221xp5_ASAP7_75t_L g932 ( 
.A1(n_922),
.A2(n_861),
.B1(n_859),
.B2(n_839),
.C(n_845),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_886),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_898),
.Y(n_934)
);

AOI221xp5_ASAP7_75t_L g935 ( 
.A1(n_922),
.A2(n_839),
.B1(n_834),
.B2(n_853),
.C(n_840),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_898),
.Y(n_936)
);

AOI221xp5_ASAP7_75t_L g937 ( 
.A1(n_922),
.A2(n_923),
.B1(n_921),
.B2(n_920),
.C(n_891),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_900),
.B(n_854),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_889),
.Y(n_939)
);

OA21x2_ASAP7_75t_L g940 ( 
.A1(n_889),
.A2(n_783),
.B(n_790),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_923),
.A2(n_843),
.B(n_847),
.Y(n_941)
);

INVxp33_ASAP7_75t_L g942 ( 
.A(n_917),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_910),
.B(n_858),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_892),
.Y(n_944)
);

AO32x2_ASAP7_75t_L g945 ( 
.A1(n_902),
.A2(n_850),
.A3(n_828),
.B1(n_860),
.B2(n_855),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_892),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_914),
.B(n_860),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_890),
.B(n_835),
.Y(n_948)
);

AO21x1_ASAP7_75t_L g949 ( 
.A1(n_923),
.A2(n_850),
.B(n_842),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_900),
.B(n_860),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_906),
.B(n_858),
.Y(n_951)
);

AO21x1_ASAP7_75t_L g952 ( 
.A1(n_921),
.A2(n_842),
.B(n_857),
.Y(n_952)
);

AO21x2_ASAP7_75t_L g953 ( 
.A1(n_911),
.A2(n_892),
.B(n_921),
.Y(n_953)
);

OAI22xp33_ASAP7_75t_L g954 ( 
.A1(n_890),
.A2(n_833),
.B1(n_828),
.B2(n_851),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_898),
.Y(n_955)
);

AO21x2_ASAP7_75t_L g956 ( 
.A1(n_911),
.A2(n_796),
.B(n_797),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_917),
.A2(n_843),
.B(n_817),
.C(n_849),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_890),
.B(n_832),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_910),
.B(n_831),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_906),
.B(n_851),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_887),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_895),
.B(n_831),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_906),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_925),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_926),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_926),
.B(n_914),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_925),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_939),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_939),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_944),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_934),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_944),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_946),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_946),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_934),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_927),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_948),
.B(n_954),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_963),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_953),
.B(n_895),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_963),
.B(n_916),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_953),
.B(n_895),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_961),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_950),
.B(n_905),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_961),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_950),
.B(n_905),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_953),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_959),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_962),
.Y(n_988)
);

OAI33xp33_ASAP7_75t_L g989 ( 
.A1(n_986),
.A2(n_947),
.A3(n_907),
.B1(n_933),
.B2(n_962),
.B3(n_916),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_964),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_976),
.B(n_938),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_965),
.B(n_938),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_964),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_R g994 ( 
.A(n_977),
.B(n_933),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_964),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_966),
.A2(n_924),
.B1(n_930),
.B2(n_935),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_971),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_965),
.B(n_987),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_987),
.B(n_934),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_988),
.B(n_936),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_968),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_983),
.B(n_958),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_971),
.Y(n_1003)
);

NAND4xp25_ASAP7_75t_SL g1004 ( 
.A(n_979),
.B(n_930),
.C(n_932),
.D(n_928),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_978),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_988),
.B(n_917),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_968),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_987),
.B(n_936),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_975),
.B(n_936),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_991),
.B(n_985),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_997),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_998),
.B(n_975),
.Y(n_1012)
);

NOR2x1_ASAP7_75t_L g1013 ( 
.A(n_1004),
.B(n_979),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_998),
.B(n_942),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_991),
.B(n_981),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_992),
.B(n_981),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_992),
.B(n_929),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1005),
.B(n_967),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_999),
.B(n_929),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_1000),
.B(n_968),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_1020),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1013),
.B(n_1019),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1013),
.B(n_1019),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_1015),
.B(n_1000),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_1011),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1010),
.B(n_1006),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1018),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_1026),
.B(n_1002),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_1021),
.B(n_1016),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1025),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_1022),
.A2(n_1004),
.B1(n_996),
.B2(n_989),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1030),
.B(n_1022),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_1029),
.B(n_1025),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1028),
.B(n_1023),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1031),
.B(n_1023),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1030),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1028),
.B(n_1027),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1028),
.B(n_1021),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1030),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1028),
.B(n_1024),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1031),
.A2(n_996),
.B1(n_989),
.B2(n_1006),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_1030),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_1033),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_1041),
.A2(n_1035),
.B1(n_1032),
.B2(n_1034),
.Y(n_1044)
);

AOI21xp33_ASAP7_75t_SL g1045 ( 
.A1(n_1038),
.A2(n_886),
.B(n_994),
.Y(n_1045)
);

INVxp33_ASAP7_75t_L g1046 ( 
.A(n_1040),
.Y(n_1046)
);

AOI32xp33_ASAP7_75t_L g1047 ( 
.A1(n_1042),
.A2(n_1017),
.A3(n_1012),
.B1(n_928),
.B2(n_1014),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1036),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1039),
.Y(n_1049)
);

AOI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_1042),
.A2(n_1024),
.B(n_915),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1037),
.A2(n_918),
.B1(n_919),
.B2(n_1003),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1041),
.A2(n_937),
.B1(n_929),
.B2(n_949),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1041),
.A2(n_918),
.B1(n_919),
.B2(n_1003),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_SL g1054 ( 
.A(n_1035),
.B(n_997),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_1041),
.A2(n_918),
.B1(n_919),
.B2(n_1018),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_1034),
.B(n_918),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1041),
.A2(n_919),
.B1(n_986),
.B2(n_957),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_SL g1058 ( 
.A(n_1033),
.B(n_912),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1043),
.B(n_1009),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1046),
.B(n_999),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1048),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_1054),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_1053),
.A2(n_941),
.B(n_952),
.C(n_949),
.Y(n_1063)
);

OAI31xp33_ASAP7_75t_L g1064 ( 
.A1(n_1057),
.A2(n_912),
.A3(n_915),
.B(n_1008),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_1049),
.Y(n_1065)
);

XNOR2xp5_ASAP7_75t_L g1066 ( 
.A(n_1044),
.B(n_943),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1047),
.B(n_1009),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1056),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1051),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1058),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_1055),
.B(n_1050),
.Y(n_1071)
);

AOI221xp5_ASAP7_75t_L g1072 ( 
.A1(n_1052),
.A2(n_952),
.B1(n_1007),
.B2(n_1001),
.C(n_990),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1045),
.B(n_1008),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1043),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_1043),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1043),
.B(n_995),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1043),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1074),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1075),
.B(n_995),
.Y(n_1079)
);

O2A1O1Ixp5_ASAP7_75t_L g1080 ( 
.A1(n_1070),
.A2(n_993),
.B(n_1007),
.C(n_1001),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1062),
.A2(n_929),
.B1(n_959),
.B2(n_943),
.Y(n_1081)
);

AOI211xp5_ASAP7_75t_L g1082 ( 
.A1(n_1077),
.A2(n_915),
.B(n_912),
.C(n_27),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1068),
.B(n_995),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1064),
.B(n_943),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_1069),
.B(n_1005),
.Y(n_1085)
);

AOI222xp33_ASAP7_75t_L g1086 ( 
.A1(n_1072),
.A2(n_931),
.B1(n_960),
.B2(n_907),
.C1(n_990),
.C2(n_29),
.Y(n_1086)
);

NAND4xp75_ASAP7_75t_L g1087 ( 
.A(n_1065),
.B(n_25),
.C(n_26),
.D(n_27),
.Y(n_1087)
);

AOI211xp5_ASAP7_75t_SL g1088 ( 
.A1(n_1073),
.A2(n_841),
.B(n_910),
.C(n_30),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_1060),
.Y(n_1089)
);

OAI211xp5_ASAP7_75t_SL g1090 ( 
.A1(n_1061),
.A2(n_26),
.B(n_28),
.C(n_31),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_1060),
.B(n_943),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_1073),
.B(n_28),
.Y(n_1092)
);

AND3x1_ASAP7_75t_L g1093 ( 
.A(n_1061),
.B(n_995),
.C(n_960),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_L g1094 ( 
.A(n_1071),
.B(n_32),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_SL g1095 ( 
.A1(n_1088),
.A2(n_1066),
.B(n_1071),
.Y(n_1095)
);

AOI21xp33_ASAP7_75t_R g1096 ( 
.A1(n_1078),
.A2(n_1067),
.B(n_1059),
.Y(n_1096)
);

AOI221x1_ASAP7_75t_L g1097 ( 
.A1(n_1092),
.A2(n_1076),
.B1(n_1065),
.B2(n_1063),
.C(n_993),
.Y(n_1097)
);

OAI211xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1094),
.A2(n_32),
.B(n_34),
.C(n_35),
.Y(n_1098)
);

AOI211xp5_ASAP7_75t_L g1099 ( 
.A1(n_1090),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_1099)
);

AOI211xp5_ASAP7_75t_SL g1100 ( 
.A1(n_1085),
.A2(n_841),
.B(n_38),
.C(n_39),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_L g1101 ( 
.A(n_1089),
.B(n_1090),
.C(n_1082),
.Y(n_1101)
);

AOI221xp5_ASAP7_75t_L g1102 ( 
.A1(n_1079),
.A2(n_993),
.B1(n_907),
.B2(n_982),
.C(n_972),
.Y(n_1102)
);

NOR4xp75_ASAP7_75t_L g1103 ( 
.A(n_1083),
.B(n_36),
.C(n_40),
.D(n_41),
.Y(n_1103)
);

AND4x1_ASAP7_75t_L g1104 ( 
.A(n_1081),
.B(n_40),
.C(n_41),
.D(n_42),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1093),
.A2(n_982),
.B1(n_967),
.B2(n_972),
.Y(n_1105)
);

AOI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_1086),
.A2(n_45),
.B(n_47),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1084),
.A2(n_959),
.B1(n_910),
.B2(n_956),
.Y(n_1107)
);

OAI221xp5_ASAP7_75t_L g1108 ( 
.A1(n_1091),
.A2(n_910),
.B1(n_838),
.B2(n_905),
.C(n_974),
.Y(n_1108)
);

AOI221xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1087),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.C(n_52),
.Y(n_1109)
);

XNOR2x1_ASAP7_75t_L g1110 ( 
.A(n_1080),
.B(n_50),
.Y(n_1110)
);

NOR4xp25_ASAP7_75t_L g1111 ( 
.A(n_1078),
.B(n_51),
.C(n_52),
.D(n_53),
.Y(n_1111)
);

AOI221x1_ASAP7_75t_L g1112 ( 
.A1(n_1078),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.C(n_58),
.Y(n_1112)
);

AOI222xp33_ASAP7_75t_L g1113 ( 
.A1(n_1094),
.A2(n_931),
.B1(n_58),
.B2(n_54),
.C1(n_908),
.C2(n_945),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1081),
.A2(n_974),
.B1(n_984),
.B2(n_973),
.Y(n_1114)
);

OAI211xp5_ASAP7_75t_L g1115 ( 
.A1(n_1094),
.A2(n_849),
.B(n_831),
.C(n_910),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_1092),
.A2(n_916),
.B1(n_951),
.B2(n_956),
.C(n_959),
.Y(n_1116)
);

OAI221xp5_ASAP7_75t_SL g1117 ( 
.A1(n_1081),
.A2(n_951),
.B1(n_980),
.B2(n_945),
.C(n_973),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1089),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1118),
.Y(n_1119)
);

AOI21xp33_ASAP7_75t_SL g1120 ( 
.A1(n_1101),
.A2(n_849),
.B(n_63),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1100),
.B(n_978),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1110),
.Y(n_1122)
);

AOI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_1095),
.A2(n_1115),
.B(n_1106),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1104),
.B(n_978),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1107),
.A2(n_984),
.B1(n_969),
.B2(n_973),
.Y(n_1125)
);

OAI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1112),
.A2(n_984),
.B1(n_970),
.B2(n_969),
.Y(n_1126)
);

NOR3xp33_ASAP7_75t_L g1127 ( 
.A(n_1098),
.B(n_819),
.C(n_905),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1111),
.B(n_980),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1099),
.A2(n_956),
.B(n_969),
.C(n_970),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1108),
.A2(n_970),
.B1(n_955),
.B2(n_838),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1109),
.A2(n_908),
.B(n_955),
.C(n_898),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1113),
.A2(n_838),
.B1(n_852),
.B2(n_955),
.Y(n_1132)
);

AOI221xp5_ASAP7_75t_L g1133 ( 
.A1(n_1096),
.A2(n_1114),
.B1(n_1116),
.B2(n_1117),
.C(n_1105),
.Y(n_1133)
);

XOR2x1_ASAP7_75t_L g1134 ( 
.A(n_1103),
.B(n_61),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_SL g1135 ( 
.A(n_1113),
.B(n_871),
.C(n_815),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1097),
.B(n_831),
.Y(n_1136)
);

AOI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_1102),
.A2(n_903),
.B1(n_899),
.B2(n_901),
.C(n_908),
.Y(n_1137)
);

AOI222xp33_ASAP7_75t_L g1138 ( 
.A1(n_1095),
.A2(n_908),
.B1(n_945),
.B2(n_904),
.C1(n_852),
.C2(n_893),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_SL g1139 ( 
.A(n_1101),
.B(n_871),
.C(n_903),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1101),
.A2(n_852),
.B1(n_899),
.B2(n_903),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_L g1141 ( 
.A1(n_1096),
.A2(n_901),
.B1(n_899),
.B2(n_903),
.C(n_893),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1118),
.B(n_899),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1119),
.B(n_901),
.Y(n_1143)
);

NAND2xp33_ASAP7_75t_L g1144 ( 
.A(n_1122),
.B(n_384),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1124),
.B(n_901),
.Y(n_1145)
);

INVxp33_ASAP7_75t_SL g1146 ( 
.A(n_1120),
.Y(n_1146)
);

NAND2x1p5_ASAP7_75t_L g1147 ( 
.A(n_1121),
.B(n_384),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1134),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1136),
.Y(n_1149)
);

OAI322xp33_ASAP7_75t_L g1150 ( 
.A1(n_1128),
.A2(n_1142),
.A3(n_1140),
.B1(n_1129),
.B2(n_1132),
.C1(n_1126),
.C2(n_1130),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_1125),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1139),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1131),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1123),
.B(n_384),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1133),
.B(n_384),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1141),
.B(n_945),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1135),
.A2(n_1138),
.B1(n_1127),
.B2(n_1137),
.Y(n_1157)
);

NAND4xp75_ASAP7_75t_L g1158 ( 
.A(n_1123),
.B(n_913),
.C(n_68),
.D(n_69),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1119),
.Y(n_1159)
);

NOR2x1_ASAP7_75t_L g1160 ( 
.A(n_1122),
.B(n_384),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1122),
.B(n_913),
.Y(n_1161)
);

NAND4xp75_ASAP7_75t_L g1162 ( 
.A(n_1123),
.B(n_913),
.C(n_71),
.D(n_72),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1119),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1119),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1148),
.B(n_66),
.Y(n_1165)
);

NOR3xp33_ASAP7_75t_L g1166 ( 
.A(n_1159),
.B(n_74),
.C(n_78),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1163),
.B(n_79),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_1164),
.B(n_384),
.C(n_389),
.Y(n_1168)
);

AOI322xp5_ASAP7_75t_L g1169 ( 
.A1(n_1153),
.A2(n_945),
.A3(n_894),
.B1(n_887),
.B2(n_909),
.C1(n_904),
.C2(n_897),
.Y(n_1169)
);

OAI221xp5_ASAP7_75t_L g1170 ( 
.A1(n_1151),
.A2(n_909),
.B1(n_897),
.B2(n_896),
.C(n_913),
.Y(n_1170)
);

AOI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1146),
.A2(n_909),
.B1(n_904),
.B2(n_894),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1149),
.B(n_909),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_L g1173 ( 
.A(n_1152),
.B(n_80),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1144),
.B(n_384),
.C(n_389),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1147),
.A2(n_1155),
.B1(n_1160),
.B2(n_1154),
.Y(n_1175)
);

NOR3xp33_ASAP7_75t_L g1176 ( 
.A(n_1150),
.B(n_83),
.C(n_87),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1143),
.B(n_896),
.Y(n_1177)
);

AOI32xp33_ASAP7_75t_L g1178 ( 
.A1(n_1145),
.A2(n_894),
.A3(n_904),
.B1(n_887),
.B2(n_897),
.Y(n_1178)
);

NOR3xp33_ASAP7_75t_L g1179 ( 
.A(n_1158),
.B(n_90),
.C(n_91),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1165),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_1167),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1176),
.B(n_1143),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1179),
.A2(n_1162),
.B1(n_1145),
.B2(n_1157),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1173),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1166),
.B(n_1168),
.C(n_1174),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1172),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1175),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_SL g1188 ( 
.A1(n_1170),
.A2(n_1161),
.B1(n_1156),
.B2(n_897),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1171),
.A2(n_904),
.B1(n_913),
.B2(n_940),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1177),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1178),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1169),
.A2(n_896),
.B1(n_888),
.B2(n_904),
.Y(n_1192)
);

XNOR2x1_ASAP7_75t_L g1193 ( 
.A(n_1165),
.B(n_93),
.Y(n_1193)
);

XNOR2x1_ASAP7_75t_L g1194 ( 
.A(n_1165),
.B(n_94),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1184),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1193),
.A2(n_888),
.B1(n_896),
.B2(n_102),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1187),
.A2(n_913),
.B1(n_940),
.B2(n_888),
.Y(n_1197)
);

AO22x2_ASAP7_75t_L g1198 ( 
.A1(n_1194),
.A2(n_888),
.B1(n_101),
.B2(n_104),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1183),
.A2(n_940),
.B1(n_399),
.B2(n_398),
.Y(n_1199)
);

AOI31xp33_ASAP7_75t_L g1200 ( 
.A1(n_1180),
.A2(n_96),
.A3(n_105),
.B(n_106),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1191),
.A2(n_1181),
.B1(n_1190),
.B2(n_1185),
.Y(n_1201)
);

INVxp67_ASAP7_75t_SL g1202 ( 
.A(n_1186),
.Y(n_1202)
);

AO22x2_ASAP7_75t_L g1203 ( 
.A1(n_1186),
.A2(n_108),
.B1(n_110),
.B2(n_113),
.Y(n_1203)
);

OAI22x1_ASAP7_75t_L g1204 ( 
.A1(n_1182),
.A2(n_940),
.B1(n_116),
.B2(n_117),
.Y(n_1204)
);

OAI22x1_ASAP7_75t_L g1205 ( 
.A1(n_1202),
.A2(n_1189),
.B1(n_1188),
.B2(n_1192),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1195),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1201),
.Y(n_1207)
);

INVxp67_ASAP7_75t_SL g1208 ( 
.A(n_1198),
.Y(n_1208)
);

AO22x2_ASAP7_75t_L g1209 ( 
.A1(n_1199),
.A2(n_114),
.B1(n_119),
.B2(n_120),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1203),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1210),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1207),
.A2(n_1208),
.B1(n_1206),
.B2(n_1205),
.Y(n_1212)
);

XNOR2xp5_ASAP7_75t_L g1213 ( 
.A(n_1209),
.B(n_1196),
.Y(n_1213)
);

OAI22x1_ASAP7_75t_L g1214 ( 
.A1(n_1209),
.A2(n_1200),
.B1(n_1204),
.B2(n_1197),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1211),
.A2(n_1214),
.B1(n_1212),
.B2(n_1213),
.Y(n_1215)
);

AO21x2_ASAP7_75t_L g1216 ( 
.A1(n_1215),
.A2(n_123),
.B(n_126),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1216),
.A2(n_128),
.B(n_129),
.Y(n_1217)
);

OAI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1217),
.A2(n_399),
.B1(n_398),
.B2(n_395),
.Y(n_1218)
);

AOI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1218),
.A2(n_399),
.B1(n_398),
.B2(n_395),
.C(n_389),
.Y(n_1219)
);

AOI211xp5_ASAP7_75t_L g1220 ( 
.A1(n_1219),
.A2(n_399),
.B(n_398),
.C(n_395),
.Y(n_1220)
);


endmodule