module fake_jpeg_1979_n_427 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_427);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_427;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx8_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g126 ( 
.A(n_61),
.Y(n_126)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_68),
.B(n_70),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_18),
.B(n_0),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_72),
.B(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_17),
.B(n_2),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_83),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_18),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_77),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_79),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_80),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_81),
.Y(n_138)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_82),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_85),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_87),
.B(n_88),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_17),
.B(n_2),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_89),
.B(n_90),
.Y(n_151)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_91),
.B(n_92),
.Y(n_152)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx16f_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_21),
.B(n_2),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

CKINVDCx12_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_21),
.B(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_98),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_44),
.B1(n_31),
.B2(n_32),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_102),
.A2(n_140),
.B1(n_146),
.B2(n_150),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_28),
.B1(n_43),
.B2(n_39),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_105),
.A2(n_129),
.B1(n_136),
.B2(n_153),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_36),
.C(n_43),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_112),
.B(n_10),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_50),
.A2(n_44),
.B1(n_34),
.B2(n_32),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_116),
.A2(n_13),
.B1(n_123),
.B2(n_138),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_36),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_134),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_39),
.B1(n_31),
.B2(n_34),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_53),
.B(n_4),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_55),
.B(n_59),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_147),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_33),
.B1(n_27),
.B2(n_24),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_57),
.A2(n_42),
.B1(n_33),
.B2(n_27),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_61),
.A2(n_42),
.B1(n_33),
.B2(n_27),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_65),
.B(n_4),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_69),
.A2(n_81),
.B1(n_77),
.B2(n_79),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_86),
.A2(n_24),
.B1(n_15),
.B2(n_6),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_76),
.A2(n_24),
.B1(n_15),
.B2(n_6),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_112),
.B1(n_126),
.B2(n_137),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_74),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_156),
.B(n_178),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_94),
.B1(n_93),
.B2(n_98),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_158),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_100),
.B(n_83),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_162),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_113),
.A2(n_15),
.B(n_5),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_165),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_80),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_182),
.Y(n_202)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_167),
.A2(n_174),
.B1(n_195),
.B2(n_133),
.Y(n_209)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_181),
.B1(n_187),
.B2(n_189),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_172),
.Y(n_228)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_176),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_116),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_134),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_175),
.A2(n_177),
.B1(n_194),
.B2(n_141),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_115),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_180),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_SL g180 ( 
.A(n_130),
.B(n_12),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_117),
.B(n_13),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_186),
.Y(n_223)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_117),
.A2(n_149),
.B1(n_110),
.B2(n_131),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_192),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_147),
.A2(n_135),
.B1(n_126),
.B2(n_142),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_104),
.A2(n_101),
.B1(n_106),
.B2(n_141),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_126),
.A3(n_144),
.B1(n_104),
.B2(n_114),
.Y(n_212)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_196),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_137),
.A2(n_103),
.B1(n_132),
.B2(n_122),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_145),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_198),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_118),
.B(n_127),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_128),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_137),
.A2(n_103),
.B1(n_122),
.B2(n_132),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_99),
.B1(n_158),
.B2(n_181),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_212),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_139),
.C(n_107),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_208),
.C(n_165),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_142),
.C(n_144),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_211),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_143),
.B(n_121),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_185),
.B(n_197),
.Y(n_251)
);

AOI32xp33_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_121),
.A3(n_108),
.B1(n_99),
.B2(n_139),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_229),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_108),
.B1(n_114),
.B2(n_120),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_159),
.A2(n_157),
.B1(n_182),
.B2(n_161),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_163),
.A2(n_184),
.B1(n_162),
.B2(n_199),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_208),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_194),
.A2(n_160),
.B1(n_186),
.B2(n_164),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_176),
.B(n_175),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_193),
.B(n_179),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_215),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_191),
.A2(n_183),
.B1(n_168),
.B2(n_173),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_235),
.A2(n_196),
.B(n_191),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_206),
.A2(n_191),
.B1(n_198),
.B2(n_192),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_254),
.B1(n_220),
.B2(n_251),
.Y(n_270)
);

BUFx2_ASAP7_75t_SL g239 ( 
.A(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_221),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_247),
.Y(n_267)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_243),
.A2(n_252),
.B(n_214),
.Y(n_286)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_245),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_248),
.Y(n_288)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_251),
.A2(n_235),
.B(n_214),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_222),
.A2(n_170),
.B(n_167),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_258),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_206),
.A2(n_169),
.B1(n_172),
.B2(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_205),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

BUFx8_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_262),
.Y(n_273)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_202),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_283),
.C(n_285),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_263),
.B1(n_244),
.B2(n_237),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_202),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_275),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_215),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_215),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_279),
.Y(n_312)
);

AOI21xp33_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_217),
.B(n_236),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_278),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_262),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_229),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_218),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_207),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_284),
.A2(n_286),
.B(n_243),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_208),
.C(n_204),
.Y(n_285)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_294),
.Y(n_317)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_238),
.C(n_252),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_300),
.C(n_301),
.Y(n_334)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_267),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_302),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_238),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_230),
.C(n_224),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_267),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_303),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_217),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_309),
.C(n_311),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_265),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_306),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_276),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_307),
.A2(n_286),
.B(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_244),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_310),
.A2(n_210),
.B1(n_249),
.B2(n_259),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_274),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_230),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_268),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_277),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_332),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_312),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_324),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_270),
.B1(n_268),
.B2(n_271),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_319),
.A2(n_328),
.B1(n_333),
.B2(n_336),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_271),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_320),
.B(n_325),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_302),
.B(n_276),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_322),
.B(n_330),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_246),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_292),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_307),
.A2(n_249),
.B(n_284),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_293),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_291),
.A2(n_259),
.B1(n_254),
.B2(n_284),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_291),
.A2(n_211),
.B1(n_289),
.B2(n_279),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_292),
.B(n_272),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_337),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_316),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_343),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_293),
.C(n_296),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_355),
.C(n_357),
.Y(n_363)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_342),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_294),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_345),
.Y(n_372)
);

OA22x2_ASAP7_75t_L g345 ( 
.A1(n_319),
.A2(n_295),
.B1(n_297),
.B2(n_303),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_321),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_347),
.A2(n_348),
.B1(n_349),
.B2(n_354),
.Y(n_359)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_312),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_350),
.Y(n_365)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_331),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_301),
.C(n_300),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_289),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_313),
.C(n_311),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_335),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_361),
.C(n_362),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_335),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_357),
.B(n_324),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_346),
.A2(n_323),
.B1(n_317),
.B2(n_327),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_364),
.A2(n_347),
.B1(n_340),
.B2(n_333),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_341),
.B(n_315),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_366),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_322),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_367),
.A2(n_368),
.B(n_370),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_342),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_338),
.B(n_299),
.Y(n_369)
);

NOR3xp33_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_354),
.C(n_349),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_327),
.C(n_323),
.Y(n_370)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_373),
.Y(n_380)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_374),
.Y(n_389)
);

OAI221xp5_ASAP7_75t_L g376 ( 
.A1(n_358),
.A2(n_351),
.B1(n_343),
.B2(n_329),
.C(n_350),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_376),
.A2(n_336),
.B1(n_308),
.B2(n_345),
.Y(n_394)
);

OAI322xp33_ASAP7_75t_L g377 ( 
.A1(n_365),
.A2(n_299),
.A3(n_344),
.B1(n_236),
.B2(n_314),
.C1(n_348),
.C2(n_356),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_381),
.Y(n_388)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_362),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_379),
.B(n_361),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_359),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_330),
.B(n_352),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_384),
.Y(n_393)
);

AO21x1_ASAP7_75t_L g384 ( 
.A1(n_371),
.A2(n_352),
.B(n_345),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_386),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_378),
.A2(n_363),
.B(n_370),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_387),
.A2(n_262),
.B(n_266),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_384),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_390),
.A2(n_398),
.B1(n_273),
.B2(n_383),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_360),
.Y(n_392)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

OAI21xp33_ASAP7_75t_SL g404 ( 
.A1(n_394),
.A2(n_266),
.B(n_248),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_380),
.A2(n_345),
.B(n_363),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_395),
.A2(n_287),
.B(n_228),
.Y(n_405)
);

NAND5xp2_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_223),
.C(n_234),
.D(n_218),
.E(n_256),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_383),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_397),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_375),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_399),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_395),
.B(n_366),
.C(n_273),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_400),
.B(n_407),
.Y(n_410)
);

FAx1_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_262),
.CI(n_272),
.CON(n_401),
.SN(n_401)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_401),
.A2(n_403),
.B(n_405),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_393),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_287),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_408),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_406),
.B(n_391),
.C(n_389),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_412),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_393),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_415),
.A2(n_255),
.B(n_250),
.Y(n_418)
);

NAND4xp25_ASAP7_75t_SL g416 ( 
.A(n_414),
.B(n_406),
.C(n_390),
.D(n_405),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_420),
.C(n_412),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_418),
.A2(n_419),
.B(n_417),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_410),
.A2(n_287),
.B(n_245),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_264),
.Y(n_420)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_421),
.A2(n_423),
.B(n_225),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_417),
.A2(n_411),
.B(n_413),
.Y(n_422)
);

AOI322xp5_ASAP7_75t_L g424 ( 
.A1(n_422),
.A2(n_223),
.A3(n_260),
.B1(n_227),
.B2(n_216),
.C1(n_212),
.C2(n_225),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_424),
.B(n_425),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_426),
.B(n_201),
.Y(n_427)
);


endmodule