module fake_aes_8592_n_1122 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1122);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1122;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_383;
wire n_288;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_236;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_1042;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_560;
wire n_517;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_1101;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_230;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_828;
wire n_767;
wire n_1063;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_1066;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_429;
wire n_488;
wire n_233;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_1069;
wire n_1021;
wire n_972;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_947;
wire n_1043;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
INVx2_ASAP7_75t_L g230 ( .A(n_139), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_165), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_112), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_157), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_65), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_179), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_45), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_202), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_35), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_25), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_96), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_79), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_64), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_21), .Y(n_243) );
INVx2_ASAP7_75t_SL g244 ( .A(n_71), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_155), .Y(n_245) );
INVxp67_ASAP7_75t_L g246 ( .A(n_135), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_42), .Y(n_247) );
INVxp67_ASAP7_75t_SL g248 ( .A(n_75), .Y(n_248) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_59), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_197), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_125), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_111), .Y(n_252) );
INVxp67_ASAP7_75t_L g253 ( .A(n_1), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_153), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_118), .Y(n_255) );
BUFx2_ASAP7_75t_SL g256 ( .A(n_93), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_191), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_98), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_208), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_46), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_211), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_29), .B(n_146), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_82), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_158), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_210), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_204), .Y(n_266) );
CKINVDCx14_ASAP7_75t_R g267 ( .A(n_218), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_156), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_194), .Y(n_269) );
BUFx10_ASAP7_75t_L g270 ( .A(n_121), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_29), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_198), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_7), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_33), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_89), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_51), .Y(n_276) );
CKINVDCx16_ASAP7_75t_R g277 ( .A(n_175), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_97), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_168), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_36), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_131), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_174), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_35), .Y(n_283) );
CKINVDCx16_ASAP7_75t_R g284 ( .A(n_10), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_101), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_115), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_201), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_167), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_13), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_7), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_17), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_32), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_176), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_196), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_85), .Y(n_295) );
CKINVDCx14_ASAP7_75t_R g296 ( .A(n_51), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_219), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_181), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_9), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_10), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_187), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_190), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_23), .Y(n_303) );
INVxp33_ASAP7_75t_SL g304 ( .A(n_22), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_164), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_162), .Y(n_306) );
CKINVDCx16_ASAP7_75t_R g307 ( .A(n_76), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_40), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_43), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_110), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_32), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_1), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_108), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_12), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_106), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_57), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_105), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_19), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_50), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_130), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_171), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_132), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_13), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_47), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_26), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_28), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_77), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_37), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_213), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_91), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_163), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_169), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_8), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_47), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_147), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_229), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_87), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_60), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_136), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_113), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_53), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_78), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_49), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_212), .Y(n_344) );
BUFx5_ASAP7_75t_L g345 ( .A(n_126), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_225), .Y(n_346) );
INVxp67_ASAP7_75t_SL g347 ( .A(n_9), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_144), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_95), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_224), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_296), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_255), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_292), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_292), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_240), .Y(n_355) );
OAI22xp5_ASAP7_75t_SL g356 ( .A1(n_343), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_273), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_345), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_236), .B(n_0), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_296), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_345), .Y(n_361) );
OAI22xp5_ASAP7_75t_SL g362 ( .A1(n_343), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_244), .B(n_4), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_286), .B(n_5), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_274), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_327), .B(n_5), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_240), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_234), .B(n_6), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_345), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_273), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_309), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_345), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_309), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_345), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_242), .A2(n_6), .B1(n_8), .B2(n_11), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_240), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_270), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_311), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_311), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_333), .B(n_12), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_333), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_345), .Y(n_382) );
INVx3_ASAP7_75t_L g383 ( .A(n_270), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_238), .B(n_14), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_380), .Y(n_385) );
INVx6_ASAP7_75t_L g386 ( .A(n_380), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_377), .B(n_235), .Y(n_387) );
OR2x6_ASAP7_75t_L g388 ( .A(n_356), .B(n_256), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_380), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_358), .Y(n_390) );
BUFx4f_ASAP7_75t_L g391 ( .A(n_377), .Y(n_391) );
INVx4_ASAP7_75t_L g392 ( .A(n_377), .Y(n_392) );
INVx4_ASAP7_75t_L g393 ( .A(n_383), .Y(n_393) );
INVx2_ASAP7_75t_SL g394 ( .A(n_351), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_358), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_351), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_360), .B(n_277), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_360), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_358), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_361), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_383), .B(n_246), .Y(n_403) );
NAND2xp33_ASAP7_75t_L g404 ( .A(n_361), .B(n_345), .Y(n_404) );
BUFx10_ASAP7_75t_L g405 ( .A(n_365), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_355), .Y(n_406) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_355), .Y(n_407) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_366), .B(n_253), .C(n_274), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_383), .B(n_307), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_356), .Y(n_410) );
BUFx4f_ASAP7_75t_L g411 ( .A(n_383), .Y(n_411) );
INVx5_ASAP7_75t_L g412 ( .A(n_355), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_371), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_369), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_379), .B(n_270), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_379), .B(n_254), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_369), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_369), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_352), .B(n_364), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_372), .Y(n_420) );
XNOR2xp5_ASAP7_75t_L g421 ( .A(n_362), .B(n_304), .Y(n_421) );
BUFx4f_ASAP7_75t_L g422 ( .A(n_357), .Y(n_422) );
BUFx10_ASAP7_75t_L g423 ( .A(n_357), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_352), .B(n_290), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_364), .B(n_243), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_366), .A2(n_247), .B1(n_276), .B2(n_271), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_355), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_372), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_372), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_374), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_392), .Y(n_431) );
INVxp67_ASAP7_75t_L g432 ( .A(n_413), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_392), .Y(n_433) );
NAND3xp33_ASAP7_75t_SL g434 ( .A(n_399), .B(n_257), .C(n_252), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_399), .Y(n_435) );
OR2x2_ASAP7_75t_SL g436 ( .A(n_421), .B(n_249), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_419), .B(n_352), .Y(n_437) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_388), .A2(n_375), .B1(n_284), .B2(n_359), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_405), .B(n_290), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_388), .A2(n_362), .B1(n_375), .B2(n_304), .Y(n_440) );
OAI22xp33_ASAP7_75t_L g441 ( .A1(n_388), .A2(n_252), .B1(n_275), .B2(n_257), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_394), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_393), .B(n_363), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_393), .B(n_363), .Y(n_444) );
BUFx2_ASAP7_75t_SL g445 ( .A(n_405), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_405), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_393), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_387), .B(n_370), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_385), .B(n_382), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_385), .B(n_382), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_386), .A2(n_373), .B1(n_381), .B2(n_378), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_403), .B(n_373), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_396), .B(n_291), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_386), .A2(n_378), .B1(n_381), .B2(n_368), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_424), .B(n_294), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_396), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_425), .B(n_291), .Y(n_457) );
NAND2x1p5_ASAP7_75t_L g458 ( .A(n_391), .B(n_283), .Y(n_458) );
AND2x2_ASAP7_75t_SL g459 ( .A(n_391), .B(n_262), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_389), .Y(n_460) );
INVx5_ASAP7_75t_L g461 ( .A(n_389), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_389), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_425), .B(n_368), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_423), .B(n_294), .Y(n_464) );
BUFx6f_ASAP7_75t_SL g465 ( .A(n_388), .Y(n_465) );
BUFx3_ASAP7_75t_L g466 ( .A(n_390), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_410), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_408), .A2(n_306), .B1(n_336), .B2(n_288), .Y(n_468) );
NOR2x2_ASAP7_75t_L g469 ( .A(n_421), .B(n_306), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_397), .B(n_312), .Y(n_470) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_423), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_426), .B(n_312), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_411), .B(n_302), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_411), .A2(n_336), .B1(n_384), .B2(n_328), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_411), .B(n_289), .Y(n_475) );
INVx5_ASAP7_75t_L g476 ( .A(n_390), .Y(n_476) );
CKINVDCx11_ASAP7_75t_R g477 ( .A(n_395), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_401), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_416), .B(n_310), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_401), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_409), .B(n_384), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_415), .B(n_299), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_422), .Y(n_483) );
INVx8_ASAP7_75t_L g484 ( .A(n_422), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_417), .B(n_232), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_417), .B(n_310), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_418), .B(n_314), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_418), .B(n_315), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_420), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_420), .A2(n_354), .B1(n_353), .B2(n_300), .Y(n_490) );
OR2x6_ASAP7_75t_L g491 ( .A(n_428), .B(n_316), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_428), .B(n_233), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_430), .B(n_314), .Y(n_493) );
NAND2xp33_ASAP7_75t_L g494 ( .A(n_430), .B(n_315), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_395), .B(n_317), .Y(n_495) );
NAND2xp33_ASAP7_75t_L g496 ( .A(n_400), .B(n_317), .Y(n_496) );
BUFx12f_ASAP7_75t_L g497 ( .A(n_412), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_402), .A2(n_354), .B1(n_353), .B2(n_318), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_404), .A2(n_341), .B1(n_328), .B2(n_239), .Y(n_499) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_414), .B(n_342), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_404), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_414), .B(n_330), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_429), .B(n_267), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_412), .B(n_267), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_412), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_412), .Y(n_506) );
NAND2x1p5_ASAP7_75t_L g507 ( .A(n_412), .B(n_323), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_463), .B(n_341), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_471), .B(n_231), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_438), .A2(n_347), .B1(n_319), .B2(n_248), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_463), .B(n_260), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_471), .B(n_261), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_462), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_487), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_454), .B(n_325), .C(n_324), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_493), .B(n_280), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_481), .B(n_326), .Y(n_517) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_471), .Y(n_518) );
AO21x1_ASAP7_75t_L g519 ( .A1(n_503), .A2(n_245), .B(n_237), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_491), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_471), .B(n_263), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_481), .B(n_334), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_432), .B(n_303), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_489), .Y(n_524) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_454), .B(n_338), .C(n_251), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_491), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_445), .B(n_308), .Y(n_527) );
NAND3xp33_ASAP7_75t_SL g528 ( .A(n_440), .B(n_348), .C(n_279), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_448), .A2(n_258), .B(n_259), .C(n_250), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_446), .B(n_278), .Y(n_530) );
XOR2xp5_ASAP7_75t_L g531 ( .A(n_434), .B(n_14), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_438), .A2(n_266), .B(n_269), .C(n_264), .Y(n_532) );
BUFx2_ASAP7_75t_L g533 ( .A(n_435), .Y(n_533) );
INVx6_ASAP7_75t_L g534 ( .A(n_497), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_439), .B(n_15), .Y(n_535) );
INVx3_ASAP7_75t_SL g536 ( .A(n_469), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_459), .A2(n_282), .B1(n_285), .B2(n_281), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_457), .B(n_15), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_461), .Y(n_539) );
INVx5_ASAP7_75t_L g540 ( .A(n_484), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_456), .B(n_293), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_477), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_459), .A2(n_297), .B1(n_298), .B2(n_295), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_443), .A2(n_305), .B1(n_313), .B2(n_301), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_456), .B(n_320), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_444), .A2(n_332), .B1(n_337), .B2(n_331), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_460), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_464), .B(n_339), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_472), .B(n_16), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_474), .A2(n_344), .B(n_346), .C(n_340), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_442), .B(n_349), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_484), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_478), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_453), .B(n_16), .Y(n_554) );
BUFx3_ASAP7_75t_L g555 ( .A(n_476), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_470), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_458), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_486), .B(n_255), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_488), .B(n_268), .Y(n_559) );
NOR2xp33_ASAP7_75t_R g560 ( .A(n_465), .B(n_18), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_458), .A2(n_241), .B1(n_287), .B2(n_230), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_476), .Y(n_562) );
INVx3_ASAP7_75t_L g563 ( .A(n_466), .Y(n_563) );
BUFx12f_ASAP7_75t_L g564 ( .A(n_436), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_502), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_475), .A2(n_335), .B1(n_350), .B2(n_322), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_475), .Y(n_567) );
OAI22x1_ASAP7_75t_L g568 ( .A1(n_468), .A2(n_350), .B1(n_335), .B2(n_20), .Y(n_568) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_484), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_482), .B(n_18), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_451), .A2(n_321), .B1(n_268), .B2(n_265), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_461), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_451), .A2(n_321), .B1(n_265), .B2(n_272), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_479), .B(n_19), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_452), .A2(n_406), .B(n_398), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_480), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_455), .B(n_20), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_499), .B(n_500), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_440), .A2(n_240), .B1(n_265), .B2(n_272), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_461), .B(n_22), .Y(n_580) );
NOR2xp33_ASAP7_75t_SL g581 ( .A(n_441), .B(n_265), .Y(n_581) );
NAND2xp33_ASAP7_75t_SL g582 ( .A(n_465), .B(n_272), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g583 ( .A1(n_437), .A2(n_272), .B(n_329), .C(n_376), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_467), .Y(n_584) );
INVx3_ASAP7_75t_L g585 ( .A(n_476), .Y(n_585) );
AOI21xp33_ASAP7_75t_L g586 ( .A1(n_494), .A2(n_329), .B(n_24), .Y(n_586) );
OR2x6_ASAP7_75t_L g587 ( .A(n_441), .B(n_329), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_485), .Y(n_588) );
A2O1A1Ixp33_ASAP7_75t_L g589 ( .A1(n_501), .A2(n_329), .B(n_376), .C(n_367), .Y(n_589) );
A2O1A1Ixp33_ASAP7_75t_L g590 ( .A1(n_431), .A2(n_376), .B(n_367), .C(n_355), .Y(n_590) );
CKINVDCx6p67_ASAP7_75t_R g591 ( .A(n_476), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_490), .B(n_24), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_483), .B(n_367), .Y(n_593) );
OAI21xp33_ASAP7_75t_SL g594 ( .A1(n_492), .A2(n_25), .B(n_26), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_495), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_498), .A2(n_367), .B1(n_376), .B2(n_30), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_498), .B(n_376), .C(n_367), .Y(n_597) );
BUFx2_ASAP7_75t_L g598 ( .A(n_507), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_492), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_433), .Y(n_600) );
INVx2_ASAP7_75t_SL g601 ( .A(n_473), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_447), .A2(n_376), .B1(n_28), .B2(n_30), .Y(n_602) );
NOR2xp33_ASAP7_75t_R g603 ( .A(n_496), .B(n_27), .Y(n_603) );
AND2x6_ASAP7_75t_L g604 ( .A(n_505), .B(n_398), .Y(n_604) );
AO22x1_ASAP7_75t_L g605 ( .A1(n_504), .A2(n_27), .B1(n_31), .B2(n_34), .Y(n_605) );
INVx8_ASAP7_75t_L g606 ( .A(n_506), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_463), .B(n_31), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_446), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_432), .B(n_34), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_489), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_432), .B(n_38), .Y(n_611) );
INVx4_ASAP7_75t_L g612 ( .A(n_471), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_432), .B(n_39), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_587), .A2(n_427), .B1(n_407), .B2(n_406), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_SL g615 ( .A1(n_583), .A2(n_123), .B(n_228), .C(n_227), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_600), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_524), .B(n_39), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_587), .A2(n_427), .B1(n_407), .B2(n_42), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_514), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_553), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_575), .A2(n_427), .B(n_407), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_581), .A2(n_427), .B1(n_407), .B2(n_43), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_576), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_SL g624 ( .A1(n_529), .A2(n_590), .B(n_586), .C(n_589), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_542), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_577), .A2(n_427), .B(n_41), .C(n_44), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_558), .A2(n_81), .B(n_80), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_607), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_SL g629 ( .A1(n_578), .A2(n_127), .B(n_223), .C(n_222), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_565), .B(n_537), .Y(n_630) );
NAND2x1_ASAP7_75t_L g631 ( .A(n_612), .B(n_83), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_559), .A2(n_86), .B(n_84), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_548), .A2(n_90), .B(n_88), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_587), .A2(n_40), .B1(n_41), .B2(n_44), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_533), .B(n_45), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_540), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_532), .A2(n_46), .B1(n_48), .B2(n_49), .C(n_50), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_537), .B(n_48), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_SL g639 ( .A1(n_592), .A2(n_141), .B(n_221), .C(n_220), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_556), .B(n_52), .Y(n_640) );
O2A1O1Ixp33_ASAP7_75t_L g641 ( .A1(n_550), .A2(n_52), .B(n_53), .C(n_54), .Y(n_641) );
AO31x2_ASAP7_75t_L g642 ( .A1(n_519), .A2(n_54), .A3(n_55), .B(n_56), .Y(n_642) );
CKINVDCx16_ASAP7_75t_R g643 ( .A(n_560), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_538), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_527), .B(n_55), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_SL g646 ( .A1(n_593), .A2(n_140), .B(n_217), .C(n_216), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_534), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_541), .A2(n_137), .B(n_215), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_523), .A2(n_56), .B1(n_57), .B2(n_58), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_545), .A2(n_138), .B(n_214), .Y(n_650) );
NOR2xp67_ASAP7_75t_L g651 ( .A(n_564), .B(n_58), .Y(n_651) );
NOR2xp67_ASAP7_75t_L g652 ( .A(n_540), .B(n_59), .Y(n_652) );
AO31x2_ASAP7_75t_L g653 ( .A1(n_573), .A2(n_60), .A3(n_61), .B(n_62), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_610), .A2(n_61), .B(n_62), .C(n_63), .Y(n_654) );
AO31x2_ASAP7_75t_L g655 ( .A1(n_571), .A2(n_63), .A3(n_64), .B(n_65), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_SL g656 ( .A1(n_597), .A2(n_148), .B(n_209), .C(n_207), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_588), .A2(n_145), .B(n_206), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_SL g658 ( .A1(n_597), .A2(n_143), .B(n_205), .C(n_203), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_528), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_659) );
AO32x2_ASAP7_75t_L g660 ( .A1(n_561), .A2(n_66), .A3(n_67), .B1(n_68), .B2(n_69), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_595), .A2(n_149), .B(n_200), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_L g662 ( .A1(n_516), .A2(n_69), .B(n_70), .C(n_71), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_534), .Y(n_663) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_574), .A2(n_70), .B(n_72), .C(n_73), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_508), .B(n_72), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_599), .A2(n_151), .B(n_199), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_510), .B(n_73), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g668 ( .A1(n_579), .A2(n_74), .B(n_92), .C(n_94), .Y(n_668) );
AO31x2_ASAP7_75t_L g669 ( .A1(n_568), .A2(n_74), .A3(n_99), .B(n_100), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_551), .A2(n_102), .B(n_103), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_609), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_579), .A2(n_104), .B(n_107), .C(n_109), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_536), .Y(n_673) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_518), .Y(n_674) );
INVx5_ASAP7_75t_L g675 ( .A(n_552), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_513), .Y(n_676) );
AO31x2_ASAP7_75t_L g677 ( .A1(n_602), .A2(n_114), .A3(n_116), .B(n_117), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_543), .B(n_119), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_554), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_547), .Y(n_680) );
AO31x2_ASAP7_75t_L g681 ( .A1(n_596), .A2(n_120), .A3(n_122), .B(n_124), .Y(n_681) );
AOI21x1_ASAP7_75t_L g682 ( .A1(n_605), .A2(n_128), .B(n_129), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_543), .A2(n_133), .B1(n_134), .B2(n_142), .Y(n_683) );
OAI22xp33_ASAP7_75t_L g684 ( .A1(n_584), .A2(n_150), .B1(n_152), .B2(n_154), .Y(n_684) );
BUFx12f_ASAP7_75t_L g685 ( .A(n_552), .Y(n_685) );
AO21x1_ASAP7_75t_L g686 ( .A1(n_570), .A2(n_566), .B(n_611), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_613), .A2(n_159), .B(n_160), .C(n_161), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_591), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_608), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_525), .A2(n_166), .B(n_170), .C(n_172), .Y(n_690) );
BUFx10_ASAP7_75t_L g691 ( .A(n_552), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_525), .A2(n_173), .B(n_177), .C(n_178), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_515), .A2(n_180), .B(n_182), .C(n_183), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_520), .B(n_226), .Y(n_694) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_518), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_511), .B(n_184), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_526), .A2(n_185), .B1(n_186), .B2(n_188), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_549), .B(n_189), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_515), .A2(n_192), .B1(n_193), .B2(n_195), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_517), .A2(n_522), .B1(n_544), .B2(n_546), .C(n_535), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_557), .B(n_567), .Y(n_701) );
INVx8_ASAP7_75t_L g702 ( .A(n_606), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_601), .B(n_530), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_594), .A2(n_582), .B(n_580), .C(n_572), .Y(n_704) );
O2A1O1Ixp33_ASAP7_75t_L g705 ( .A1(n_509), .A2(n_512), .B(n_521), .C(n_539), .Y(n_705) );
OR2x6_ASAP7_75t_L g706 ( .A(n_569), .B(n_606), .Y(n_706) );
O2A1O1Ixp33_ASAP7_75t_SL g707 ( .A1(n_585), .A2(n_563), .B(n_612), .C(n_604), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_563), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_518), .A2(n_606), .B(n_598), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_531), .B(n_569), .Y(n_710) );
AOI31xp67_ASAP7_75t_L g711 ( .A1(n_604), .A2(n_603), .A3(n_555), .B(n_562), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_604), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_604), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_514), .B(n_463), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_533), .Y(n_715) );
O2A1O1Ixp33_ASAP7_75t_SL g716 ( .A1(n_583), .A2(n_529), .B(n_590), .C(n_586), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_577), .A2(n_574), .B(n_579), .C(n_532), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_534), .Y(n_718) );
OR2x2_ASAP7_75t_L g719 ( .A(n_524), .B(n_432), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_575), .A2(n_450), .B(n_449), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_542), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g722 ( .A1(n_577), .A2(n_574), .B(n_579), .C(n_532), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_537), .A2(n_489), .B1(n_543), .B2(n_491), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_556), .B(n_432), .Y(n_724) );
NOR2xp33_ASAP7_75t_SL g725 ( .A(n_542), .B(n_445), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_600), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_514), .Y(n_727) );
CKINVDCx11_ASAP7_75t_R g728 ( .A(n_536), .Y(n_728) );
BUFx2_ASAP7_75t_L g729 ( .A(n_533), .Y(n_729) );
A2O1A1Ixp33_ASAP7_75t_L g730 ( .A1(n_577), .A2(n_574), .B(n_579), .C(n_532), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_587), .A2(n_581), .B1(n_388), .B2(n_440), .Y(n_731) );
OR2x6_ASAP7_75t_L g732 ( .A(n_587), .B(n_445), .Y(n_732) );
INVx3_ASAP7_75t_SL g733 ( .A(n_542), .Y(n_733) );
BUFx10_ASAP7_75t_L g734 ( .A(n_534), .Y(n_734) );
INVx3_ASAP7_75t_L g735 ( .A(n_702), .Y(n_735) );
AOI22xp33_ASAP7_75t_SL g736 ( .A1(n_723), .A2(n_702), .B1(n_732), .B2(n_643), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_630), .B(n_714), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_731), .A2(n_732), .B1(n_634), .B2(n_694), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_685), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_730), .A2(n_720), .B(n_698), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_700), .A2(n_724), .B1(n_686), .B2(n_645), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_620), .B(n_623), .Y(n_742) );
AO31x2_ASAP7_75t_L g743 ( .A1(n_672), .A2(n_704), .A3(n_668), .B(n_626), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_664), .B(n_618), .C(n_662), .Y(n_744) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_729), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_619), .B(n_727), .Y(n_746) );
AOI222xp33_ASAP7_75t_L g747 ( .A1(n_667), .A2(n_671), .B1(n_710), .B2(n_651), .C1(n_638), .C2(n_637), .Y(n_747) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_674), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_640), .B(n_679), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_716), .A2(n_624), .B(n_628), .Y(n_750) );
INVx1_ASAP7_75t_SL g751 ( .A(n_715), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_675), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_676), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_629), .A2(n_639), .B(n_658), .Y(n_754) );
OAI21x1_ASAP7_75t_SL g755 ( .A1(n_682), .A2(n_709), .B(n_683), .Y(n_755) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_644), .A2(n_654), .B1(n_641), .B2(n_703), .C(n_617), .Y(n_756) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_675), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_680), .B(n_616), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_701), .B(n_719), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_726), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_635), .A2(n_665), .B1(n_694), .B2(n_678), .Y(n_761) );
BUFx3_ASAP7_75t_L g762 ( .A(n_734), .Y(n_762) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_627), .A2(n_632), .B(n_648), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_706), .B(n_689), .Y(n_764) );
OAI21xp5_ASAP7_75t_L g765 ( .A1(n_650), .A2(n_661), .B(n_696), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_675), .B(n_706), .Y(n_766) );
BUFx2_ASAP7_75t_R g767 ( .A(n_733), .Y(n_767) );
OA21x2_ASAP7_75t_L g768 ( .A1(n_690), .A2(n_692), .B(n_693), .Y(n_768) );
AO21x2_ASAP7_75t_L g769 ( .A1(n_656), .A2(n_622), .B(n_687), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_642), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_707), .A2(n_615), .B(n_705), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_642), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_649), .A2(n_659), .B1(n_652), .B2(n_725), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_642), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_666), .A2(n_614), .B(n_646), .Y(n_775) );
INVx11_ASAP7_75t_L g776 ( .A(n_734), .Y(n_776) );
INVx4_ASAP7_75t_SL g777 ( .A(n_669), .Y(n_777) );
INVx2_ASAP7_75t_SL g778 ( .A(n_691), .Y(n_778) );
AO21x2_ASAP7_75t_L g779 ( .A1(n_713), .A2(n_684), .B(n_699), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_636), .B(n_688), .Y(n_780) );
OA21x2_ASAP7_75t_L g781 ( .A1(n_633), .A2(n_670), .B(n_697), .Y(n_781) );
OA21x2_ASAP7_75t_L g782 ( .A1(n_712), .A2(n_708), .B(n_681), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_674), .A2(n_695), .B(n_631), .Y(n_783) );
AO31x2_ASAP7_75t_L g784 ( .A1(n_681), .A2(n_677), .A3(n_711), .B(n_655), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_636), .A2(n_718), .B1(n_663), .B2(n_728), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_691), .B(n_695), .Y(n_786) );
INVx3_ASAP7_75t_L g787 ( .A(n_647), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_673), .A2(n_625), .B1(n_721), .B2(n_660), .Y(n_788) );
A2O1A1Ixp33_ASAP7_75t_L g789 ( .A1(n_669), .A2(n_660), .B(n_677), .C(n_655), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_660), .Y(n_790) );
INVx4_ASAP7_75t_L g791 ( .A(n_653), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_620), .Y(n_792) );
NOR2xp67_ASAP7_75t_L g793 ( .A(n_685), .B(n_432), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_723), .A2(n_581), .B1(n_587), .B2(n_524), .Y(n_794) );
OR2x6_ASAP7_75t_L g795 ( .A(n_702), .B(n_732), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_620), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_620), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_630), .B(n_620), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_731), .A2(n_510), .B1(n_440), .B2(n_723), .C(n_432), .Y(n_799) );
OAI21x1_ASAP7_75t_SL g800 ( .A1(n_731), .A2(n_723), .B(n_657), .Y(n_800) );
A2O1A1Ixp33_ASAP7_75t_L g801 ( .A1(n_717), .A2(n_722), .B(n_730), .C(n_577), .Y(n_801) );
AOI221xp5_ASAP7_75t_L g802 ( .A1(n_723), .A2(n_438), .B1(n_532), .B2(n_510), .C(n_514), .Y(n_802) );
BUFx5_ASAP7_75t_L g803 ( .A(n_685), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_630), .B(n_620), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_630), .B(n_620), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_620), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_620), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_630), .B(n_620), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_630), .B(n_620), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_620), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_723), .B(n_432), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_621), .A2(n_575), .B(n_717), .Y(n_812) );
INVx2_ASAP7_75t_SL g813 ( .A(n_702), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_728), .Y(n_814) );
AND2x4_ASAP7_75t_L g815 ( .A(n_706), .B(n_540), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_621), .A2(n_575), .B(n_717), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_723), .B(n_441), .Y(n_817) );
INVx2_ASAP7_75t_SL g818 ( .A(n_702), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_620), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_630), .B(n_723), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_620), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_630), .B(n_620), .Y(n_822) );
NOR2x1_ASAP7_75t_R g823 ( .A(n_728), .B(n_445), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_723), .B(n_432), .Y(n_824) );
INVxp67_ASAP7_75t_L g825 ( .A(n_729), .Y(n_825) );
OR2x6_ASAP7_75t_L g826 ( .A(n_702), .B(n_732), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_723), .B(n_432), .Y(n_827) );
BUFx3_ASAP7_75t_L g828 ( .A(n_685), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_723), .B(n_432), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_620), .Y(n_830) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_729), .Y(n_831) );
INVx4_ASAP7_75t_R g832 ( .A(n_647), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_620), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_719), .B(n_432), .Y(n_834) );
AOI221xp5_ASAP7_75t_L g835 ( .A1(n_723), .A2(n_438), .B1(n_532), .B2(n_510), .C(n_514), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_630), .B(n_620), .Y(n_836) );
AOI21xp5_ASAP7_75t_SL g837 ( .A1(n_738), .A2(n_801), .B(n_789), .Y(n_837) );
BUFx2_ASAP7_75t_L g838 ( .A(n_748), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_770), .Y(n_839) );
INVx2_ASAP7_75t_SL g840 ( .A(n_803), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_817), .A2(n_794), .B1(n_799), .B2(n_800), .Y(n_841) );
AND2x4_ASAP7_75t_L g842 ( .A(n_795), .B(n_826), .Y(n_842) );
NAND2x1_ASAP7_75t_L g843 ( .A(n_755), .B(n_791), .Y(n_843) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_751), .Y(n_844) );
BUFx2_ASAP7_75t_L g845 ( .A(n_795), .Y(n_845) );
OA21x2_ASAP7_75t_L g846 ( .A1(n_812), .A2(n_816), .B(n_772), .Y(n_846) );
AO21x2_ASAP7_75t_L g847 ( .A1(n_774), .A2(n_740), .B(n_754), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_790), .Y(n_848) );
AOI221xp5_ASAP7_75t_L g849 ( .A1(n_802), .A2(n_835), .B1(n_741), .B2(n_756), .C(n_749), .Y(n_849) );
AND2x4_ASAP7_75t_L g850 ( .A(n_795), .B(n_826), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_746), .Y(n_851) );
INVx3_ASAP7_75t_SL g852 ( .A(n_803), .Y(n_852) );
OA21x2_ASAP7_75t_L g853 ( .A1(n_750), .A2(n_771), .B(n_763), .Y(n_853) );
OA21x2_ASAP7_75t_L g854 ( .A1(n_763), .A2(n_775), .B(n_765), .Y(n_854) );
INVx4_ASAP7_75t_L g855 ( .A(n_826), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_758), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_811), .B(n_824), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_827), .B(n_829), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_742), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_820), .B(n_836), .Y(n_860) );
INVxp67_ASAP7_75t_SL g861 ( .A(n_738), .Y(n_861) );
OR2x6_ASAP7_75t_L g862 ( .A(n_815), .B(n_766), .Y(n_862) );
BUFx3_ASAP7_75t_L g863 ( .A(n_828), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_792), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_796), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_797), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_806), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_807), .Y(n_868) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_751), .Y(n_869) );
OR2x6_ASAP7_75t_L g870 ( .A(n_815), .B(n_752), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_810), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_761), .A2(n_736), .B1(n_737), .B2(n_773), .Y(n_872) );
AND2x4_ASAP7_75t_L g873 ( .A(n_819), .B(n_821), .Y(n_873) );
AO21x2_ASAP7_75t_L g874 ( .A1(n_744), .A2(n_788), .B(n_769), .Y(n_874) );
NAND2x1p5_ASAP7_75t_L g875 ( .A(n_753), .B(n_760), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_836), .B(n_808), .Y(n_876) );
OR2x2_ASAP7_75t_L g877 ( .A(n_798), .B(n_809), .Y(n_877) );
AOI222xp33_ASAP7_75t_SL g878 ( .A1(n_825), .A2(n_745), .B1(n_831), .B2(n_739), .C1(n_830), .C2(n_833), .Y(n_878) );
AO21x2_ASAP7_75t_L g879 ( .A1(n_779), .A2(n_805), .B(n_808), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_804), .B(n_822), .Y(n_880) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_793), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_804), .Y(n_882) );
OR2x2_ASAP7_75t_L g883 ( .A(n_805), .B(n_809), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_784), .Y(n_884) );
AO21x2_ASAP7_75t_L g885 ( .A1(n_779), .A2(n_783), .B(n_773), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_784), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_759), .B(n_747), .Y(n_887) );
OA21x2_ASAP7_75t_L g888 ( .A1(n_777), .A2(n_782), .B(n_786), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_834), .A2(n_757), .B1(n_787), .B2(n_785), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_803), .Y(n_890) );
OAI321xp33_ASAP7_75t_L g891 ( .A1(n_780), .A2(n_764), .A3(n_778), .B1(n_813), .B2(n_818), .C(n_747), .Y(n_891) );
BUFx3_ASAP7_75t_L g892 ( .A(n_803), .Y(n_892) );
OAI221xp5_ASAP7_75t_L g893 ( .A1(n_787), .A2(n_735), .B1(n_762), .B2(n_768), .C(n_781), .Y(n_893) );
AOI22xp33_ASAP7_75t_SL g894 ( .A1(n_803), .A2(n_735), .B1(n_832), .B2(n_781), .Y(n_894) );
OA21x2_ASAP7_75t_L g895 ( .A1(n_743), .A2(n_823), .B(n_814), .Y(n_895) );
BUFx3_ASAP7_75t_L g896 ( .A(n_776), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_743), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_767), .B(n_817), .Y(n_898) );
AND2x4_ASAP7_75t_L g899 ( .A(n_795), .B(n_826), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_746), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_746), .Y(n_901) );
INVxp67_ASAP7_75t_L g902 ( .A(n_834), .Y(n_902) );
AOI31xp33_ASAP7_75t_L g903 ( .A1(n_823), .A2(n_736), .A3(n_794), .B(n_723), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_811), .B(n_829), .Y(n_904) );
INVxp67_ASAP7_75t_SL g905 ( .A(n_758), .Y(n_905) );
AOI21xp5_ASAP7_75t_SL g906 ( .A1(n_738), .A2(n_732), .B(n_694), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_811), .B(n_829), .Y(n_907) );
HB1xp67_ASAP7_75t_L g908 ( .A(n_751), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_770), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_770), .Y(n_910) );
AOI221xp5_ASAP7_75t_L g911 ( .A1(n_799), .A2(n_438), .B1(n_802), .B2(n_835), .C(n_817), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_839), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_911), .A2(n_887), .B1(n_849), .B2(n_872), .Y(n_913) );
INVx3_ASAP7_75t_L g914 ( .A(n_843), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_897), .B(n_848), .Y(n_915) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_905), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_909), .B(n_910), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_909), .B(n_910), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_884), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_903), .B(n_898), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_879), .B(n_886), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_879), .B(n_886), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_880), .B(n_882), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_880), .B(n_882), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_879), .B(n_861), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_857), .B(n_904), .Y(n_926) );
INVxp67_ASAP7_75t_SL g927 ( .A(n_875), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_860), .B(n_859), .Y(n_928) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_844), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_857), .B(n_904), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_841), .A2(n_887), .B1(n_907), .B2(n_858), .Y(n_931) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_869), .Y(n_932) );
OR2x2_ASAP7_75t_L g933 ( .A(n_907), .B(n_877), .Y(n_933) );
INVx4_ASAP7_75t_SL g934 ( .A(n_852), .Y(n_934) );
INVx4_ASAP7_75t_L g935 ( .A(n_852), .Y(n_935) );
BUFx2_ASAP7_75t_L g936 ( .A(n_838), .Y(n_936) );
OR2x2_ASAP7_75t_L g937 ( .A(n_877), .B(n_883), .Y(n_937) );
OR2x2_ASAP7_75t_L g938 ( .A(n_883), .B(n_876), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_837), .B(n_846), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_856), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_837), .B(n_846), .Y(n_941) );
HB1xp67_ASAP7_75t_L g942 ( .A(n_908), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_870), .Y(n_943) );
AOI221xp5_ASAP7_75t_L g944 ( .A1(n_891), .A2(n_906), .B1(n_902), .B2(n_901), .C(n_900), .Y(n_944) );
OR2x2_ASAP7_75t_L g945 ( .A(n_906), .B(n_851), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_854), .B(n_847), .Y(n_946) );
INVx2_ASAP7_75t_SL g947 ( .A(n_935), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_926), .B(n_873), .Y(n_948) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_944), .B(n_878), .C(n_893), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_926), .B(n_885), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_926), .B(n_873), .Y(n_951) );
INVxp67_ASAP7_75t_L g952 ( .A(n_929), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_919), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_930), .B(n_885), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_930), .B(n_885), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_930), .B(n_854), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_917), .B(n_854), .Y(n_957) );
OR2x2_ASAP7_75t_L g958 ( .A(n_933), .B(n_916), .Y(n_958) );
OR2x2_ASAP7_75t_L g959 ( .A(n_933), .B(n_874), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_938), .B(n_873), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_912), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_912), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_917), .B(n_888), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_938), .B(n_864), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_918), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_923), .B(n_866), .Y(n_966) );
AND2x4_ASAP7_75t_L g967 ( .A(n_914), .B(n_847), .Y(n_967) );
INVx3_ASAP7_75t_L g968 ( .A(n_914), .Y(n_968) );
OR2x2_ASAP7_75t_L g969 ( .A(n_937), .B(n_895), .Y(n_969) );
NAND2xp5_ASAP7_75t_SL g970 ( .A(n_935), .B(n_899), .Y(n_970) );
INVx2_ASAP7_75t_SL g971 ( .A(n_935), .Y(n_971) );
OR2x2_ASAP7_75t_L g972 ( .A(n_937), .B(n_895), .Y(n_972) );
INVx2_ASAP7_75t_SL g973 ( .A(n_935), .Y(n_973) );
AND2x4_ASAP7_75t_SL g974 ( .A(n_943), .B(n_899), .Y(n_974) );
AND3x1_ASAP7_75t_L g975 ( .A(n_920), .B(n_881), .C(n_840), .Y(n_975) );
NOR2xp33_ASAP7_75t_L g976 ( .A(n_913), .B(n_863), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_915), .B(n_867), .Y(n_977) );
NOR2xp33_ASAP7_75t_L g978 ( .A(n_913), .B(n_863), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_915), .B(n_871), .Y(n_979) );
AND2x4_ASAP7_75t_L g980 ( .A(n_914), .B(n_899), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_921), .B(n_865), .Y(n_981) );
BUFx3_ASAP7_75t_L g982 ( .A(n_936), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_921), .B(n_868), .Y(n_983) );
INVx1_ASAP7_75t_SL g984 ( .A(n_934), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_921), .B(n_853), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_922), .B(n_853), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_961), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_961), .Y(n_988) );
INVx2_ASAP7_75t_SL g989 ( .A(n_947), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_956), .B(n_946), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g991 ( .A(n_976), .B(n_855), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_965), .B(n_925), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_956), .B(n_925), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_985), .B(n_946), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_950), .B(n_925), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_953), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_965), .B(n_922), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_962), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_985), .B(n_946), .Y(n_999) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_958), .B(n_929), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_981), .B(n_922), .Y(n_1001) );
OR2x2_ASAP7_75t_L g1002 ( .A(n_958), .B(n_932), .Y(n_1002) );
INVx2_ASAP7_75t_SL g1003 ( .A(n_947), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_981), .B(n_932), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_950), .B(n_939), .Y(n_1005) );
OR2x2_ASAP7_75t_L g1006 ( .A(n_959), .B(n_942), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_983), .B(n_942), .Y(n_1007) );
OR2x2_ASAP7_75t_L g1008 ( .A(n_959), .B(n_923), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_983), .B(n_940), .Y(n_1009) );
INVx1_ASAP7_75t_SL g1010 ( .A(n_982), .Y(n_1010) );
INVxp33_ASAP7_75t_L g1011 ( .A(n_978), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_954), .B(n_940), .Y(n_1012) );
INVx3_ASAP7_75t_SL g1013 ( .A(n_971), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_954), .B(n_939), .Y(n_1014) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_967), .B(n_939), .Y(n_1015) );
NOR2x1_ASAP7_75t_L g1016 ( .A(n_970), .B(n_895), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_955), .B(n_941), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_955), .B(n_941), .Y(n_1018) );
INVxp67_ASAP7_75t_SL g1019 ( .A(n_952), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_986), .B(n_941), .Y(n_1020) );
NAND2xp5_ASAP7_75t_SL g1021 ( .A(n_1013), .B(n_975), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1000), .Y(n_1022) );
NOR2xp33_ASAP7_75t_L g1023 ( .A(n_1011), .B(n_948), .Y(n_1023) );
NOR2x1_ASAP7_75t_L g1024 ( .A(n_1016), .B(n_984), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_990), .B(n_986), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_1004), .B(n_977), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_1004), .B(n_977), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_987), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_990), .B(n_957), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_991), .A2(n_949), .B1(n_945), .B2(n_944), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_987), .Y(n_1031) );
INVx1_ASAP7_75t_SL g1032 ( .A(n_1013), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1000), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1002), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_1013), .A2(n_973), .B1(n_971), .B2(n_945), .Y(n_1035) );
AND2x4_ASAP7_75t_L g1036 ( .A(n_1015), .B(n_967), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_988), .Y(n_1037) );
INVxp67_ASAP7_75t_L g1038 ( .A(n_1019), .Y(n_1038) );
INVxp67_ASAP7_75t_L g1039 ( .A(n_1019), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_988), .Y(n_1040) );
NOR2xp33_ASAP7_75t_L g1041 ( .A(n_1002), .B(n_951), .Y(n_1041) );
INVx2_ASAP7_75t_L g1042 ( .A(n_996), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_998), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_990), .B(n_957), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1007), .B(n_979), .Y(n_1045) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_989), .Y(n_1046) );
BUFx2_ASAP7_75t_L g1047 ( .A(n_989), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_1006), .B(n_969), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_994), .B(n_963), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1007), .Y(n_1050) );
AND2x2_ASAP7_75t_SL g1051 ( .A(n_1015), .B(n_974), .Y(n_1051) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_1023), .A2(n_1020), .B1(n_1014), .B2(n_1005), .C(n_1018), .Y(n_1052) );
AOI211x1_ASAP7_75t_L g1053 ( .A1(n_1021), .A2(n_1009), .B(n_1020), .C(n_964), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_1050), .B(n_995), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1022), .B(n_995), .Y(n_1055) );
NAND2x1_ASAP7_75t_L g1056 ( .A(n_1047), .B(n_989), .Y(n_1056) );
AOI21xp33_ASAP7_75t_SL g1057 ( .A1(n_1051), .A2(n_1003), .B(n_973), .Y(n_1057) );
NAND2xp5_ASAP7_75t_SL g1058 ( .A(n_1032), .B(n_1003), .Y(n_1058) );
AOI22xp5_ASAP7_75t_L g1059 ( .A1(n_1030), .A2(n_1020), .B1(n_1017), .B2(n_1014), .Y(n_1059) );
INVx2_ASAP7_75t_L g1060 ( .A(n_1042), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1028), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1025), .B(n_993), .Y(n_1062) );
NOR2xp33_ASAP7_75t_L g1063 ( .A(n_1038), .B(n_1010), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1028), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1031), .Y(n_1065) );
AND2x4_ASAP7_75t_L g1066 ( .A(n_1036), .B(n_1015), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1031), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1025), .B(n_993), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g1069 ( .A1(n_1039), .A2(n_1018), .B1(n_1017), .B2(n_1005), .C(n_999), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1033), .B(n_994), .Y(n_1070) );
INVx2_ASAP7_75t_L g1071 ( .A(n_1042), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1037), .Y(n_1072) );
AOI22xp5_ASAP7_75t_L g1073 ( .A1(n_1059), .A2(n_1034), .B1(n_1036), .B2(n_1051), .Y(n_1073) );
AOI21xp5_ASAP7_75t_L g1074 ( .A1(n_1056), .A2(n_1047), .B(n_1035), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1060), .Y(n_1075) );
OAI221xp5_ASAP7_75t_L g1076 ( .A1(n_1069), .A2(n_1046), .B1(n_1048), .B2(n_1024), .C(n_1016), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1061), .Y(n_1077) );
A2O1A1Ixp33_ASAP7_75t_L g1078 ( .A1(n_1057), .A2(n_1046), .B(n_1036), .C(n_1041), .Y(n_1078) );
AOI222xp33_ASAP7_75t_L g1079 ( .A1(n_1052), .A2(n_931), .B1(n_999), .B2(n_994), .C1(n_1049), .C2(n_1044), .Y(n_1079) );
AOI221xp5_ASAP7_75t_L g1080 ( .A1(n_1053), .A2(n_1026), .B1(n_1027), .B2(n_1045), .C(n_1049), .Y(n_1080) );
AOI322xp5_ASAP7_75t_L g1081 ( .A1(n_1062), .A2(n_1044), .A3(n_1029), .B1(n_999), .B2(n_1001), .C1(n_960), .C2(n_992), .Y(n_1081) );
AOI21xp33_ASAP7_75t_L g1082 ( .A1(n_1063), .A2(n_889), .B(n_890), .Y(n_1082) );
AOI322xp5_ASAP7_75t_L g1083 ( .A1(n_1068), .A2(n_1029), .A3(n_1001), .B1(n_992), .B2(n_842), .C1(n_850), .C2(n_997), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1064), .Y(n_1084) );
NOR3xp33_ASAP7_75t_L g1085 ( .A(n_1058), .B(n_894), .C(n_855), .Y(n_1085) );
AOI22xp5_ASAP7_75t_L g1086 ( .A1(n_1063), .A2(n_1015), .B1(n_1048), .B2(n_1012), .Y(n_1086) );
AOI22xp5_ASAP7_75t_L g1087 ( .A1(n_1079), .A2(n_1058), .B1(n_1066), .B2(n_1054), .Y(n_1087) );
AOI221xp5_ASAP7_75t_L g1088 ( .A1(n_1076), .A2(n_1072), .B1(n_1065), .B2(n_1067), .C(n_1070), .Y(n_1088) );
NAND4xp25_ASAP7_75t_L g1089 ( .A(n_1085), .B(n_842), .C(n_850), .D(n_855), .Y(n_1089) );
NOR2xp33_ASAP7_75t_R g1090 ( .A(n_1077), .B(n_896), .Y(n_1090) );
OAI21xp5_ASAP7_75t_L g1091 ( .A1(n_1074), .A2(n_1066), .B(n_1003), .Y(n_1091) );
O2A1O1Ixp33_ASAP7_75t_L g1092 ( .A1(n_1078), .A2(n_845), .B(n_842), .C(n_850), .Y(n_1092) );
AND2x2_ASAP7_75t_SL g1093 ( .A(n_1073), .B(n_1066), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1084), .Y(n_1094) );
OAI22xp33_ASAP7_75t_L g1095 ( .A1(n_1086), .A2(n_1010), .B1(n_1055), .B2(n_969), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1094), .Y(n_1096) );
OAI211xp5_ASAP7_75t_L g1097 ( .A1(n_1089), .A2(n_1083), .B(n_1081), .C(n_1082), .Y(n_1097) );
NAND3xp33_ASAP7_75t_SL g1098 ( .A(n_1092), .B(n_1080), .C(n_845), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1087), .B(n_1075), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_1088), .A2(n_1082), .B1(n_1071), .B2(n_1060), .C(n_966), .Y(n_1100) );
NAND4xp25_ASAP7_75t_L g1101 ( .A(n_1091), .B(n_896), .C(n_972), .D(n_980), .Y(n_1101) );
NOR2x1p5_ASAP7_75t_L g1102 ( .A(n_1099), .B(n_1090), .Y(n_1102) );
NAND4xp75_ASAP7_75t_L g1103 ( .A(n_1100), .B(n_1093), .C(n_840), .D(n_1095), .Y(n_1103) );
AND2x4_ASAP7_75t_L g1104 ( .A(n_1096), .B(n_1071), .Y(n_1104) );
NOR3xp33_ASAP7_75t_SL g1105 ( .A(n_1098), .B(n_928), .C(n_1012), .Y(n_1105) );
NAND5xp2_ASAP7_75t_L g1106 ( .A(n_1097), .B(n_875), .C(n_927), .D(n_928), .E(n_934), .Y(n_1106) );
AND3x1_ASAP7_75t_L g1107 ( .A(n_1106), .B(n_1101), .C(n_968), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_1102), .B(n_1037), .Y(n_1108) );
OR3x1_ASAP7_75t_L g1109 ( .A(n_1105), .B(n_1043), .C(n_1040), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1104), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1110), .B(n_1104), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1108), .Y(n_1112) );
OA22x2_ASAP7_75t_L g1113 ( .A1(n_1108), .A2(n_1103), .B1(n_974), .B2(n_870), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1111), .Y(n_1114) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_1112), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_1113), .A2(n_1109), .B1(n_1107), .B2(n_1006), .Y(n_1116) );
XNOR2xp5_ASAP7_75t_L g1117 ( .A(n_1114), .B(n_1107), .Y(n_1117) );
AOI222xp33_ASAP7_75t_L g1118 ( .A1(n_1115), .A2(n_892), .B1(n_1040), .B2(n_1043), .C1(n_934), .C2(n_980), .Y(n_1118) );
OAI21xp5_ASAP7_75t_L g1119 ( .A1(n_1117), .A2(n_1116), .B(n_892), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_1118), .B(n_1008), .Y(n_1120) );
AO221x2_ASAP7_75t_L g1121 ( .A1(n_1119), .A2(n_1120), .B1(n_924), .B2(n_1009), .C(n_997), .Y(n_1121) );
AOI22xp5_ASAP7_75t_L g1122 ( .A1(n_1121), .A2(n_862), .B1(n_934), .B2(n_979), .Y(n_1122) );
endmodule