module fake_jpeg_29213_n_223 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_223);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_40),
.B(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_10),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_48),
.Y(n_66)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_1),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_16),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_20),
.B(n_15),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_18),
.B1(n_32),
.B2(n_29),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_80),
.B1(n_83),
.B2(n_1),
.Y(n_114)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_39),
.A2(n_17),
.B1(n_22),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_85),
.B1(n_48),
.B2(n_40),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_19),
.B1(n_32),
.B2(n_28),
.Y(n_80)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_24),
.B1(n_28),
.B2(n_19),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_17),
.B1(n_22),
.B2(n_36),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_26),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_27),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_27),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_22),
.Y(n_105)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_94),
.B(n_107),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_110),
.B(n_102),
.Y(n_125)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_46),
.B1(n_42),
.B2(n_51),
.Y(n_99)
);

AO22x1_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_101),
.B1(n_89),
.B2(n_70),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_84),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_56),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_64),
.B(n_35),
.Y(n_106)
);

OR2x6_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_73),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_26),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_22),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_14),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_23),
.B1(n_2),
.B2(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_114),
.B1(n_73),
.B2(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_61),
.B(n_23),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_61),
.B(n_11),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_11),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_120),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_84),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_95),
.B1(n_100),
.B2(n_99),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_125),
.B1(n_132),
.B2(n_134),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_67),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_117),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_131),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_135),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_81),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_99),
.A2(n_82),
.B1(n_68),
.B2(n_91),
.Y(n_134)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

AOI32xp33_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_70),
.A3(n_78),
.B1(n_13),
.B2(n_12),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_111),
.Y(n_152)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

OA22x2_ASAP7_75t_SL g143 ( 
.A1(n_99),
.A2(n_91),
.B1(n_92),
.B2(n_71),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_143),
.A2(n_104),
.B(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_154),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_101),
.B(n_107),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

NOR4xp25_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_94),
.C(n_120),
.D(n_111),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_148),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_125),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_160),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_130),
.C(n_121),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_112),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_159),
.B(n_138),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_96),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_129),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_166),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_146),
.B(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_167),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_130),
.B1(n_135),
.B2(n_143),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_151),
.B1(n_161),
.B2(n_154),
.C(n_144),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_149),
.B(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_191),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_153),
.C(n_158),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_167),
.C(n_174),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_151),
.B1(n_149),
.B2(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

OAI322xp33_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_171),
.A3(n_191),
.B1(n_180),
.B2(n_177),
.C1(n_186),
.C2(n_181),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_171),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_161),
.B(n_162),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_195),
.C(n_197),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_194),
.B(n_200),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_170),
.C(n_175),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_184),
.B(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_196),
.B(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_168),
.C(n_166),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_164),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_181),
.B1(n_186),
.B2(n_190),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_98),
.B1(n_71),
.B2(n_78),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

AOI31xp67_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_157),
.A3(n_112),
.B(n_145),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_207),
.Y(n_210)
);

AOI31xp67_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_96),
.A3(n_136),
.B(n_141),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_SL g208 ( 
.A(n_202),
.B(n_103),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_211),
.B(n_212),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_98),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_209),
.A2(n_201),
.B(n_202),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_215),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_87),
.B1(n_6),
.B2(n_7),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

AOI21x1_ASAP7_75t_SL g215 ( 
.A1(n_208),
.A2(n_2),
.B(n_7),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_87),
.C(n_2),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_8),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_218),
.Y(n_223)
);


endmodule