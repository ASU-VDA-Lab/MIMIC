module real_jpeg_1377_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_1),
.B(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_1),
.B(n_28),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_1),
.B(n_51),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_1),
.B(n_26),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_2),
.B(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_4),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_4),
.B(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_4),
.B(n_36),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_51),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_28),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_4),
.B(n_26),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_5),
.B(n_32),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_61),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_5),
.B(n_53),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_8),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_8),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_8),
.B(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_8),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_8),
.B(n_53),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_8),
.B(n_51),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_9),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_9),
.B(n_53),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_9),
.B(n_26),
.Y(n_122)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_11),
.B(n_28),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_14),
.B(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_14),
.B(n_61),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_14),
.B(n_28),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_92),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_20),
.B(n_92),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_56),
.C(n_81),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_21),
.B(n_204),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_21),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_38),
.CI(n_42),
.CON(n_21),
.SN(n_21)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_22),
.B(n_38),
.C(n_42),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_31),
.C(n_35),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_23),
.A2(n_24),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_25),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_25),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_161)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_27),
.A2(n_71),
.B1(n_74),
.B2(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_29),
.B(n_127),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_31),
.B(n_35),
.Y(n_200)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_41),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_41),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_43),
.B(n_50),
.C(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_44),
.B(n_72),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_44),
.B(n_103),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_45),
.B(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_56),
.B(n_81),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_68),
.B2(n_80),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_69),
.C(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_65),
.C(n_67),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.C(n_79),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.C(n_90),
.Y(n_81)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_82),
.B(n_86),
.CI(n_90),
.CON(n_194),
.SN(n_194)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.C(n_89),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_89),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_140),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g209 ( 
.A(n_92),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_114),
.CI(n_115),
.CON(n_92),
.SN(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_104),
.B2(n_105),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_112),
.B2(n_113),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_110),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_122),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_125),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_202),
.B(n_206),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_190),
.B(n_201),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_162),
.B(n_189),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_153),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_153),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_143),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.C(n_138),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_137),
.CI(n_138),
.CON(n_154),
.SN(n_154)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_141),
.C(n_143),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_149),
.C(n_150),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.C(n_161),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_186),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_154),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_156),
.B1(n_161),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_183),
.B(n_188),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_174),
.B(n_182),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_170),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_168),
.C(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_177),
.B(n_181),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_185),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_191),
.B(n_192),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_197),
.C(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_205),
.Y(n_206)
);


endmodule