module fake_netlist_5_2073_n_1741 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_1741);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1741;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_144;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_146;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_149;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_147;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_145;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_27),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_141),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

BUFx8_ASAP7_75t_SL g147 ( 
.A(n_4),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_105),
.Y(n_148)
);

BUFx10_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_96),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_11),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_10),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_111),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_16),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_51),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_4),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_60),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_63),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_53),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_87),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_85),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_7),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_79),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_48),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_45),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_20),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_115),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_7),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_1),
.Y(n_175)
);

BUFx2_ASAP7_75t_SL g176 ( 
.A(n_19),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_32),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_56),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_68),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_77),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_74),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_41),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_54),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_82),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_71),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_37),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_1),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_94),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_124),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_45),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_20),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_131),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_84),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_83),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_81),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_48),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_17),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_12),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_25),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_129),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_93),
.Y(n_204)
);

BUFx2_ASAP7_75t_SL g205 ( 
.A(n_134),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_28),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_25),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_100),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_58),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_65),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_139),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_47),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_136),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_75),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_118),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_143),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_21),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_15),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_142),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_128),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_12),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_8),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_70),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_14),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_50),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_18),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_69),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_14),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_10),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_62),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_109),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_49),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_138),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_106),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_91),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_3),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_36),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_11),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_112),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_59),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_28),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_55),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_110),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_27),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_90),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_18),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_97),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_46),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_78),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_61),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_21),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_13),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_113),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_107),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_16),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_114),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_43),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_9),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_108),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_117),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_86),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_43),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_22),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_22),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_103),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_140),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_17),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_123),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_13),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_36),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_26),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_33),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_47),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_132),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_0),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_42),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_80),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_26),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_49),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_38),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_38),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_66),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_122),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_72),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_37),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_30),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_41),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_9),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_46),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_6),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_192),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_183),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_192),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_252),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_164),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_152),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_147),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_168),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_145),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_152),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_203),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_167),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_167),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_169),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_146),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_169),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_148),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_188),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_188),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_224),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_224),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_226),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_237),
.Y(n_320)
);

BUFx2_ASAP7_75t_SL g321 ( 
.A(n_284),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_238),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_150),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_238),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_267),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_151),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_153),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_176),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_155),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_157),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_144),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_183),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_153),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_165),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_209),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_165),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_173),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_173),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_289),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_210),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_182),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_182),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_269),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_158),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_286),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_286),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_277),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_181),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_181),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_186),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_215),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_215),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_186),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_189),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_234),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_189),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_299),
.Y(n_363)
);

NOR2x1_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_282),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_301),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_282),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_357),
.A2(n_187),
.B1(n_288),
.B2(n_200),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_301),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_240),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_292),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_352),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_317),
.A2(n_229),
.B1(n_228),
.B2(n_257),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_305),
.Y(n_377)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_355),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_240),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_295),
.Y(n_381)
);

AND3x1_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_278),
.C(n_198),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_329),
.B(n_284),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_307),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

AND2x6_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_163),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_307),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_361),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_303),
.A2(n_236),
.B1(n_217),
.B2(n_290),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_304),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_359),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_321),
.B(n_161),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_306),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_335),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_343),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_291),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_321),
.B(n_166),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_336),
.B(n_235),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_291),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_310),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_309),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_309),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_311),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_353),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_338),
.B(n_339),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_294),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_311),
.Y(n_413)
);

OA21x2_ASAP7_75t_L g414 ( 
.A1(n_340),
.A2(n_201),
.B(n_190),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_294),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_296),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_296),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_313),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_313),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_172),
.Y(n_420)
);

BUFx12f_ASAP7_75t_L g421 ( 
.A(n_302),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_314),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_360),
.A2(n_202),
.B1(n_285),
.B2(n_281),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_293),
.A2(n_199),
.B1(n_280),
.B2(n_279),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_345),
.B(n_235),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_374),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_374),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_380),
.B(n_312),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_380),
.B(n_334),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_324),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_362),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_374),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_367),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_367),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_328),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_367),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_374),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

OAI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_420),
.A2(n_356),
.B1(n_190),
.B2(n_201),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_383),
.B(n_331),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_376),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_397),
.B(n_332),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_383),
.B(n_348),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_394),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_366),
.B(n_160),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_376),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_406),
.B(n_346),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_376),
.Y(n_459)
);

INVx6_ASAP7_75t_L g460 ( 
.A(n_378),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

NOR3xp33_ASAP7_75t_L g462 ( 
.A(n_368),
.B(n_278),
.C(n_198),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_410),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_403),
.B(n_149),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

INVx5_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_379),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_384),
.B(n_345),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_366),
.B(n_219),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_379),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_410),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_371),
.Y(n_472)
);

INVx6_ASAP7_75t_L g473 ( 
.A(n_378),
.Y(n_473)
);

BUFx10_ASAP7_75t_L g474 ( 
.A(n_424),
.Y(n_474)
);

AOI21x1_ASAP7_75t_L g475 ( 
.A1(n_414),
.A2(n_420),
.B(n_404),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_379),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_366),
.B(n_204),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_403),
.B(n_347),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_387),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_L g483 ( 
.A(n_424),
.B(n_163),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_370),
.B(n_347),
.Y(n_484)
);

BUFx4f_ASAP7_75t_L g485 ( 
.A(n_414),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_387),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_387),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_384),
.B(n_349),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_387),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_388),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_388),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_366),
.B(n_378),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_425),
.B(n_149),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_370),
.A2(n_265),
.B1(n_266),
.B2(n_242),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_388),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_388),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_378),
.B(n_231),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_425),
.B(n_149),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_411),
.Y(n_501)
);

OR2x6_ASAP7_75t_L g502 ( 
.A(n_421),
.B(n_205),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_395),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_381),
.B(n_349),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_395),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_395),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_395),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_363),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_381),
.B(n_350),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_395),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_378),
.Y(n_514)
);

INVx8_ASAP7_75t_L g515 ( 
.A(n_389),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_399),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_411),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_399),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_399),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_399),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_371),
.B(n_350),
.Y(n_521)
);

BUFx8_ASAP7_75t_SL g522 ( 
.A(n_398),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_412),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_378),
.B(n_233),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_412),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_415),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_423),
.B(n_382),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_404),
.A2(n_176),
.B1(n_205),
.B2(n_254),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_399),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_415),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_399),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_R g534 ( 
.A(n_414),
.B(n_154),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_423),
.B(n_149),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_415),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_378),
.B(n_253),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_417),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_417),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_414),
.Y(n_541)
);

NAND3xp33_ASAP7_75t_L g542 ( 
.A(n_382),
.B(n_159),
.C(n_156),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_414),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_372),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_384),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_417),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_384),
.B(n_297),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_372),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_417),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_368),
.B(n_162),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_372),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_364),
.Y(n_552)
);

INVx4_ASAP7_75t_SL g553 ( 
.A(n_389),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_364),
.B(n_171),
.C(n_170),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_385),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_385),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_385),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_391),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_404),
.B(n_391),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_404),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_391),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_392),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_392),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_392),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_426),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_426),
.B(n_268),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_401),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_402),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_375),
.B(n_314),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_365),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_426),
.B(n_163),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_402),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_365),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_369),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_439),
.B(n_426),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_453),
.B(n_219),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_474),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_545),
.B(n_209),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_479),
.B(n_223),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_485),
.B(n_163),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_431),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_565),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_565),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_429),
.A2(n_254),
.B1(n_230),
.B2(n_283),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_574),
.B(n_230),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_L g586 ( 
.A(n_462),
.B(n_375),
.C(n_175),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_574),
.B(n_274),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_431),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_560),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_431),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_432),
.B(n_393),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_574),
.B(n_274),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_485),
.B(n_163),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_430),
.B(n_401),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_430),
.B(n_393),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_557),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_552),
.B(n_283),
.Y(n_597)
);

INVx8_ASAP7_75t_L g598 ( 
.A(n_502),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_570),
.B(n_369),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_534),
.A2(n_245),
.B1(n_195),
.B2(n_194),
.Y(n_600)
);

NOR2x1p5_ASAP7_75t_L g601 ( 
.A(n_569),
.B(n_421),
.Y(n_601)
);

AOI22x1_ASAP7_75t_L g602 ( 
.A1(n_543),
.A2(n_422),
.B1(n_419),
.B2(n_418),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_480),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_570),
.B(n_373),
.Y(n_604)
);

INVxp33_ASAP7_75t_L g605 ( 
.A(n_472),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_573),
.B(n_373),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_573),
.B(n_377),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_557),
.Y(n_608)
);

INVx8_ASAP7_75t_L g609 ( 
.A(n_502),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_502),
.B(n_421),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_469),
.B(n_377),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_472),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_560),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_433),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_469),
.B(n_386),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_485),
.B(n_209),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_469),
.B(n_386),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_485),
.B(n_209),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_474),
.B(n_390),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_512),
.B(n_390),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_541),
.B(n_209),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_512),
.B(n_526),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_541),
.A2(n_422),
.B1(n_419),
.B2(n_418),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_512),
.B(n_396),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_512),
.B(n_396),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_557),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_541),
.B(n_209),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_563),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_455),
.B(n_400),
.Y(n_629)
);

BUFx6f_ASAP7_75t_SL g630 ( 
.A(n_502),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_526),
.B(n_400),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_526),
.B(n_538),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_526),
.B(n_407),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_538),
.B(n_407),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_468),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_SL g636 ( 
.A(n_550),
.B(n_535),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_501),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_560),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_538),
.B(n_408),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_538),
.B(n_209),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_521),
.B(n_174),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_456),
.B(n_209),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_563),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_484),
.B(n_408),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g645 ( 
.A(n_480),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_501),
.B(n_409),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_524),
.B(n_178),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_504),
.B(n_409),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_493),
.A2(n_533),
.B(n_520),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_433),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_440),
.Y(n_651)
);

BUFx5_ASAP7_75t_L g652 ( 
.A(n_427),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_478),
.B(n_179),
.Y(n_653)
);

AND2x4_ASAP7_75t_SL g654 ( 
.A(n_502),
.B(n_162),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_559),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_501),
.B(n_413),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_513),
.B(n_413),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_569),
.B(n_177),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_571),
.B(n_180),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_513),
.B(n_402),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_524),
.B(n_184),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_513),
.B(n_405),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_509),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_440),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_517),
.B(n_405),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_566),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_L g667 ( 
.A(n_571),
.B(n_185),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_517),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_571),
.B(n_191),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_440),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_547),
.A2(n_322),
.B(n_315),
.C(n_342),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_468),
.B(n_405),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_446),
.A2(n_322),
.B(n_342),
.C(n_341),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_449),
.B(n_193),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_494),
.A2(n_232),
.B1(n_323),
.B2(n_341),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_523),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_563),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_488),
.B(n_416),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_454),
.B(n_206),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_488),
.B(n_416),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_458),
.B(n_232),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_463),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_463),
.B(n_471),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_464),
.A2(n_214),
.B1(n_196),
.B2(n_261),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_542),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_524),
.B(n_197),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_463),
.B(n_416),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_529),
.A2(n_496),
.B1(n_500),
.B2(n_524),
.Y(n_688)
);

AND2x2_ASAP7_75t_SL g689 ( 
.A(n_530),
.B(n_316),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_471),
.B(n_389),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_471),
.B(n_389),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_475),
.B(n_208),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_564),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_547),
.B(n_389),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_436),
.B(n_437),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_522),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_475),
.B(n_207),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_436),
.B(n_389),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_433),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_554),
.B(n_212),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_435),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_436),
.B(n_389),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_508),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_437),
.B(n_211),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_523),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_R g706 ( 
.A(n_567),
.B(n_213),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_523),
.B(n_216),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_527),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_437),
.B(n_220),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_564),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_483),
.B(n_218),
.C(n_287),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_564),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_556),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_499),
.Y(n_714)
);

BUFx12f_ASAP7_75t_SL g715 ( 
.A(n_480),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_438),
.B(n_225),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_527),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_527),
.B(n_232),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_525),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_438),
.B(n_227),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_537),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_528),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_528),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_528),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_556),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_532),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_571),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_532),
.B(n_232),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_532),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_536),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_536),
.B(n_318),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_536),
.B(n_221),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_539),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_480),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_539),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_438),
.B(n_243),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_539),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_540),
.B(n_162),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_441),
.B(n_319),
.Y(n_739)
);

NOR3xp33_ASAP7_75t_SL g740 ( 
.A(n_586),
.B(n_241),
.C(n_222),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_655),
.B(n_544),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_731),
.Y(n_742)
);

AND2x6_ASAP7_75t_L g743 ( 
.A(n_637),
.B(n_540),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_663),
.B(n_319),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_612),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_637),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_688),
.B(n_466),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_596),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_731),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_623),
.B(n_544),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_623),
.B(n_548),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_637),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_575),
.B(n_548),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_576),
.A2(n_549),
.B1(n_546),
.B2(n_540),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_594),
.B(n_320),
.Y(n_755)
);

INVx5_ASAP7_75t_L g756 ( 
.A(n_734),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_605),
.B(n_447),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_635),
.B(n_320),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_619),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_703),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_676),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_595),
.A2(n_591),
.B1(n_579),
.B2(n_689),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_598),
.B(n_515),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_637),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_705),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_666),
.B(n_551),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_591),
.B(n_447),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_697),
.A2(n_546),
.B1(n_549),
.B2(n_558),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_596),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_608),
.Y(n_770)
);

CKINVDCx8_ASAP7_75t_R g771 ( 
.A(n_610),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_SL g772 ( 
.A1(n_595),
.A2(n_276),
.B1(n_275),
.B2(n_272),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_608),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_651),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_598),
.B(n_515),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_626),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_666),
.B(n_555),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_651),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_641),
.B(n_447),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_685),
.A2(n_516),
.B1(n_518),
.B2(n_519),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_714),
.B(n_555),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_648),
.B(n_558),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_644),
.B(n_561),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_672),
.B(n_561),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_708),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_678),
.B(n_562),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_641),
.B(n_323),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_658),
.B(n_447),
.Y(n_788)
);

INVx5_ASAP7_75t_L g789 ( 
.A(n_734),
.Y(n_789)
);

BUFx8_ASAP7_75t_L g790 ( 
.A(n_630),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_636),
.A2(n_516),
.B1(n_518),
.B2(n_519),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_717),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_723),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_629),
.B(n_466),
.Y(n_794)
);

BUFx4f_ASAP7_75t_L g795 ( 
.A(n_598),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_726),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_664),
.B(n_325),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_718),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_626),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_689),
.B(n_466),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_680),
.B(n_562),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_577),
.B(n_466),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_729),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_628),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_628),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_582),
.B(n_435),
.Y(n_806)
);

BUFx4f_ASAP7_75t_L g807 ( 
.A(n_609),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_583),
.B(n_599),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_734),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_SL g810 ( 
.A1(n_658),
.A2(n_262),
.B1(n_258),
.B2(n_255),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_730),
.Y(n_811)
);

AO22x1_ASAP7_75t_L g812 ( 
.A1(n_674),
.A2(n_264),
.B1(n_244),
.B2(n_263),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_735),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_737),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_643),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_604),
.B(n_435),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_664),
.B(n_325),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_589),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_606),
.B(n_428),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_679),
.B(n_466),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_643),
.Y(n_821)
);

AND2x6_ASAP7_75t_SL g822 ( 
.A(n_679),
.B(n_326),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_613),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_681),
.B(n_428),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_SL g825 ( 
.A1(n_675),
.A2(n_251),
.B1(n_246),
.B2(n_248),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_677),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_706),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_728),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_706),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_607),
.B(n_434),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_697),
.A2(n_571),
.B1(n_531),
.B2(n_444),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_638),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_739),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_677),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_621),
.A2(n_627),
.B(n_593),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_734),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_620),
.B(n_434),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_624),
.B(n_443),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_670),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_670),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_700),
.B(n_443),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_682),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_668),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_625),
.B(n_444),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_682),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_646),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_656),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_683),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_630),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_671),
.A2(n_572),
.B(n_568),
.C(n_459),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_657),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_693),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_631),
.B(n_445),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_609),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_693),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_597),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_611),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_700),
.B(n_445),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_615),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_617),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_603),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_621),
.A2(n_627),
.B1(n_584),
.B2(n_602),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_633),
.B(n_452),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_600),
.B(n_452),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_713),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_696),
.B(n_675),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_601),
.B(n_327),
.Y(n_867)
);

XNOR2xp5_ASAP7_75t_L g868 ( 
.A(n_610),
.B(n_52),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_710),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_654),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_732),
.A2(n_571),
.B1(n_531),
.B2(n_476),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_722),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_610),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_634),
.B(n_457),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_639),
.B(n_457),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_707),
.A2(n_459),
.B1(n_476),
.B2(n_503),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_609),
.A2(n_239),
.B1(n_162),
.B2(n_571),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_585),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_710),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_715),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_724),
.B(n_481),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_732),
.B(n_327),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_707),
.A2(n_503),
.B1(n_498),
.B2(n_481),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_L g884 ( 
.A(n_652),
.B(n_515),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_722),
.Y(n_885)
);

NAND2x1p5_ASAP7_75t_L g886 ( 
.A(n_733),
.B(n_505),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_684),
.B(n_480),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_671),
.B(n_553),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_R g889 ( 
.A(n_653),
.B(n_505),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_713),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_711),
.B(n_660),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_725),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_622),
.B(n_490),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_738),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_632),
.B(n_490),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_652),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_580),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_662),
.Y(n_898)
);

AND2x6_ASAP7_75t_L g899 ( 
.A(n_694),
.B(n_441),
.Y(n_899)
);

INVx5_ASAP7_75t_L g900 ( 
.A(n_712),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_665),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_712),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_581),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_588),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_580),
.A2(n_441),
.B(n_442),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_652),
.B(n_497),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_587),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_590),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_687),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_614),
.Y(n_910)
);

OAI22xp33_ASAP7_75t_L g911 ( 
.A1(n_592),
.A2(n_442),
.B1(n_497),
.B2(n_498),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_738),
.Y(n_912)
);

AND2x6_ASAP7_75t_SL g913 ( 
.A(n_704),
.B(n_298),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_647),
.B(n_482),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_647),
.B(n_482),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_652),
.B(n_593),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_650),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_699),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_661),
.B(n_300),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_856),
.B(n_661),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_896),
.A2(n_692),
.B(n_645),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_896),
.A2(n_692),
.B(n_649),
.Y(n_922)
);

OAI21x1_ASAP7_75t_L g923 ( 
.A1(n_905),
.A2(n_695),
.B(n_616),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_762),
.A2(n_686),
.B(n_673),
.C(n_642),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_787),
.B(n_686),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_884),
.A2(n_616),
.B(n_618),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_L g927 ( 
.A(n_762),
.B(n_719),
.C(n_721),
.Y(n_927)
);

OAI21xp33_ASAP7_75t_L g928 ( 
.A1(n_755),
.A2(n_618),
.B(n_640),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_782),
.A2(n_727),
.B1(n_690),
.B2(n_691),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_763),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_759),
.B(n_640),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_756),
.A2(n_515),
.B(n_578),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_880),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_828),
.B(n_652),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_756),
.A2(n_515),
.B(n_669),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_905),
.A2(n_698),
.B(n_702),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_767),
.A2(n_736),
.B(n_720),
.C(n_716),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_742),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_760),
.Y(n_939)
);

O2A1O1Ixp5_ASAP7_75t_L g940 ( 
.A1(n_841),
.A2(n_858),
.B(n_887),
.C(n_914),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_824),
.A2(n_709),
.B(n_701),
.C(n_667),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_756),
.A2(n_659),
.B(n_482),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_854),
.B(n_442),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_882),
.B(n_828),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_798),
.B(n_239),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_SL g946 ( 
.A1(n_747),
.A2(n_489),
.B(n_451),
.C(n_448),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_846),
.B(n_652),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_746),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_847),
.B(n_448),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_854),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_749),
.Y(n_951)
);

AOI33xp33_ASAP7_75t_L g952 ( 
.A1(n_744),
.A2(n_572),
.A3(n_568),
.B1(n_511),
.B2(n_506),
.B3(n_495),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_857),
.A2(n_571),
.B1(n_239),
.B2(n_487),
.Y(n_953)
);

OAI22x1_ASAP7_75t_L g954 ( 
.A1(n_868),
.A2(n_511),
.B1(n_448),
.B2(n_450),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_840),
.B(n_505),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_745),
.B(n_827),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_756),
.A2(n_482),
.B(n_514),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_829),
.B(n_505),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_778),
.B(n_482),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_890),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_835),
.A2(n_489),
.B(n_450),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_782),
.A2(n_572),
.B1(n_568),
.B2(n_511),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_789),
.A2(n_514),
.B(n_507),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_865),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_750),
.A2(n_451),
.B1(n_450),
.B2(n_461),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_894),
.A2(n_487),
.B(n_451),
.C(n_461),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_850),
.A2(n_489),
.B(n_465),
.Y(n_967)
);

AOI21x1_ASAP7_75t_L g968 ( 
.A1(n_820),
.A2(n_486),
.B(n_465),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_890),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_892),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_766),
.B(n_467),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_789),
.A2(n_514),
.B(n_507),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_854),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_851),
.B(n_492),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_746),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_750),
.A2(n_491),
.B1(n_467),
.B2(n_470),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_866),
.B(n_510),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_SL g978 ( 
.A1(n_772),
.A2(n_239),
.B1(n_2),
.B2(n_5),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_859),
.B(n_492),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_860),
.B(n_492),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_746),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_840),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_751),
.A2(n_486),
.B1(n_467),
.B2(n_470),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_797),
.B(n_495),
.Y(n_984)
);

O2A1O1Ixp5_ASAP7_75t_L g985 ( 
.A1(n_915),
.A2(n_495),
.B(n_477),
.C(n_486),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_748),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_808),
.B(n_506),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_751),
.A2(n_491),
.B1(n_470),
.B2(n_506),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_761),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_769),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_836),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_789),
.A2(n_514),
.B(n_510),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_765),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_808),
.A2(n_878),
.B(n_907),
.C(n_912),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_822),
.B(n_507),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_788),
.A2(n_477),
.B(n_491),
.C(n_510),
.Y(n_996)
);

NOR2x1_ASAP7_75t_L g997 ( 
.A(n_774),
.B(n_477),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_864),
.A2(n_510),
.B(n_2),
.C(n_5),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_836),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_797),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_810),
.B(n_757),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_862),
.A2(n_460),
.B1(n_473),
.B2(n_8),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_835),
.A2(n_779),
.B(n_901),
.C(n_898),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_778),
.B(n_553),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_781),
.A2(n_0),
.B(n_6),
.C(n_15),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_817),
.B(n_19),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_770),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_817),
.B(n_23),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_785),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_SL g1010 ( 
.A(n_740),
.B(n_877),
.C(n_771),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_SL g1011 ( 
.A1(n_916),
.A2(n_76),
.B(n_135),
.C(n_133),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_766),
.B(n_553),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_789),
.A2(n_553),
.B(n_473),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_792),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_916),
.A2(n_460),
.B1(n_473),
.B2(n_29),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_793),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_777),
.B(n_23),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_777),
.B(n_24),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_836),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_809),
.A2(n_553),
.B(n_473),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_781),
.B(n_24),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_773),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_818),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_783),
.A2(n_473),
.B1(n_460),
.B2(n_33),
.Y(n_1024)
);

BUFx4f_ASAP7_75t_L g1025 ( 
.A(n_778),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_758),
.A2(n_31),
.B(n_32),
.Y(n_1026)
);

OR2x6_ASAP7_75t_L g1027 ( 
.A(n_763),
.B(n_460),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_840),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_913),
.B(n_34),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_919),
.A2(n_833),
.B(n_909),
.C(n_891),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_SL g1031 ( 
.A(n_873),
.B(n_34),
.C(n_35),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_867),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_850),
.A2(n_88),
.B(n_130),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_796),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_803),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_823),
.A2(n_35),
.B(n_39),
.C(n_40),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_SL g1037 ( 
.A(n_877),
.B(n_39),
.C(n_40),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_776),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_867),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_812),
.B(n_42),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_842),
.Y(n_1041)
);

BUFx4f_ASAP7_75t_L g1042 ( 
.A(n_870),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_758),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_799),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_790),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_774),
.A2(n_95),
.B1(n_57),
.B2(n_67),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_783),
.B(n_44),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_861),
.B(n_125),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_832),
.A2(n_73),
.B(n_92),
.C(n_102),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_R g1050 ( 
.A(n_849),
.B(n_104),
.Y(n_1050)
);

CKINVDCx16_ASAP7_75t_R g1051 ( 
.A(n_825),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_842),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_843),
.B(n_120),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_842),
.B(n_809),
.Y(n_1054)
);

BUFx4f_ASAP7_75t_L g1055 ( 
.A(n_763),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_809),
.A2(n_753),
.B(n_906),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_848),
.B(n_800),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_775),
.B(n_752),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_804),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_809),
.A2(n_753),
.B(n_906),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_930),
.Y(n_1061)
);

AO31x2_ASAP7_75t_L g1062 ( 
.A1(n_1030),
.A2(n_897),
.A3(n_784),
.B(n_786),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_967),
.A2(n_895),
.B(n_893),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_940),
.A2(n_784),
.B(n_801),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_922),
.A2(n_845),
.B(n_839),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_944),
.B(n_741),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_925),
.B(n_741),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_987),
.B(n_819),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_926),
.A2(n_845),
.B(n_839),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_936),
.A2(n_895),
.B(n_893),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1043),
.B(n_807),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_923),
.A2(n_806),
.B(n_768),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_986),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_SL g1074 ( 
.A(n_939),
.B(n_900),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_989),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_924),
.A2(n_1001),
.B(n_927),
.C(n_920),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_993),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_933),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1009),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1003),
.A2(n_801),
.B(n_786),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1014),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1025),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_968),
.A2(n_806),
.B(n_874),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_1025),
.Y(n_1084)
);

AND2x2_ASAP7_75t_SL g1085 ( 
.A(n_1051),
.B(n_807),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_937),
.A2(n_816),
.B(n_830),
.Y(n_1086)
);

O2A1O1Ixp5_ASAP7_75t_L g1087 ( 
.A1(n_1033),
.A2(n_911),
.B(n_802),
.C(n_830),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_921),
.A2(n_853),
.B(n_874),
.Y(n_1088)
);

OAI22x1_ASAP7_75t_L g1089 ( 
.A1(n_1040),
.A2(n_1018),
.B1(n_1017),
.B2(n_1029),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_1000),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1021),
.B(n_848),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_961),
.A2(n_985),
.B(n_976),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_1032),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_991),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1006),
.B(n_1008),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_961),
.A2(n_976),
.B(n_965),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_965),
.A2(n_875),
.B(n_837),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1033),
.A2(n_780),
.B(n_795),
.C(n_791),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1050),
.Y(n_1099)
);

AO21x1_ASAP7_75t_L g1100 ( 
.A1(n_1002),
.A2(n_819),
.B(n_897),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1002),
.A2(n_1016),
.B1(n_1035),
.B2(n_1034),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_983),
.A2(n_853),
.B(n_875),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_983),
.A2(n_844),
.B(n_863),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_931),
.B(n_848),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_996),
.A2(n_863),
.B(n_837),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_988),
.A2(n_844),
.B(n_838),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_SL g1107 ( 
.A1(n_998),
.A2(n_1049),
.B(n_1037),
.C(n_934),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_988),
.A2(n_838),
.B(n_886),
.Y(n_1108)
);

CKINVDCx11_ASAP7_75t_R g1109 ( 
.A(n_1045),
.Y(n_1109)
);

INVx5_ASAP7_75t_SL g1110 ( 
.A(n_950),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_945),
.B(n_1039),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_942),
.A2(n_886),
.B(n_881),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_956),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_964),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_941),
.A2(n_816),
.B(n_831),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1056),
.A2(n_900),
.B(n_872),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_938),
.B(n_811),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1057),
.B(n_814),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_994),
.B(n_752),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_966),
.A2(n_813),
.A3(n_881),
.B(n_821),
.Y(n_1120)
);

OAI22x1_ASAP7_75t_L g1121 ( 
.A1(n_995),
.A2(n_764),
.B1(n_888),
.B2(n_876),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_929),
.A2(n_754),
.B(n_899),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1042),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1047),
.B(n_764),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_950),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_928),
.A2(n_795),
.B(n_871),
.C(n_883),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_990),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_977),
.B(n_885),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1060),
.A2(n_879),
.B(n_869),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_970),
.Y(n_1130)
);

OR2x2_ASAP7_75t_L g1131 ( 
.A(n_951),
.B(n_917),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_SL g1132 ( 
.A(n_1023),
.B(n_889),
.C(n_794),
.Y(n_1132)
);

AO32x2_ASAP7_75t_L g1133 ( 
.A1(n_1024),
.A2(n_899),
.A3(n_743),
.B1(n_900),
.B2(n_805),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1007),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1053),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_962),
.A2(n_826),
.B(n_852),
.Y(n_1136)
);

AOI211x1_ASAP7_75t_L g1137 ( 
.A1(n_1026),
.A2(n_888),
.B(n_899),
.C(n_790),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_929),
.A2(n_899),
.B(n_902),
.Y(n_1138)
);

OAI21xp33_ASAP7_75t_L g1139 ( 
.A1(n_1036),
.A2(n_918),
.B(n_904),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_971),
.B(n_885),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_973),
.B(n_775),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1022),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_962),
.A2(n_815),
.B(n_834),
.Y(n_1143)
);

NAND3xp33_ASAP7_75t_L g1144 ( 
.A(n_1005),
.B(n_908),
.C(n_903),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1038),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_1024),
.A2(n_855),
.A3(n_899),
.B(n_743),
.Y(n_1146)
);

AO32x2_ASAP7_75t_L g1147 ( 
.A1(n_1015),
.A2(n_743),
.A3(n_900),
.B1(n_910),
.B2(n_872),
.Y(n_1147)
);

OR2x6_ASAP7_75t_L g1148 ( 
.A(n_1041),
.B(n_775),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1044),
.Y(n_1149)
);

AO22x2_ASAP7_75t_L g1150 ( 
.A1(n_1010),
.A2(n_910),
.B1(n_743),
.B2(n_872),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_973),
.B(n_872),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_947),
.A2(n_1015),
.B(n_974),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_935),
.A2(n_932),
.B(n_997),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1059),
.Y(n_1154)
);

O2A1O1Ixp5_ASAP7_75t_SL g1155 ( 
.A1(n_959),
.A2(n_981),
.B(n_948),
.C(n_975),
.Y(n_1155)
);

AO32x2_ASAP7_75t_L g1156 ( 
.A1(n_978),
.A2(n_952),
.A3(n_954),
.B1(n_1041),
.B2(n_946),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_949),
.B(n_980),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_979),
.B(n_969),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_R g1159 ( 
.A(n_973),
.B(n_982),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_960),
.B(n_958),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_930),
.Y(n_1161)
);

AND3x4_ASAP7_75t_L g1162 ( 
.A(n_1031),
.B(n_1058),
.C(n_984),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_991),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1042),
.B(n_943),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_SL g1165 ( 
.A(n_930),
.B(n_1027),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_943),
.B(n_1052),
.Y(n_1166)
);

OAI21xp33_ASAP7_75t_L g1167 ( 
.A1(n_1046),
.A2(n_953),
.B(n_1048),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1012),
.B(n_1058),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_963),
.A2(n_972),
.B(n_992),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_948),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_975),
.B(n_981),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_991),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_957),
.A2(n_955),
.B(n_1020),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_955),
.A2(n_1013),
.B(n_1054),
.Y(n_1174)
);

OAI22x1_ASAP7_75t_L g1175 ( 
.A1(n_982),
.A2(n_1052),
.B1(n_1028),
.B2(n_1004),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1028),
.B(n_999),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1055),
.A2(n_1011),
.B1(n_1027),
.B2(n_1019),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1055),
.B(n_999),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_999),
.B(n_1019),
.C(n_1027),
.Y(n_1179)
);

BUFx2_ASAP7_75t_SL g1180 ( 
.A(n_1019),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_989),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1030),
.A2(n_762),
.B(n_591),
.C(n_535),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1025),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1043),
.B(n_854),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_940),
.A2(n_1033),
.B(n_1030),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_922),
.A2(n_896),
.B(n_884),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1030),
.A2(n_996),
.A3(n_1003),
.B(n_966),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1030),
.A2(n_996),
.A3(n_1003),
.B(n_966),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_930),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_933),
.Y(n_1190)
);

OAI22x1_ASAP7_75t_L g1191 ( 
.A1(n_1001),
.A2(n_688),
.B1(n_591),
.B2(n_595),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_920),
.B(n_594),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1030),
.A2(n_762),
.B(n_591),
.C(n_535),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_939),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1001),
.A2(n_762),
.B1(n_591),
.B2(n_595),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_925),
.B(n_762),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_930),
.B(n_1055),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1025),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_922),
.A2(n_896),
.B(n_884),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_944),
.B(n_787),
.Y(n_1200)
);

AOI221x1_ASAP7_75t_L g1201 ( 
.A1(n_927),
.A2(n_762),
.B1(n_1033),
.B2(n_1037),
.C(n_998),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_967),
.A2(n_936),
.B(n_923),
.Y(n_1202)
);

BUFx10_ASAP7_75t_L g1203 ( 
.A(n_939),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1000),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1201),
.A2(n_1076),
.A3(n_1121),
.B(n_1100),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1202),
.A2(n_1153),
.B(n_1169),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1186),
.A2(n_1199),
.B(n_1112),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1195),
.B(n_1111),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1090),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1195),
.A2(n_1193),
.B(n_1182),
.C(n_1098),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1086),
.A2(n_1065),
.B(n_1068),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1070),
.A2(n_1173),
.B(n_1129),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1069),
.A2(n_1088),
.B(n_1063),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1141),
.B(n_1148),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1075),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1136),
.A2(n_1143),
.B(n_1083),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1167),
.A2(n_1087),
.B(n_1196),
.Y(n_1217)
);

BUFx12f_ASAP7_75t_L g1218 ( 
.A(n_1109),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1066),
.B(n_1067),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1077),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1079),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1167),
.A2(n_1196),
.B(n_1152),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1116),
.A2(n_1108),
.B(n_1072),
.Y(n_1223)
);

BUFx8_ASAP7_75t_L g1224 ( 
.A(n_1183),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1081),
.Y(n_1225)
);

AO21x2_ASAP7_75t_L g1226 ( 
.A1(n_1138),
.A2(n_1122),
.B(n_1064),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1092),
.A2(n_1115),
.B(n_1097),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1102),
.A2(n_1106),
.B(n_1103),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1126),
.A2(n_1191),
.A3(n_1089),
.B(n_1101),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_1113),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1096),
.A2(n_1138),
.B(n_1122),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1174),
.A2(n_1080),
.B(n_1064),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1119),
.A2(n_1150),
.B(n_1124),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1181),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1117),
.Y(n_1235)
);

OR2x6_ASAP7_75t_L g1236 ( 
.A(n_1197),
.B(n_1137),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1190),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1114),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_1183),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1093),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_1194),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1183),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1067),
.B(n_1135),
.Y(n_1243)
);

O2A1O1Ixp5_ASAP7_75t_L g1244 ( 
.A1(n_1152),
.A2(n_1080),
.B(n_1101),
.C(n_1178),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1155),
.A2(n_1105),
.B(n_1185),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1130),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1131),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1099),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1135),
.A2(n_1185),
.B1(n_1085),
.B2(n_1118),
.Y(n_1249)
);

BUFx12f_ASAP7_75t_L g1250 ( 
.A(n_1203),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1120),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1145),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1105),
.A2(n_1168),
.B(n_1128),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1149),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1168),
.A2(n_1157),
.B(n_1177),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1157),
.A2(n_1177),
.B(n_1068),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1120),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_1104),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_1203),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1118),
.A2(n_1091),
.B1(n_1162),
.B2(n_1104),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1154),
.Y(n_1261)
);

NOR2x1_ASAP7_75t_L g1262 ( 
.A(n_1179),
.B(n_1061),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1078),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1132),
.A2(n_1139),
.B1(n_1144),
.B2(n_1204),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1144),
.A2(n_1107),
.B(n_1160),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1071),
.A2(n_1164),
.B1(n_1204),
.B2(n_1184),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1161),
.A2(n_1189),
.B(n_1197),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1141),
.B(n_1148),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1158),
.A2(n_1140),
.B(n_1139),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1123),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1158),
.A2(n_1179),
.B(n_1160),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1120),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1082),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1146),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1084),
.A2(n_1150),
.B1(n_1184),
.B2(n_1198),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1148),
.B(n_1166),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1073),
.B(n_1127),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1134),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1142),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1165),
.A2(n_1198),
.B1(n_1147),
.B2(n_1110),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1094),
.Y(n_1281)
);

CKINVDCx16_ASAP7_75t_R g1282 ( 
.A(n_1159),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_SL g1283 ( 
.A1(n_1171),
.A2(n_1176),
.B(n_1170),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1062),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1125),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1163),
.B(n_1172),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1176),
.A2(n_1188),
.B(n_1187),
.Y(n_1287)
);

BUFx4f_ASAP7_75t_SL g1288 ( 
.A(n_1163),
.Y(n_1288)
);

AO22x1_ASAP7_75t_SL g1289 ( 
.A1(n_1151),
.A2(n_1074),
.B1(n_1156),
.B2(n_1110),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1094),
.B(n_1175),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1133),
.A2(n_1147),
.A3(n_1062),
.B(n_1146),
.Y(n_1291)
);

CKINVDCx11_ASAP7_75t_R g1292 ( 
.A(n_1180),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1094),
.B(n_1062),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1147),
.A2(n_1133),
.B(n_1146),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1187),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1188),
.B(n_1156),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1195),
.A2(n_762),
.B1(n_1076),
.B2(n_1001),
.Y(n_1297)
);

AND2x4_ASAP7_75t_SL g1298 ( 
.A(n_1203),
.B(n_1183),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1192),
.B(n_1200),
.Y(n_1299)
);

BUFx8_ASAP7_75t_SL g1300 ( 
.A(n_1194),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1195),
.A2(n_1193),
.B(n_1182),
.C(n_762),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1203),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1075),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1095),
.B(n_594),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1195),
.A2(n_1051),
.B1(n_1113),
.B2(n_978),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1104),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1075),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1192),
.B(n_1200),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1195),
.A2(n_1191),
.B1(n_762),
.B2(n_1201),
.Y(n_1309)
);

NOR2x1_ASAP7_75t_L g1310 ( 
.A(n_1113),
.B(n_1179),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1202),
.A2(n_1153),
.B(n_1169),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1076),
.A2(n_1195),
.B(n_641),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1200),
.B(n_1066),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1195),
.A2(n_762),
.B1(n_1076),
.B2(n_1001),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1195),
.B(n_762),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1075),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1195),
.B(n_762),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1075),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1136),
.Y(n_1319)
);

NAND3xp33_ASAP7_75t_SL g1320 ( 
.A(n_1195),
.B(n_1076),
.C(n_1182),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1096),
.A2(n_1092),
.B(n_1201),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1200),
.B(n_1066),
.Y(n_1322)
);

OR2x4_ASAP7_75t_L g1323 ( 
.A(n_1183),
.B(n_1010),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1075),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1203),
.Y(n_1325)
);

INVx5_ASAP7_75t_L g1326 ( 
.A(n_1183),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1075),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1153),
.A2(n_1202),
.B(n_1065),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1113),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1136),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1075),
.Y(n_1331)
);

O2A1O1Ixp5_ASAP7_75t_L g1332 ( 
.A1(n_1312),
.A2(n_1314),
.B(n_1297),
.C(n_1309),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1315),
.B(n_1317),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1315),
.B(n_1317),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1225),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1208),
.B(n_1296),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1296),
.B(n_1229),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1320),
.A2(n_1210),
.B(n_1309),
.C(n_1301),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1313),
.B(n_1322),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1306),
.B(n_1258),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1296),
.B(n_1229),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1219),
.B(n_1243),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1230),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1236),
.B(n_1214),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1258),
.B(n_1299),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1237),
.Y(n_1346)
);

AOI21x1_ASAP7_75t_SL g1347 ( 
.A1(n_1293),
.A2(n_1295),
.B(n_1304),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1236),
.B(n_1214),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1305),
.A2(n_1260),
.B1(n_1323),
.B2(n_1266),
.Y(n_1349)
);

O2A1O1Ixp5_ASAP7_75t_L g1350 ( 
.A1(n_1217),
.A2(n_1222),
.B(n_1301),
.C(n_1244),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1308),
.B(n_1306),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1235),
.B(n_1247),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1229),
.B(n_1205),
.Y(n_1353)
);

AOI21x1_ASAP7_75t_SL g1354 ( 
.A1(n_1268),
.A2(n_1274),
.B(n_1276),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1277),
.B(n_1209),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1240),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1229),
.B(n_1205),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1209),
.B(n_1278),
.Y(n_1358)
);

NOR2xp67_ASAP7_75t_L g1359 ( 
.A(n_1302),
.B(n_1325),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1245),
.A2(n_1228),
.B(n_1227),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1361)
);

NAND2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1262),
.B(n_1256),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1265),
.A2(n_1275),
.B(n_1264),
.C(n_1283),
.Y(n_1363)
);

NOR2xp67_ASAP7_75t_L g1364 ( 
.A(n_1250),
.B(n_1270),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1268),
.A2(n_1274),
.B(n_1276),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1245),
.A2(n_1216),
.B(n_1213),
.Y(n_1366)
);

O2A1O1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1264),
.A2(n_1310),
.B(n_1303),
.C(n_1307),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1281),
.A2(n_1268),
.B(n_1276),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1323),
.A2(n_1249),
.B1(n_1282),
.B2(n_1259),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1249),
.A2(n_1259),
.B1(n_1273),
.B2(n_1288),
.Y(n_1370)
);

O2A1O1Ixp5_ASAP7_75t_L g1371 ( 
.A1(n_1233),
.A2(n_1284),
.B(n_1272),
.C(n_1257),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1205),
.B(n_1215),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1236),
.B(n_1267),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1280),
.A2(n_1255),
.B(n_1271),
.C(n_1253),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1224),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1286),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1220),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1329),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_SL g1379 ( 
.A1(n_1289),
.A2(n_1250),
.B(n_1280),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1205),
.B(n_1331),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1273),
.A2(n_1288),
.B1(n_1263),
.B2(n_1290),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1221),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1287),
.B(n_1226),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1234),
.Y(n_1384)
);

O2A1O1Ixp5_ASAP7_75t_L g1385 ( 
.A1(n_1284),
.A2(n_1251),
.B(n_1257),
.C(n_1272),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1238),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1279),
.B(n_1261),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1207),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1285),
.Y(n_1389)
);

NOR2xp67_ASAP7_75t_L g1390 ( 
.A(n_1252),
.B(n_1254),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1271),
.A2(n_1269),
.B(n_1287),
.C(n_1318),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1231),
.B(n_1321),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1246),
.A2(n_1327),
.B(n_1324),
.C(n_1316),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1223),
.A2(n_1212),
.B(n_1206),
.Y(n_1394)
);

O2A1O1Ixp5_ASAP7_75t_L g1395 ( 
.A1(n_1319),
.A2(n_1330),
.B(n_1290),
.C(n_1231),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1212),
.A2(n_1206),
.B(n_1311),
.Y(n_1396)
);

AOI21x1_ASAP7_75t_SL g1397 ( 
.A1(n_1292),
.A2(n_1218),
.B(n_1224),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1263),
.A2(n_1326),
.B1(n_1239),
.B2(n_1298),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1300),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1242),
.B(n_1239),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1321),
.B(n_1294),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1239),
.A2(n_1326),
.B1(n_1242),
.B2(n_1241),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1321),
.B(n_1294),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1326),
.A2(n_1242),
.B1(n_1241),
.B2(n_1281),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1242),
.B(n_1224),
.Y(n_1405)
);

CKINVDCx16_ASAP7_75t_R g1406 ( 
.A(n_1218),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1292),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1248),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1281),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1281),
.A2(n_1248),
.B1(n_1330),
.B2(n_1300),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1291),
.B(n_1328),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1291),
.A2(n_1195),
.B1(n_1113),
.B2(n_1305),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1312),
.A2(n_1211),
.B(n_1297),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1225),
.Y(n_1414)
);

O2A1O1Ixp5_ASAP7_75t_L g1415 ( 
.A1(n_1312),
.A2(n_1297),
.B(n_1314),
.C(n_1309),
.Y(n_1415)
);

AOI21x1_ASAP7_75t_SL g1416 ( 
.A1(n_1293),
.A2(n_576),
.B(n_579),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1312),
.A2(n_1076),
.B(n_762),
.C(n_1297),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1315),
.B(n_1317),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1313),
.B(n_1322),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1312),
.A2(n_1195),
.B(n_1193),
.C(n_1182),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1312),
.A2(n_1076),
.B(n_762),
.C(n_1297),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1313),
.B(n_1322),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1315),
.B(n_1317),
.Y(n_1423)
);

BUFx4f_ASAP7_75t_SL g1424 ( 
.A(n_1218),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1225),
.Y(n_1425)
);

OAI31xp33_ASAP7_75t_L g1426 ( 
.A1(n_1297),
.A2(n_636),
.A3(n_1076),
.B(n_978),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1313),
.B(n_1322),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1313),
.B(n_1322),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1315),
.B(n_1317),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1312),
.A2(n_1195),
.B(n_1193),
.C(n_1182),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1336),
.B(n_1337),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1372),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1380),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1343),
.B(n_1378),
.Y(n_1434)
);

CKINVDCx14_ASAP7_75t_R g1435 ( 
.A(n_1399),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1390),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1395),
.A2(n_1385),
.B(n_1371),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1413),
.A2(n_1430),
.B(n_1420),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1416),
.A2(n_1360),
.B(n_1366),
.Y(n_1439)
);

AO21x2_ASAP7_75t_L g1440 ( 
.A1(n_1420),
.A2(n_1430),
.B(n_1391),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1346),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1373),
.B(n_1344),
.Y(n_1442)
);

OAI211xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1426),
.A2(n_1338),
.B(n_1421),
.C(n_1417),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1332),
.A2(n_1415),
.B(n_1350),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1336),
.B(n_1337),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1391),
.A2(n_1374),
.B(n_1392),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1373),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1401),
.A2(n_1403),
.B(n_1357),
.Y(n_1448)
);

NAND2xp33_ASAP7_75t_SL g1449 ( 
.A(n_1399),
.B(n_1349),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1335),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1411),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1414),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1425),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1377),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1333),
.B(n_1334),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1341),
.B(n_1353),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1341),
.B(n_1353),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1382),
.Y(n_1458)
);

OR2x6_ASAP7_75t_L g1459 ( 
.A(n_1368),
.B(n_1344),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1384),
.Y(n_1460)
);

OR2x6_ASAP7_75t_L g1461 ( 
.A(n_1344),
.B(n_1348),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1348),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1386),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1393),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1387),
.Y(n_1465)
);

OR2x6_ASAP7_75t_L g1466 ( 
.A(n_1348),
.B(n_1362),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1340),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1361),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1383),
.A2(n_1363),
.B(n_1345),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1351),
.B(n_1376),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1358),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1388),
.A2(n_1429),
.B(n_1334),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1333),
.B(n_1429),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1418),
.B(n_1423),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1418),
.B(n_1423),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1356),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1352),
.Y(n_1477)
);

BUFx12f_ASAP7_75t_L g1478 ( 
.A(n_1375),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1367),
.B(n_1404),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1412),
.A2(n_1339),
.B1(n_1427),
.B2(n_1422),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1396),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1370),
.A2(n_1369),
.B(n_1360),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1355),
.B(n_1342),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1451),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1447),
.B(n_1375),
.Y(n_1485)
);

AOI21xp33_ASAP7_75t_L g1486 ( 
.A1(n_1438),
.A2(n_1428),
.B(n_1419),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1458),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1458),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1431),
.B(n_1394),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1448),
.B(n_1389),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1445),
.B(n_1394),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1471),
.B(n_1409),
.Y(n_1492)
);

AOI211x1_ASAP7_75t_L g1493 ( 
.A1(n_1480),
.A2(n_1381),
.B(n_1410),
.C(n_1405),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1478),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1478),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1448),
.B(n_1396),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1454),
.Y(n_1497)
);

AND2x4_ASAP7_75t_SL g1498 ( 
.A(n_1459),
.B(n_1354),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1432),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1467),
.B(n_1359),
.Y(n_1500)
);

AOI222xp33_ASAP7_75t_L g1501 ( 
.A1(n_1443),
.A2(n_1424),
.B1(n_1408),
.B2(n_1407),
.C1(n_1364),
.C2(n_1402),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1456),
.B(n_1400),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1448),
.B(n_1398),
.Y(n_1503)
);

NOR2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1464),
.B(n_1379),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1448),
.B(n_1406),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1459),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1467),
.B(n_1347),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1469),
.B(n_1365),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1456),
.B(n_1457),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1457),
.B(n_1397),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1447),
.Y(n_1511)
);

NAND4xp25_ASAP7_75t_L g1512 ( 
.A(n_1493),
.B(n_1443),
.C(n_1444),
.D(n_1480),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1490),
.B(n_1470),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1504),
.A2(n_1438),
.B1(n_1449),
.B2(n_1440),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1502),
.B(n_1442),
.Y(n_1515)
);

OAI31xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1510),
.A2(n_1442),
.A3(n_1476),
.B(n_1441),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1508),
.A2(n_1481),
.B(n_1472),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1484),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_R g1519 ( 
.A(n_1494),
.B(n_1435),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1493),
.A2(n_1479),
.B1(n_1444),
.B2(n_1459),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1506),
.B(n_1459),
.Y(n_1521)
);

INVx4_ASAP7_75t_L g1522 ( 
.A(n_1494),
.Y(n_1522)
);

OAI211xp5_ASAP7_75t_L g1523 ( 
.A1(n_1486),
.A2(n_1508),
.B(n_1501),
.C(n_1505),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1497),
.B(n_1483),
.Y(n_1524)
);

NAND2x1_ASAP7_75t_L g1525 ( 
.A(n_1511),
.B(n_1459),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1487),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1504),
.A2(n_1438),
.B1(n_1440),
.B2(n_1479),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1494),
.Y(n_1528)
);

OAI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1505),
.A2(n_1479),
.B1(n_1441),
.B2(n_1476),
.C(n_1436),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1500),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1500),
.A2(n_1479),
.B1(n_1461),
.B2(n_1473),
.Y(n_1531)
);

BUFx4f_ASAP7_75t_L g1532 ( 
.A(n_1485),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1492),
.B(n_1483),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1501),
.A2(n_1479),
.B1(n_1440),
.B2(n_1442),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1488),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1484),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1506),
.B(n_1466),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1506),
.B(n_1447),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1509),
.B(n_1462),
.Y(n_1539)
);

OAI33xp33_ASAP7_75t_L g1540 ( 
.A1(n_1507),
.A2(n_1463),
.A3(n_1460),
.B1(n_1477),
.B2(n_1433),
.B3(n_1432),
.Y(n_1540)
);

AOI33xp33_ASAP7_75t_L g1541 ( 
.A1(n_1510),
.A2(n_1477),
.A3(n_1460),
.B1(n_1463),
.B2(n_1465),
.B3(n_1433),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1507),
.A2(n_1455),
.B1(n_1474),
.B2(n_1475),
.C(n_1465),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1499),
.Y(n_1543)
);

AOI33xp33_ASAP7_75t_L g1544 ( 
.A1(n_1498),
.A2(n_1468),
.A3(n_1475),
.B1(n_1452),
.B2(n_1450),
.B3(n_1453),
.Y(n_1544)
);

AOI222xp33_ASAP7_75t_L g1545 ( 
.A1(n_1498),
.A2(n_1424),
.B1(n_1434),
.B2(n_1474),
.C1(n_1455),
.C2(n_1468),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1525),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1512),
.A2(n_1498),
.B(n_1506),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1518),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1542),
.B(n_1491),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1537),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1536),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1527),
.A2(n_1482),
.B(n_1446),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1517),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1517),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1513),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1539),
.B(n_1509),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1526),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1532),
.Y(n_1558)
);

BUFx12f_ASAP7_75t_L g1559 ( 
.A(n_1522),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1538),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1521),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1535),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1541),
.B(n_1491),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1543),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1531),
.A2(n_1437),
.B(n_1439),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1541),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1544),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1538),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1523),
.B(n_1496),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1538),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1557),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1566),
.B(n_1567),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1560),
.B(n_1532),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1553),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1550),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1566),
.B(n_1530),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1553),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1567),
.B(n_1533),
.Y(n_1578)
);

INVx4_ASAP7_75t_L g1579 ( 
.A(n_1559),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1569),
.A2(n_1527),
.B1(n_1520),
.B2(n_1534),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1559),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1569),
.B(n_1524),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1550),
.B(n_1516),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1548),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1550),
.B(n_1489),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1553),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1564),
.B(n_1544),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1561),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1561),
.B(n_1537),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1557),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1553),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1554),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_L g1593 ( 
.A(n_1569),
.B(n_1522),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1557),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1537),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1562),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1560),
.B(n_1568),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1568),
.B(n_1515),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1563),
.B(n_1503),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1563),
.B(n_1469),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1559),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1562),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1561),
.B(n_1546),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1547),
.A2(n_1514),
.B(n_1529),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1568),
.B(n_1521),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1559),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1587),
.B(n_1549),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1597),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1583),
.B(n_1568),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1571),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1587),
.B(n_1549),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_SL g1612 ( 
.A1(n_1593),
.A2(n_1561),
.B1(n_1546),
.B2(n_1552),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1571),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1583),
.B(n_1570),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1590),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1572),
.B(n_1556),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1582),
.B(n_1555),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1590),
.Y(n_1618)
);

AOI211xp5_ASAP7_75t_L g1619 ( 
.A1(n_1604),
.A2(n_1547),
.B(n_1565),
.C(n_1558),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1594),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1594),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1596),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1603),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1593),
.B(n_1519),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1589),
.B(n_1570),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1584),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1572),
.B(n_1556),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1596),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1583),
.B(n_1570),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1576),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1579),
.B(n_1495),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1602),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1597),
.Y(n_1633)
);

A2O1A1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1604),
.A2(n_1514),
.B(n_1565),
.C(n_1558),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1575),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1602),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1573),
.B(n_1570),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1576),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1573),
.B(n_1546),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_L g1640 ( 
.A(n_1580),
.B(n_1545),
.C(n_1554),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_SL g1641 ( 
.A(n_1580),
.B(n_1519),
.C(n_1554),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1635),
.Y(n_1642)
);

AND2x2_ASAP7_75t_SL g1643 ( 
.A(n_1607),
.B(n_1579),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1641),
.A2(n_1600),
.B1(n_1575),
.B2(n_1578),
.C(n_1588),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1623),
.B(n_1589),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1617),
.Y(n_1646)
);

AOI222xp33_ASAP7_75t_L g1647 ( 
.A1(n_1630),
.A2(n_1578),
.B1(n_1600),
.B2(n_1588),
.C1(n_1540),
.C2(n_1581),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1626),
.B(n_1638),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1609),
.B(n_1581),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1617),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1609),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1614),
.B(n_1606),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1610),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1610),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1624),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1631),
.B(n_1579),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1616),
.B(n_1582),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1607),
.B(n_1579),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1614),
.Y(n_1659)
);

AOI22x1_ASAP7_75t_L g1660 ( 
.A1(n_1611),
.A2(n_1606),
.B1(n_1601),
.B2(n_1589),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1618),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1629),
.B(n_1606),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1623),
.Y(n_1663)
);

OA21x2_ASAP7_75t_L g1664 ( 
.A1(n_1634),
.A2(n_1574),
.B(n_1554),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1618),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1627),
.B(n_1599),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1649),
.B(n_1629),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1664),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1650),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1646),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1644),
.A2(n_1634),
.B1(n_1612),
.B2(n_1619),
.C(n_1640),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1651),
.Y(n_1672)
);

OAI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1664),
.A2(n_1611),
.B1(n_1599),
.B2(n_1601),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1663),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1664),
.A2(n_1601),
.B1(n_1589),
.B2(n_1606),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1649),
.B(n_1637),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1647),
.B(n_1637),
.C(n_1625),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1655),
.A2(n_1639),
.B1(n_1605),
.B2(n_1595),
.C(n_1613),
.Y(n_1678)
);

O2A1O1Ixp33_ASAP7_75t_SL g1679 ( 
.A1(n_1642),
.A2(n_1558),
.B(n_1551),
.C(n_1548),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1652),
.B(n_1639),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1648),
.B(n_1625),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1664),
.A2(n_1589),
.B1(n_1625),
.B2(n_1603),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1646),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1658),
.A2(n_1603),
.B(n_1495),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1642),
.B(n_1598),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1671),
.A2(n_1660),
.B1(n_1648),
.B2(n_1663),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1667),
.B(n_1676),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1672),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1685),
.B(n_1646),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1672),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1680),
.Y(n_1691)
);

NAND2x1p5_ASAP7_75t_L g1692 ( 
.A(n_1669),
.B(n_1643),
.Y(n_1692)
);

NAND2x1p5_ASAP7_75t_L g1693 ( 
.A(n_1674),
.B(n_1643),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1678),
.B(n_1652),
.Y(n_1694)
);

OAI21xp33_ASAP7_75t_L g1695 ( 
.A1(n_1681),
.A2(n_1647),
.B(n_1677),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1684),
.B(n_1656),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1670),
.B(n_1643),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1686),
.A2(n_1668),
.B(n_1673),
.Y(n_1698)
);

AOI211xp5_ASAP7_75t_L g1699 ( 
.A1(n_1695),
.A2(n_1679),
.B(n_1668),
.C(n_1683),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1697),
.A2(n_1675),
.B(n_1660),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1693),
.B(n_1645),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1694),
.A2(n_1651),
.B1(n_1659),
.B2(n_1662),
.C(n_1645),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1691),
.A2(n_1651),
.B1(n_1659),
.B2(n_1662),
.C(n_1645),
.Y(n_1703)
);

AOI222xp33_ASAP7_75t_L g1704 ( 
.A1(n_1690),
.A2(n_1657),
.B1(n_1666),
.B2(n_1659),
.C1(n_1661),
.C2(n_1665),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1696),
.B(n_1692),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1688),
.A2(n_1687),
.B(n_1689),
.Y(n_1706)
);

NAND4xp25_ASAP7_75t_L g1707 ( 
.A(n_1688),
.B(n_1682),
.C(n_1657),
.D(n_1663),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1699),
.B(n_1645),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1698),
.A2(n_1666),
.B1(n_1603),
.B2(n_1546),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1701),
.Y(n_1710)
);

NAND2xp33_ASAP7_75t_L g1711 ( 
.A(n_1703),
.B(n_1653),
.Y(n_1711)
);

OAI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1707),
.A2(n_1546),
.B1(n_1608),
.B2(n_1633),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_L g1713 ( 
.A(n_1711),
.B(n_1705),
.C(n_1706),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1710),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1708),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1712),
.Y(n_1716)
);

NOR2x1_ASAP7_75t_L g1717 ( 
.A(n_1709),
.B(n_1700),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1711),
.Y(n_1718)
);

AOI211xp5_ASAP7_75t_L g1719 ( 
.A1(n_1713),
.A2(n_1702),
.B(n_1654),
.C(n_1665),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1714),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1718),
.B(n_1704),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1715),
.B(n_1653),
.Y(n_1722)
);

XNOR2xp5_ASAP7_75t_L g1723 ( 
.A(n_1717),
.B(n_1603),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1722),
.Y(n_1724)
);

OAI31xp33_ASAP7_75t_L g1725 ( 
.A1(n_1721),
.A2(n_1716),
.A3(n_1661),
.B(n_1654),
.Y(n_1725)
);

NOR2xp67_ASAP7_75t_L g1726 ( 
.A(n_1723),
.B(n_1615),
.Y(n_1726)
);

NAND2x1_ASAP7_75t_L g1727 ( 
.A(n_1726),
.B(n_1720),
.Y(n_1727)
);

OAI211xp5_ASAP7_75t_SL g1728 ( 
.A1(n_1727),
.A2(n_1725),
.B(n_1724),
.C(n_1719),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1728),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1729),
.Y(n_1730)
);

OR5x1_ASAP7_75t_L g1731 ( 
.A(n_1730),
.B(n_1574),
.C(n_1608),
.D(n_1633),
.E(n_1577),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1731),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1731),
.A2(n_1632),
.B1(n_1636),
.B2(n_1628),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1732),
.A2(n_1632),
.B1(n_1622),
.B2(n_1621),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1733),
.A2(n_1620),
.B(n_1592),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1734),
.A2(n_1586),
.B(n_1591),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1735),
.A2(n_1592),
.B(n_1577),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_SL g1738 ( 
.A1(n_1736),
.A2(n_1597),
.B1(n_1595),
.B2(n_1605),
.Y(n_1738)
);

AOI322xp5_ASAP7_75t_L g1739 ( 
.A1(n_1737),
.A2(n_1577),
.A3(n_1586),
.B1(n_1592),
.B2(n_1591),
.C1(n_1546),
.C2(n_1585),
.Y(n_1739)
);

AOI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1738),
.A2(n_1586),
.B1(n_1591),
.B2(n_1585),
.Y(n_1740)
);

AOI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1740),
.A2(n_1739),
.B(n_1528),
.C(n_1585),
.Y(n_1741)
);


endmodule