module fake_netlist_1_7402_n_740 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_740);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_740;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g82 ( .A(n_10), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_21), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_74), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_33), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_64), .Y(n_86) );
INVxp33_ASAP7_75t_L g87 ( .A(n_71), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_47), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_63), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_51), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_13), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_50), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_48), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_15), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_61), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_45), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_8), .Y(n_97) );
INVx1_ASAP7_75t_SL g98 ( .A(n_6), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_32), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_37), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_72), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_23), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_31), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_19), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_57), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_4), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_46), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_76), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_10), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_1), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_8), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_38), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_73), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_41), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_66), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_9), .Y(n_117) );
INVxp33_ASAP7_75t_L g118 ( .A(n_62), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_28), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_34), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_54), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_2), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_18), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_4), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_5), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_79), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_26), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_25), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_36), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_30), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_2), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_114), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_114), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_114), .Y(n_134) );
NAND2x1_ASAP7_75t_L g135 ( .A(n_91), .B(n_0), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_105), .B(n_0), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_116), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_92), .B(n_1), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_83), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_83), .Y(n_141) );
NOR2xp67_ASAP7_75t_L g142 ( .A(n_122), .B(n_3), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_97), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_92), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_111), .B(n_3), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_95), .Y(n_146) );
INVxp67_ASAP7_75t_L g147 ( .A(n_107), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_94), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_125), .A2(n_131), .B1(n_94), .B2(n_119), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_110), .B(n_5), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_108), .B(n_6), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_88), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_108), .Y(n_154) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_88), .B(n_43), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_129), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_95), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_129), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_119), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_82), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_86), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_89), .B(n_7), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_86), .Y(n_163) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_89), .A2(n_44), .B(n_80), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_121), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_121), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_93), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_93), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_96), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_96), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_128), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_126), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_130), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_84), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_87), .B(n_7), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_139), .B(n_106), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_161), .B(n_103), .Y(n_178) );
OR2x6_ASAP7_75t_L g179 ( .A(n_148), .B(n_117), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_139), .Y(n_180) );
NAND2xp33_ASAP7_75t_L g181 ( .A(n_163), .B(n_127), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_161), .B(n_118), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_148), .B(n_127), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_132), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_132), .Y(n_186) );
BUFx4f_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_139), .Y(n_188) );
AND2x6_ASAP7_75t_L g189 ( .A(n_152), .B(n_104), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_132), .Y(n_190) );
NAND3xp33_ASAP7_75t_L g191 ( .A(n_176), .B(n_126), .C(n_123), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_132), .Y(n_194) );
AND2x6_ASAP7_75t_L g195 ( .A(n_176), .B(n_120), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_160), .B(n_98), .Y(n_196) );
BUFx4f_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_168), .B(n_102), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_168), .B(n_101), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_168), .B(n_109), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_147), .B(n_112), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_133), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_156), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_133), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_156), .Y(n_205) );
INVx4_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_156), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_167), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_153), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_170), .B(n_115), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_134), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_175), .B(n_113), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_138), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_153), .B(n_171), .Y(n_215) );
AND2x2_ASAP7_75t_SL g216 ( .A(n_136), .B(n_85), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_170), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_163), .B(n_117), .Y(n_218) );
AND2x6_ASAP7_75t_L g219 ( .A(n_172), .B(n_100), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_165), .B(n_99), .Y(n_220) );
INVx4_ASAP7_75t_SL g221 ( .A(n_167), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_172), .B(n_90), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_172), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_156), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_169), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_169), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_143), .B(n_42), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_144), .Y(n_228) );
INVx4_ASAP7_75t_L g229 ( .A(n_165), .Y(n_229) );
OR2x2_ASAP7_75t_L g230 ( .A(n_151), .B(n_9), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_166), .B(n_11), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_167), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_166), .B(n_11), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_144), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_156), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_173), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_154), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_154), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_173), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_174), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_174), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_137), .B(n_12), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_216), .B(n_137), .Y(n_243) );
OR2x6_ASAP7_75t_L g244 ( .A(n_179), .B(n_145), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_180), .A2(n_164), .B(n_162), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_206), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_190), .Y(n_247) );
AND2x6_ASAP7_75t_SL g248 ( .A(n_179), .B(n_145), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_216), .B(n_150), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_206), .B(n_174), .Y(n_250) );
NAND3xp33_ASAP7_75t_L g251 ( .A(n_188), .B(n_174), .C(n_167), .Y(n_251) );
NOR2xp67_ASAP7_75t_L g252 ( .A(n_229), .B(n_149), .Y(n_252) );
OR2x6_ASAP7_75t_L g253 ( .A(n_179), .B(n_135), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_190), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_188), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_217), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_183), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_236), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_229), .B(n_142), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_184), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_222), .B(n_174), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_187), .A2(n_167), .B1(n_158), .B2(n_164), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_222), .B(n_164), .Y(n_263) );
AO22x1_ASAP7_75t_L g264 ( .A1(n_236), .A2(n_157), .B1(n_141), .B2(n_159), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_187), .A2(n_158), .B1(n_159), .B2(n_157), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_223), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_202), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_188), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_222), .B(n_146), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_197), .A2(n_146), .B1(n_141), .B2(n_140), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_202), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_177), .B(n_140), .Y(n_272) );
INVxp67_ASAP7_75t_L g273 ( .A(n_239), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_201), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_207), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_178), .B(n_158), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_197), .A2(n_158), .B1(n_13), .B2(n_14), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_207), .Y(n_278) );
INVx4_ASAP7_75t_L g279 ( .A(n_189), .Y(n_279) );
NAND2x1p5_ASAP7_75t_L g280 ( .A(n_230), .B(n_158), .Y(n_280) );
NOR2xp67_ASAP7_75t_L g281 ( .A(n_191), .B(n_12), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_215), .B(n_53), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_185), .Y(n_283) );
NOR2x1_ASAP7_75t_L g284 ( .A(n_242), .B(n_14), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_204), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_185), .Y(n_286) );
AND2x4_ASAP7_75t_SL g287 ( .A(n_218), .B(n_15), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_212), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_182), .B(n_16), .Y(n_289) );
INVx5_ASAP7_75t_L g290 ( .A(n_189), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_228), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_198), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_234), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_182), .B(n_17), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_237), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_186), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_220), .B(n_20), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_198), .B(n_22), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_177), .B(n_24), .Y(n_299) );
OAI22xp33_ASAP7_75t_L g300 ( .A1(n_231), .A2(n_27), .B1(n_29), .B2(n_35), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_186), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_198), .B(n_39), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_196), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_225), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_SL g306 ( .A1(n_227), .A2(n_40), .B(n_49), .C(n_52), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_177), .B(n_55), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_192), .A2(n_56), .B1(n_58), .B2(n_59), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_193), .B(n_60), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_199), .B(n_65), .Y(n_310) );
NOR2x2_ASAP7_75t_L g311 ( .A(n_181), .B(n_67), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_226), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_199), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_244), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_279), .B(n_233), .Y(n_315) );
OAI21xp33_ASAP7_75t_L g316 ( .A1(n_274), .A2(n_181), .B(n_213), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_268), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_290), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_279), .B(n_199), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_290), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_290), .B(n_211), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_261), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_256), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_274), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_272), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_249), .B(n_195), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_266), .Y(n_327) );
INVx3_ASAP7_75t_SL g328 ( .A(n_244), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_290), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_302), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_292), .A2(n_211), .B1(n_210), .B2(n_214), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_291), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_261), .Y(n_333) );
AND2x6_ASAP7_75t_L g334 ( .A(n_310), .B(n_211), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_305), .Y(n_335) );
AOI21x1_ASAP7_75t_L g336 ( .A1(n_263), .A2(n_241), .B(n_240), .Y(n_336) );
AOI21x1_ASAP7_75t_L g337 ( .A1(n_263), .A2(n_194), .B(n_208), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_312), .Y(n_338) );
INVx5_ASAP7_75t_L g339 ( .A(n_254), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_313), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_304), .B(n_195), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_285), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_260), .B(n_195), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_254), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_273), .B(n_195), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_243), .B(n_195), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_254), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_293), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_269), .B(n_210), .Y(n_350) );
INVx6_ASAP7_75t_L g351 ( .A(n_272), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_295), .B(n_189), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_244), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_257), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_276), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_255), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_267), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_252), .B(n_189), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_255), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_253), .A2(n_189), .B1(n_200), .B2(n_219), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_275), .Y(n_361) );
OR2x6_ASAP7_75t_L g362 ( .A(n_253), .B(n_227), .Y(n_362) );
NOR2xp33_ASAP7_75t_SL g363 ( .A(n_258), .B(n_200), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_246), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_280), .B(n_200), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_278), .Y(n_366) );
INVx6_ASAP7_75t_L g367 ( .A(n_253), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_271), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_245), .A2(n_194), .B(n_235), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_319), .B(n_299), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_337), .A2(n_262), .B(n_310), .Y(n_371) );
OAI22xp33_ASAP7_75t_SL g372 ( .A1(n_324), .A2(n_308), .B1(n_311), .B2(n_277), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_336), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_369), .A2(n_282), .B(n_303), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_323), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_323), .Y(n_376) );
OAI21x1_ASAP7_75t_L g377 ( .A1(n_315), .A2(n_282), .B(n_298), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_339), .Y(n_378) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_355), .A2(n_309), .B(n_307), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_327), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_315), .A2(n_308), .B(n_280), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_327), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_352), .A2(n_284), .B(n_294), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g384 ( .A1(n_324), .A2(n_259), .B(n_289), .C(n_265), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_351), .A2(n_287), .B1(n_270), .B2(n_281), .Y(n_385) );
OA21x2_ASAP7_75t_L g386 ( .A1(n_326), .A2(n_297), .B(n_251), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_339), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_365), .A2(n_251), .B(n_250), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_SL g389 ( .A1(n_332), .A2(n_306), .B(n_300), .C(n_250), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_332), .Y(n_390) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_316), .A2(n_368), .B(n_349), .Y(n_391) );
OAI21x1_ASAP7_75t_L g392 ( .A1(n_368), .A2(n_235), .B(n_208), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_335), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_354), .A2(n_247), .B(n_296), .Y(n_394) );
AO31x2_ASAP7_75t_L g395 ( .A1(n_338), .A2(n_205), .A3(n_224), .B(n_283), .Y(n_395) );
AOI21x1_ASAP7_75t_L g396 ( .A1(n_357), .A2(n_224), .B(n_205), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_351), .A2(n_219), .B1(n_200), .B2(n_248), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_367), .A2(n_264), .B1(n_200), .B2(n_219), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_325), .Y(n_399) );
OAI222xp33_ASAP7_75t_L g400 ( .A1(n_362), .A2(n_232), .B1(n_209), .B2(n_219), .C1(n_301), .C2(n_286), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_342), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_367), .A2(n_219), .B1(n_183), .B2(n_257), .Y(n_402) );
OAI21x1_ASAP7_75t_L g403 ( .A1(n_329), .A2(n_232), .B(n_209), .Y(n_403) );
A2O1A1Ixp33_ASAP7_75t_L g404 ( .A1(n_350), .A2(n_183), .B(n_203), .C(n_257), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_372), .A2(n_353), .B1(n_314), .B2(n_348), .C(n_350), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_399), .A2(n_328), .B1(n_353), .B2(n_367), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_372), .A2(n_351), .B1(n_358), .B2(n_362), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_378), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_385), .A2(n_358), .B1(n_362), .B2(n_328), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_393), .B(n_341), .Y(n_411) );
AOI21xp33_ASAP7_75t_L g412 ( .A1(n_384), .A2(n_362), .B(n_346), .Y(n_412) );
CKINVDCx11_ASAP7_75t_R g413 ( .A(n_378), .Y(n_413) );
AND2x6_ASAP7_75t_L g414 ( .A(n_375), .B(n_319), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g415 ( .A1(n_375), .A2(n_343), .B1(n_363), .B2(n_360), .Y(n_415) );
AO21x1_ASAP7_75t_L g416 ( .A1(n_373), .A2(n_346), .B(n_331), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_376), .B(n_333), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_380), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_376), .A2(n_330), .B1(n_345), .B2(n_340), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_389), .A2(n_354), .B(n_321), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_382), .B(n_322), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g422 ( .A1(n_379), .A2(n_358), .B(n_330), .C(n_364), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_382), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_378), .B(n_339), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g425 ( .A1(n_397), .A2(n_317), .B(n_361), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_390), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_390), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_393), .B(n_319), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_401), .A2(n_334), .B1(n_359), .B2(n_356), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_401), .B(n_366), .Y(n_431) );
CKINVDCx11_ASAP7_75t_R g432 ( .A(n_387), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_398), .A2(n_334), .B1(n_321), .B2(n_357), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_387), .B(n_366), .Y(n_434) );
NOR2xp33_ASAP7_75t_SL g435 ( .A(n_414), .B(n_400), .Y(n_435) );
INVx4_ASAP7_75t_L g436 ( .A(n_414), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_405), .A2(n_334), .B1(n_381), .B2(n_370), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_423), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_417), .B(n_391), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_418), .Y(n_440) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_426), .B(n_373), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_408), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_417), .B(n_391), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_423), .Y(n_444) );
OAI211xp5_ASAP7_75t_L g445 ( .A1(n_407), .A2(n_402), .B(n_404), .C(n_381), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_418), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_414), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_421), .B(n_391), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_409), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_427), .B(n_395), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_427), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_409), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_428), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_414), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_408), .Y(n_455) );
INVx5_ASAP7_75t_L g456 ( .A(n_414), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_406), .B(n_413), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_428), .A2(n_370), .B1(n_386), .B2(n_339), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_421), .B(n_395), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_424), .B(n_370), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_412), .A2(n_334), .B1(n_383), .B2(n_386), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_434), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_424), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_426), .B(n_383), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_431), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_434), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_411), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_424), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_429), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_450), .Y(n_471) );
OAI21xp33_ASAP7_75t_L g472 ( .A1(n_435), .A2(n_410), .B(n_433), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_440), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_440), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_459), .B(n_416), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_450), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_462), .B(n_432), .Y(n_477) );
AOI211xp5_ASAP7_75t_L g478 ( .A1(n_457), .A2(n_419), .B(n_415), .C(n_416), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_459), .B(n_395), .Y(n_479) );
AO31x2_ASAP7_75t_L g480 ( .A1(n_458), .A2(n_422), .A3(n_420), .B(n_361), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_451), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_463), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_451), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_467), .B(n_395), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_453), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g486 ( .A(n_437), .B(n_430), .C(n_425), .D(n_394), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_467), .B(n_395), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_453), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_467), .B(n_414), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_449), .B(n_452), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_446), .Y(n_492) );
AOI211xp5_ASAP7_75t_L g493 ( .A1(n_435), .A2(n_403), .B(n_377), .C(n_392), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_449), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_464), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_449), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_452), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_462), .B(n_334), .Y(n_498) );
NOR3xp33_ASAP7_75t_SL g499 ( .A(n_445), .B(n_68), .C(n_70), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_452), .Y(n_500) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_461), .A2(n_386), .B1(n_318), .B2(n_344), .C(n_329), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_438), .B(n_386), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_438), .B(n_371), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_444), .B(n_371), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_442), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_466), .B(n_388), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g507 ( .A1(n_454), .A2(n_377), .B1(n_344), .B2(n_347), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_444), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_466), .B(n_388), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_439), .B(n_392), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_446), .Y(n_511) );
BUFx3_ASAP7_75t_L g512 ( .A(n_464), .Y(n_512) );
INVx1_ASAP7_75t_SL g513 ( .A(n_455), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_468), .B(n_347), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_436), .A2(n_374), .B1(n_347), .B2(n_329), .Y(n_515) );
OAI31xp33_ASAP7_75t_L g516 ( .A1(n_454), .A2(n_318), .A3(n_320), .B(n_221), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_448), .B(n_374), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_443), .B(n_403), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_446), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_448), .B(n_347), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_465), .B(n_396), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_468), .B(n_75), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_513), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_495), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_482), .B(n_470), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_481), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_481), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_477), .B(n_442), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_483), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_479), .B(n_465), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_483), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_508), .B(n_470), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_494), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_494), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_471), .B(n_476), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_485), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_479), .B(n_470), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_475), .B(n_465), .Y(n_538) );
INVx3_ASAP7_75t_L g539 ( .A(n_521), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_485), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_488), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_488), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_496), .Y(n_543) );
AND2x4_ASAP7_75t_SL g544 ( .A(n_489), .B(n_436), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_475), .B(n_465), .Y(n_545) );
OAI32xp33_ASAP7_75t_L g546 ( .A1(n_505), .A2(n_436), .A3(n_455), .B1(n_447), .B2(n_469), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_471), .B(n_468), .Y(n_547) );
INVx4_ASAP7_75t_SL g548 ( .A(n_495), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_476), .B(n_455), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_497), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_490), .B(n_464), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_490), .B(n_447), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_484), .B(n_447), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_484), .B(n_447), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_472), .B(n_436), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_496), .B(n_460), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_500), .Y(n_557) );
BUFx12f_ASAP7_75t_L g558 ( .A(n_512), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_517), .B(n_456), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_500), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_512), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_473), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_517), .B(n_502), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_489), .B(n_456), .Y(n_564) );
AND2x4_ASAP7_75t_SL g565 ( .A(n_487), .B(n_460), .Y(n_565) );
AND2x2_ASAP7_75t_SL g566 ( .A(n_521), .B(n_456), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_487), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_520), .B(n_456), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_473), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_502), .B(n_456), .Y(n_570) );
OAI21x1_ASAP7_75t_L g571 ( .A1(n_515), .A2(n_441), .B(n_458), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_472), .B(n_460), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_520), .B(n_460), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_474), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_503), .B(n_441), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_474), .B(n_492), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_491), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_491), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_498), .B(n_460), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_492), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_511), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_511), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_503), .B(n_456), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_563), .B(n_538), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_563), .B(n_506), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_537), .B(n_518), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_548), .B(n_493), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_526), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_527), .Y(n_589) );
NAND4xp25_ASAP7_75t_L g590 ( .A(n_555), .B(n_478), .C(n_493), .D(n_486), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_533), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_528), .B(n_509), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_567), .B(n_518), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_529), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_535), .B(n_478), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_525), .B(n_519), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_531), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_532), .B(n_510), .Y(n_598) );
INVxp67_ASAP7_75t_L g599 ( .A(n_523), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_574), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_536), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_550), .B(n_510), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_558), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_538), .B(n_521), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_533), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_540), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_541), .B(n_519), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_547), .B(n_504), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_542), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_545), .B(n_521), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_545), .B(n_553), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_554), .B(n_504), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_530), .B(n_480), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_534), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_557), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_530), .B(n_480), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_575), .B(n_480), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_575), .B(n_480), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_539), .B(n_480), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_534), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_543), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_543), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_539), .B(n_507), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_549), .B(n_514), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_539), .B(n_583), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_583), .B(n_522), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_560), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_560), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_559), .B(n_522), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_559), .B(n_499), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_574), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_569), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_561), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_562), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_558), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_559), .B(n_203), .Y(n_636) );
OAI31xp33_ASAP7_75t_L g637 ( .A1(n_555), .A2(n_501), .A3(n_516), .B(n_320), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_562), .Y(n_638) );
AOI21xp33_ASAP7_75t_SL g639 ( .A1(n_603), .A2(n_566), .B(n_524), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_606), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_606), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_609), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_609), .Y(n_643) );
AOI21xp33_ASAP7_75t_SL g644 ( .A1(n_603), .A2(n_566), .B(n_524), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_588), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_635), .A2(n_572), .B1(n_565), .B2(n_528), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_595), .B(n_572), .Y(n_647) );
NAND4xp25_ASAP7_75t_SL g648 ( .A(n_633), .B(n_570), .C(n_573), .D(n_551), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_590), .A2(n_556), .B1(n_552), .B2(n_579), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_592), .B(n_584), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_591), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_589), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_594), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_597), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_599), .A2(n_565), .B1(n_544), .B2(n_579), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_630), .A2(n_568), .B1(n_544), .B2(n_564), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_584), .B(n_548), .Y(n_657) );
AOI31xp33_ASAP7_75t_L g658 ( .A1(n_587), .A2(n_548), .A3(n_546), .B(n_582), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_601), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_615), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_625), .B(n_578), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_602), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_602), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_600), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_632), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_625), .B(n_577), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_632), .Y(n_667) );
O2A1O1Ixp5_ASAP7_75t_L g668 ( .A1(n_630), .A2(n_576), .B(n_580), .C(n_581), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_631), .B(n_581), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_585), .B(n_580), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_593), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_623), .A2(n_571), .B(n_203), .C(n_183), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_611), .B(n_571), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_604), .B(n_203), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_586), .B(n_77), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_631), .B(n_354), .C(n_81), .Y(n_676) );
NOR4xp25_ASAP7_75t_SL g677 ( .A(n_614), .B(n_78), .C(n_396), .D(n_221), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_647), .B(n_616), .Y(n_678) );
NOR2x1_ASAP7_75t_L g679 ( .A(n_658), .B(n_648), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_651), .Y(n_680) );
NOR2x1_ASAP7_75t_L g681 ( .A(n_676), .B(n_623), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_664), .Y(n_682) );
OAI21xp5_ASAP7_75t_SL g683 ( .A1(n_639), .A2(n_637), .B(n_616), .Y(n_683) );
INVxp67_ASAP7_75t_L g684 ( .A(n_647), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_661), .Y(n_685) );
NOR3xp33_ASAP7_75t_L g686 ( .A(n_649), .B(n_636), .C(n_624), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_650), .B(n_611), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_651), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_649), .A2(n_613), .B1(n_618), .B2(n_617), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_662), .B(n_663), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_669), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_669), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_666), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_644), .B(n_628), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g695 ( .A1(n_668), .A2(n_636), .B(n_610), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_657), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_640), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_675), .Y(n_698) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_674), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_673), .A2(n_613), .B1(n_618), .B2(n_617), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_671), .B(n_593), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_697), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_700), .B(n_673), .Y(n_703) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_679), .A2(n_656), .B(n_672), .C(n_646), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_683), .A2(n_668), .B(n_655), .C(n_610), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_684), .A2(n_659), .B1(n_653), .B2(n_654), .C(n_660), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_691), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_691), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_686), .A2(n_652), .B1(n_645), .B2(n_643), .C(n_641), .Y(n_709) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_692), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_689), .A2(n_642), .B1(n_670), .B2(n_665), .C(n_667), .Y(n_711) );
INVx1_ASAP7_75t_SL g712 ( .A(n_696), .Y(n_712) );
INVx1_ASAP7_75t_SL g713 ( .A(n_698), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_699), .A2(n_604), .B1(n_619), .B2(n_629), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_694), .A2(n_586), .B1(n_598), .B2(n_612), .Y(n_715) );
OAI211xp5_ASAP7_75t_L g716 ( .A1(n_681), .A2(n_619), .B(n_598), .C(n_612), .Y(n_716) );
AOI221x1_ASAP7_75t_L g717 ( .A1(n_705), .A2(n_692), .B1(n_682), .B2(n_695), .C(n_690), .Y(n_717) );
OAI211xp5_ASAP7_75t_SL g718 ( .A1(n_704), .A2(n_694), .B(n_678), .C(n_701), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_716), .A2(n_685), .B(n_693), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_703), .A2(n_687), .B1(n_680), .B2(n_688), .C(n_596), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_709), .A2(n_680), .B1(n_688), .B2(n_608), .C(n_607), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_707), .A2(n_614), .B(n_620), .C(n_621), .Y(n_722) );
AOI211xp5_ASAP7_75t_SL g723 ( .A1(n_715), .A2(n_608), .B(n_629), .C(n_626), .Y(n_723) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_711), .A2(n_622), .B1(n_628), .B2(n_591), .C(n_605), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g725 ( .A(n_707), .B(n_677), .C(n_627), .Y(n_725) );
AND2x4_ASAP7_75t_L g726 ( .A(n_719), .B(n_713), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_718), .B(n_712), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_722), .B(n_710), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_721), .B(n_702), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_723), .B(n_714), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_727), .B(n_717), .C(n_725), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_726), .A2(n_720), .B1(n_708), .B2(n_724), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_730), .B(n_706), .Y(n_733) );
OAI21xp5_ASAP7_75t_L g734 ( .A1(n_731), .A2(n_729), .B(n_728), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_733), .B(n_605), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_735), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_736), .Y(n_737) );
AOI222xp33_ASAP7_75t_L g738 ( .A1(n_737), .A2(n_734), .B1(n_732), .B2(n_627), .C1(n_634), .C2(n_638), .Y(n_738) );
OA22x2_ASAP7_75t_L g739 ( .A1(n_738), .A2(n_634), .B1(n_638), .B2(n_626), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_739), .A2(n_354), .B(n_221), .Y(n_740) );
endmodule