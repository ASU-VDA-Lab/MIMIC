module fake_jpeg_29565_n_500 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_500);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_500;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_15),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_56),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g140 ( 
.A(n_53),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_65),
.Y(n_112)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_88),
.Y(n_121)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_67),
.Y(n_133)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_72),
.Y(n_136)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_78),
.Y(n_119)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_49),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_30),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_8),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_9),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_50),
.Y(n_126)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_91),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_93),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_40),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_97),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_39),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_98),
.Y(n_129)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_45),
.B1(n_37),
.B2(n_44),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_101),
.A2(n_145),
.B1(n_149),
.B2(n_27),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_66),
.B(n_50),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_41),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_37),
.B1(n_36),
.B2(n_44),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_107),
.A2(n_110),
.B1(n_111),
.B2(n_47),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_56),
.A2(n_37),
.B1(n_48),
.B2(n_27),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_126),
.B(n_130),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_59),
.B(n_46),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_45),
.C(n_33),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_72),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_82),
.B(n_43),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_137),
.B(n_39),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_54),
.A2(n_32),
.B1(n_43),
.B2(n_42),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_32),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_31),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_70),
.A2(n_31),
.B1(n_42),
.B2(n_41),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_60),
.A2(n_13),
.B(n_14),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_39),
.B(n_29),
.Y(n_175)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_156),
.Y(n_240)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_47),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_174),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_159),
.B(n_162),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_160),
.B(n_167),
.Y(n_229)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_176),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_110),
.A2(n_124),
.B1(n_118),
.B2(n_141),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_164),
.A2(n_186),
.B1(n_136),
.B2(n_103),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_165),
.Y(n_214)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_166),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g167 ( 
.A(n_105),
.B(n_77),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_105),
.A2(n_81),
.B1(n_87),
.B2(n_96),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_SL g247 ( 
.A1(n_168),
.A2(n_192),
.B(n_201),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_169),
.A2(n_202),
.B(n_195),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_170),
.A2(n_197),
.B1(n_203),
.B2(n_205),
.Y(n_239)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

OR2x2_ASAP7_75t_SL g174 ( 
.A(n_110),
.B(n_55),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_181),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_98),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_177),
.B(n_178),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_98),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_23),
.C(n_90),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_195),
.C(n_206),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_129),
.B(n_99),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_180),
.B(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_23),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_80),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_84),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_183),
.B(n_193),
.Y(n_245)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_123),
.A2(n_79),
.B1(n_58),
.B2(n_61),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_100),
.Y(n_189)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_191),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_140),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_116),
.A2(n_64),
.B1(n_83),
.B2(n_74),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_140),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_101),
.A2(n_39),
.B1(n_76),
.B2(n_91),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_194),
.A2(n_139),
.B1(n_122),
.B2(n_123),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_120),
.B(n_29),
.Y(n_195)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_115),
.B1(n_116),
.B2(n_109),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_125),
.A2(n_69),
.B1(n_11),
.B2(n_12),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_139),
.B1(n_122),
.B2(n_133),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_132),
.B(n_63),
.Y(n_202)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_242)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_125),
.B(n_150),
.Y(n_206)
);

OAI22x1_ASAP7_75t_SL g207 ( 
.A1(n_174),
.A2(n_107),
.B1(n_109),
.B2(n_102),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g267 ( 
.A1(n_207),
.A2(n_186),
.B(n_204),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_208),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_220),
.A2(n_230),
.B1(n_237),
.B2(n_199),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_115),
.B1(n_148),
.B2(n_132),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_160),
.A2(n_131),
.B1(n_109),
.B2(n_147),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_222),
.A2(n_244),
.B1(n_158),
.B2(n_199),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_170),
.A2(n_131),
.B1(n_103),
.B2(n_133),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_226),
.A2(n_197),
.B1(n_203),
.B2(n_166),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_151),
.B1(n_144),
.B2(n_136),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_179),
.B(n_151),
.C(n_144),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_246),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_63),
.B1(n_53),
.B2(n_29),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_163),
.B1(n_198),
.B2(n_184),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_169),
.A2(n_53),
.B1(n_29),
.B2(n_2),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_242),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_169),
.A2(n_7),
.B1(n_13),
.B2(n_11),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_175),
.B(n_196),
.C(n_201),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_162),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_248),
.A2(n_6),
.B1(n_10),
.B2(n_15),
.Y(n_279)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_249),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_207),
.A2(n_193),
.B1(n_161),
.B2(n_185),
.Y(n_250)
);

OAI22x1_ASAP7_75t_L g316 ( 
.A1(n_250),
.A2(n_266),
.B1(n_241),
.B2(n_216),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_172),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_252),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_209),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_171),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_253),
.B(n_256),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_167),
.B(n_200),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_254),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_255),
.A2(n_257),
.B1(n_271),
.B2(n_285),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_157),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_210),
.A2(n_158),
.B(n_198),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_261),
.A2(n_269),
.B(n_242),
.C(n_234),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_210),
.B(n_212),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_262),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_213),
.B(n_177),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_264),
.B(n_273),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_165),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_270),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_214),
.A2(n_228),
.B1(n_235),
.B2(n_216),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_267),
.A2(n_239),
.B1(n_236),
.B2(n_228),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_268),
.A2(n_279),
.B1(n_283),
.B2(n_241),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_210),
.A2(n_190),
.B(n_205),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_156),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_245),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_272),
.B(n_274),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_173),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_229),
.B(n_0),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_212),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_275),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_212),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_277),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_3),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_278),
.B(n_281),
.Y(n_322)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_3),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_224),
.A2(n_239),
.B1(n_225),
.B2(n_226),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_217),
.B(n_3),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_248),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_239),
.A2(n_204),
.B1(n_187),
.B2(n_4),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_211),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_252),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_294),
.C(n_295),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_237),
.C(n_215),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_233),
.C(n_234),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_296),
.A2(n_298),
.B1(n_308),
.B2(n_285),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_310),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_239),
.B1(n_244),
.B2(n_221),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_260),
.A2(n_208),
.B1(n_235),
.B2(n_233),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_305),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_273),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_311),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_314),
.A2(n_262),
.B(n_278),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_316),
.A2(n_243),
.B1(n_218),
.B2(n_10),
.Y(n_342)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_253),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_320),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_249),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_318),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_249),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_319),
.Y(n_345)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_255),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_284),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_321),
.Y(n_350)
);

OAI21xp33_ASAP7_75t_L g325 ( 
.A1(n_302),
.A2(n_272),
.B(n_274),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_325),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_326),
.A2(n_328),
.B1(n_351),
.B2(n_352),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_276),
.B1(n_254),
.B2(n_259),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_327),
.B(n_329),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_308),
.A2(n_257),
.B1(n_277),
.B2(n_275),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_300),
.A2(n_283),
.B1(n_268),
.B2(n_259),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_330),
.A2(n_347),
.B(n_306),
.Y(n_358)
);

XOR2x1_ASAP7_75t_SL g331 ( 
.A(n_314),
.B(n_261),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_331),
.B(n_330),
.Y(n_368)
);

A2O1A1O1Ixp25_ASAP7_75t_L g332 ( 
.A1(n_293),
.A2(n_269),
.B(n_256),
.C(n_265),
.D(n_281),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_332),
.B(n_294),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_291),
.A2(n_267),
.B1(n_266),
.B2(n_264),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_335),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_320),
.A2(n_267),
.B1(n_279),
.B2(n_270),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_291),
.B(n_267),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_336),
.B(n_289),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_288),
.B(n_223),
.C(n_219),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_346),
.C(n_349),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_317),
.A2(n_204),
.B1(n_218),
.B2(n_223),
.Y(n_340)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_243),
.B(n_6),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_341),
.A2(n_312),
.B(n_299),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_342),
.A2(n_355),
.B1(n_319),
.B2(n_318),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_287),
.B(n_218),
.C(n_4),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_309),
.A2(n_6),
.B(n_15),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_6),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_298),
.A2(n_4),
.B1(n_311),
.B2(n_313),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_313),
.A2(n_4),
.B1(n_309),
.B2(n_292),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_290),
.Y(n_354)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_354),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_321),
.A2(n_306),
.B1(n_303),
.B2(n_315),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_293),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_374),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_357),
.B(n_368),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_358),
.A2(n_380),
.B1(n_350),
.B2(n_353),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_324),
.B(n_295),
.C(n_315),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_362),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_322),
.C(n_289),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_333),
.Y(n_364)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_322),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_375),
.Y(n_391)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_338),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_373),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_370),
.A2(n_327),
.B1(n_329),
.B2(n_338),
.Y(n_404)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_301),
.C(n_304),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_331),
.C(n_346),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_301),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_305),
.C(n_299),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_352),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_290),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_328),
.Y(n_400)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_343),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_345),
.Y(n_396)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_383),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_336),
.A2(n_312),
.B(n_310),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_384),
.Y(n_388)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_351),
.Y(n_385)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_385),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_384),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_387),
.B(n_393),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_356),
.B(n_350),
.Y(n_393)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_396),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_360),
.B(n_339),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_398),
.B(n_407),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_402),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_334),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_404),
.A2(n_326),
.B1(n_378),
.B2(n_371),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_362),
.B(n_323),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_408),
.C(n_359),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_374),
.B(n_323),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_409),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_363),
.B(n_339),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_411),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_363),
.B(n_345),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_401),
.A2(n_377),
.B1(n_385),
.B2(n_379),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_414),
.A2(n_371),
.B1(n_365),
.B2(n_342),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_431),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_382),
.Y(n_418)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_418),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_396),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_422),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_359),
.C(n_376),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_421),
.B(n_429),
.C(n_406),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_388),
.A2(n_378),
.B(n_380),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_375),
.Y(n_424)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_424),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_411),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_428),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_361),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_427),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_395),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_386),
.B(n_373),
.C(n_368),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_377),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_388),
.B(n_361),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_SL g432 ( 
.A(n_405),
.B(n_402),
.C(n_358),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_432),
.B(n_400),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_443),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_435),
.B(n_447),
.Y(n_453)
);

AO21x1_ASAP7_75t_L g451 ( 
.A1(n_439),
.A2(n_432),
.B(n_416),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_394),
.C(n_408),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_441),
.B(n_442),
.C(n_444),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_405),
.C(n_407),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_391),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_391),
.C(n_401),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_404),
.C(n_366),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_446),
.B(n_365),
.C(n_424),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_403),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_430),
.Y(n_452)
);

NAND4xp25_ASAP7_75t_SL g449 ( 
.A(n_414),
.B(n_422),
.C(n_418),
.D(n_413),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_449),
.B(n_415),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_412),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_450),
.A2(n_458),
.B(n_341),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_451),
.B(n_452),
.Y(n_477)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_436),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_456),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_440),
.B(n_428),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_449),
.A2(n_413),
.B(n_431),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_459),
.B(n_464),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_433),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_462),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_461),
.B(n_427),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_415),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_392),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_463),
.A2(n_425),
.B1(n_445),
.B2(n_409),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_435),
.A2(n_412),
.B(n_425),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_SL g467 ( 
.A(n_451),
.B(n_457),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_467),
.B(n_474),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_468),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_444),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_469),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_475),
.Y(n_480)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_471),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_453),
.A2(n_442),
.B(n_446),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_472),
.A2(n_476),
.B(n_450),
.Y(n_485)
);

FAx1_ASAP7_75t_SL g474 ( 
.A(n_459),
.B(n_434),
.CI(n_443),
.CON(n_474),
.SN(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_458),
.A2(n_390),
.B1(n_389),
.B2(n_348),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_454),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_457),
.C(n_455),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_474),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_473),
.B(n_348),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_485),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_477),
.A2(n_340),
.B1(n_347),
.B2(n_471),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_486),
.B(n_468),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_481),
.B(n_466),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_488),
.B(n_490),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_489),
.Y(n_493)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_478),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_483),
.A2(n_465),
.B1(n_476),
.B2(n_466),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_491),
.A2(n_492),
.B(n_478),
.Y(n_494)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_494),
.Y(n_497)
);

AOI21x1_ASAP7_75t_L g496 ( 
.A1(n_495),
.A2(n_487),
.B(n_480),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_496),
.B(n_479),
.C(n_493),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_498),
.B(n_497),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_482),
.Y(n_500)
);


endmodule