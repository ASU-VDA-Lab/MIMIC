module fake_jpeg_3670_n_222 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_222);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_3),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_32),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_85),
.Y(n_88)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_65),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_61),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_62),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_64),
.B1(n_68),
.B2(n_58),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_68),
.B1(n_54),
.B2(n_78),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_78),
.B1(n_69),
.B2(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_55),
.B1(n_61),
.B2(n_69),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_79),
.B1(n_73),
.B2(n_60),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_0),
.Y(n_139)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_97),
.B(n_91),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_87),
.Y(n_121)
);

BUFx2_ASAP7_75t_SL g112 ( 
.A(n_96),
.Y(n_112)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_26),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_63),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_139),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_135),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_133),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_116),
.C(n_114),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_24),
.C(n_50),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_86),
.B1(n_71),
.B2(n_75),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_132),
.B1(n_60),
.B2(n_70),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_86),
.B1(n_71),
.B2(n_75),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_115),
.B(n_107),
.C(n_73),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_136),
.B(n_73),
.Y(n_148)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_27),
.B1(n_45),
.B2(n_44),
.Y(n_163)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

BUFx2_ASAP7_75t_SL g141 ( 
.A(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_1),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_1),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_9),
.B(n_10),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_149),
.A2(n_150),
.B1(n_7),
.B2(n_8),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_60),
.B1(n_66),
.B2(n_5),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_163),
.B1(n_131),
.B2(n_8),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_161),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_4),
.B(n_6),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_150),
.B(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_22),
.C(n_48),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_6),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_177),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_160),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_175),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_180),
.B1(n_13),
.B2(n_14),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_181),
.Y(n_188)
);

AOI22x1_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_20),
.B1(n_42),
.B2(n_40),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_183),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_175),
.B(n_169),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_186),
.B(n_189),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_29),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_30),
.C(n_38),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_180),
.C(n_170),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_192)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_199),
.C(n_203),
.Y(n_208)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

NOR2x1_ASAP7_75t_R g201 ( 
.A(n_193),
.B(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_194),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_202),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_187),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_173),
.C(n_174),
.Y(n_204)
);

XNOR2x1_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_176),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_193),
.B1(n_191),
.B2(n_195),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_184),
.B1(n_164),
.B2(n_166),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_196),
.B(n_197),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_207),
.B(n_200),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_212),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_214),
.Y(n_216)
);

NOR3xp33_ASAP7_75t_SL g214 ( 
.A(n_209),
.B(n_15),
.C(n_16),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_208),
.C(n_210),
.Y(n_217)
);

OAI21x1_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_216),
.B(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_53),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_18),
.C(n_35),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_36),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_17),
.Y(n_222)
);


endmodule