module fake_jpeg_8116_n_186 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_31),
.Y(n_35)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_43),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_21),
.B1(n_15),
.B2(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_21),
.B1(n_15),
.B2(n_16),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_34),
.B1(n_17),
.B2(n_13),
.Y(n_75)
);

BUFx12f_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_25),
.B1(n_17),
.B2(n_12),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_21),
.B1(n_33),
.B2(n_24),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_43),
.B1(n_34),
.B2(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_21),
.B(n_25),
.C(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_61),
.Y(n_66)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_14),
.B(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_57),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_22),
.B1(n_13),
.B2(n_17),
.Y(n_81)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_0),
.Y(n_73)
);

A2O1A1O1Ixp25_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_11),
.B(n_1),
.C(n_2),
.D(n_4),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_75),
.B1(n_51),
.B2(n_34),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_54),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_79),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_22),
.B(n_13),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_49),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_52),
.B1(n_59),
.B2(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_91),
.Y(n_100)
);

XNOR2x2_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_11),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_53),
.C(n_41),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_63),
.C(n_67),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_94),
.C(n_95),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_65),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_65),
.C(n_63),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_80),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_70),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_91),
.C(n_79),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_107),
.B1(n_22),
.B2(n_20),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_70),
.B(n_76),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_99),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_112),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_87),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_119),
.C(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_88),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_101),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_106),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_53),
.B1(n_37),
.B2(n_44),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_96),
.B1(n_93),
.B2(n_104),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_18),
.B(n_19),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_132),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_120),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_121),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_44),
.Y(n_146)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_111),
.C(n_109),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_136),
.C(n_26),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_96),
.B1(n_119),
.B2(n_95),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_144),
.B1(n_133),
.B2(n_123),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_110),
.B1(n_114),
.B2(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_147),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_130),
.A2(n_118),
.B(n_20),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_145),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_41),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_148),
.C(n_126),
.Y(n_151)
);

AOI21x1_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_44),
.B(n_19),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_14),
.B(n_1),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_153),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_155),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_125),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_149),
.B(n_158),
.Y(n_159)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_148),
.B(n_143),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_161),
.A2(n_0),
.B(n_4),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_125),
.B1(n_77),
.B2(n_36),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_18),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_77),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_165),
.C(n_164),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_169),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_168),
.A2(n_0),
.B(n_4),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_19),
.B1(n_36),
.B2(n_18),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_162),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_173),
.B(n_18),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_36),
.Y(n_173)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_26),
.C(n_18),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_177),
.A3(n_170),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_5),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_37),
.C2(n_30),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_178),
.C(n_37),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.C(n_5),
.Y(n_184)
);

OAI221xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_180),
.B1(n_8),
.B2(n_9),
.C(n_5),
.Y(n_185)
);

XNOR2x2_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_28),
.Y(n_186)
);


endmodule