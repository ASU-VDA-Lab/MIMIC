module fake_jpeg_21245_n_254 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_32),
.B1(n_25),
.B2(n_26),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_52),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_32),
.B1(n_29),
.B2(n_30),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_25),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_15),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_48),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_32),
.B1(n_25),
.B2(n_26),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_11),
.B1(n_15),
.B2(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_24),
.B1(n_31),
.B2(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_60),
.Y(n_87)
);

AO21x2_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_33),
.B(n_24),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_54),
.B1(n_31),
.B2(n_27),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_47),
.B1(n_24),
.B2(n_46),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_66),
.B1(n_27),
.B2(n_31),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_33),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_33),
.B(n_28),
.C(n_31),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_52),
.B(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_28),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_33),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_82),
.B1(n_83),
.B2(n_86),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_95),
.B(n_71),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_71),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_45),
.B1(n_48),
.B2(n_30),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_58),
.B1(n_29),
.B2(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_88),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_31),
.B1(n_27),
.B2(n_49),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_27),
.B1(n_53),
.B2(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_61),
.A2(n_53),
.B1(n_11),
.B2(n_15),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_80),
.B1(n_69),
.B2(n_79),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_14),
.B1(n_28),
.B2(n_22),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_61),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_17),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_65),
.B(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_96),
.B(n_106),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_111),
.B1(n_90),
.B2(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_63),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_95),
.B(n_63),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_71),
.B1(n_64),
.B2(n_67),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_75),
.B(n_69),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_33),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_84),
.B(n_81),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_21),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_84),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_128),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_121),
.B1(n_142),
.B2(n_103),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_71),
.B1(n_64),
.B2(n_76),
.Y(n_121)
);

OAI22x1_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_73),
.B1(n_57),
.B2(n_76),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_124),
.B1(n_127),
.B2(n_135),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_107),
.B1(n_100),
.B2(n_110),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_14),
.B1(n_73),
.B2(n_28),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_57),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_14),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_136),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_137),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_14),
.B1(n_22),
.B2(n_23),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_17),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_97),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_96),
.B1(n_99),
.B2(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_16),
.B1(n_23),
.B2(n_21),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_17),
.C(n_33),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_33),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_12),
.B1(n_23),
.B2(n_21),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_33),
.C(n_19),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_98),
.C(n_33),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_103),
.B1(n_105),
.B2(n_104),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_109),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_143),
.C(n_136),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_106),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_98),
.B1(n_97),
.B2(n_2),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_162),
.B1(n_121),
.B2(n_142),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_20),
.B1(n_16),
.B2(n_12),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_17),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_164),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_16),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_130),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_167),
.B(n_13),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_131),
.B(n_120),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g193 ( 
.A(n_169),
.B(n_146),
.Y(n_193)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_174),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_127),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_164),
.B(n_153),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_182),
.B1(n_152),
.B2(n_156),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_162),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_183),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_141),
.C(n_137),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_180),
.C(n_166),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_19),
.C(n_13),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_9),
.B1(n_10),
.B2(n_8),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_152),
.B1(n_144),
.B2(n_150),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_195),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_13),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_197),
.B(n_201),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_177),
.B1(n_169),
.B2(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_159),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_196),
.A2(n_181),
.B(n_171),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_167),
.C(n_160),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_166),
.C(n_19),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_19),
.C(n_13),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_8),
.B(n_10),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_168),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_213),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_168),
.C(n_181),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_199),
.C(n_198),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_197),
.A2(n_12),
.B(n_20),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_211),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_187),
.A2(n_20),
.B(n_8),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_6),
.B(n_10),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_201),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_217),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_186),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_223),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_206),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_SL g233 ( 
.A1(n_222),
.A2(n_214),
.B(n_6),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_200),
.C(n_19),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_213),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_224),
.B(n_203),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_225),
.B(n_232),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_R g227 ( 
.A(n_218),
.B(n_204),
.Y(n_227)
);

AOI21x1_ASAP7_75t_SL g237 ( 
.A1(n_227),
.A2(n_233),
.B(n_5),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_204),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_231),
.Y(n_239)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_223),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_207),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_6),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_238),
.B(n_10),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_5),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_241),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_1),
.B(n_3),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_5),
.B(n_7),
.C(n_9),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_5),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_7),
.C(n_9),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_245),
.B(n_1),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_240),
.A2(n_236),
.B(n_241),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_247),
.B(n_246),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_1),
.B(n_3),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_250),
.B(n_3),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_3),
.B(n_4),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_4),
.B(n_238),
.Y(n_254)
);


endmodule