module fake_jpeg_30572_n_86 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_34),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_51),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_35),
.B1(n_30),
.B2(n_29),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_61),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_31),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_60),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_3),
.Y(n_60)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_18),
.B(n_5),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_10),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_53),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_46),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_71),
.C(n_12),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_3),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_74),
.Y(n_78)
);

NOR4xp25_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_63),
.C(n_68),
.D(n_65),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_75),
.B1(n_73),
.B2(n_78),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_67),
.B1(n_74),
.B2(n_17),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_27),
.B(n_15),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_13),
.C(n_19),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_20),
.C(n_22),
.Y(n_84)
);

NAND2xp67_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_23),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_24),
.Y(n_86)
);


endmodule