module fake_jpeg_10606_n_116 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_116);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_20),
.Y(n_30)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_11),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_11),
.B1(n_10),
.B2(n_14),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_36),
.B1(n_14),
.B2(n_17),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_14),
.B1(n_17),
.B2(n_20),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_37),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_34),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_26),
.B1(n_24),
.B2(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_50),
.B1(n_61),
.B2(n_53),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_30),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_46),
.B(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_47),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_70),
.B1(n_44),
.B2(n_13),
.Y(n_80)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_67),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_21),
.B(n_36),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_42),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_41),
.B1(n_40),
.B2(n_43),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_41),
.B1(n_26),
.B2(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_72),
.Y(n_77)
);

A2O1A1O1Ixp25_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_60),
.B(n_45),
.C(n_48),
.D(n_51),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_12),
.B(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_62),
.C(n_66),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_12),
.B1(n_18),
.B2(n_2),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_18),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_90),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_74),
.C(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_76),
.C(n_82),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_0),
.B(n_1),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_18),
.C(n_9),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_97),
.C(n_90),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_8),
.C(n_1),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_100),
.C(n_98),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_87),
.B(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_87),
.B1(n_85),
.B2(n_2),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

NAND4xp25_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_92),
.C(n_3),
.D(n_4),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_107),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_0),
.C(n_3),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_5),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_5),
.B(n_109),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_112),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_108),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g115 ( 
.A(n_114),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_5),
.Y(n_116)
);


endmodule