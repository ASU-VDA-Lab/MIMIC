module fake_jpeg_11309_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_23),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_11),
.B1(n_15),
.B2(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_17),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_22),
.B1(n_19),
.B2(n_15),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_35),
.B1(n_24),
.B2(n_26),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_34),
.C(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_33),
.B1(n_35),
.B2(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_2),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_30),
.C(n_27),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_40),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_25),
.C(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_12),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_35),
.B(n_25),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_12),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_50),
.B(n_3),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_3),
.B(n_14),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_45),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_53),
.B1(n_49),
.B2(n_14),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_13),
.C(n_20),
.Y(n_55)
);


endmodule