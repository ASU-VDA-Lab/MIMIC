module fake_jpeg_11965_n_560 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_560);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_560;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_2),
.B(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_60),
.A2(n_59),
.B1(n_58),
.B2(n_52),
.Y(n_179)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_62),
.Y(n_182)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_63),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_64),
.B(n_81),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g186 ( 
.A(n_65),
.Y(n_186)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_66),
.Y(n_184)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_69),
.Y(n_197)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_73),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_75),
.B(n_97),
.Y(n_157)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_77),
.Y(n_181)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_20),
.B(n_3),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_83),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_19),
.B(n_16),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_88),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_25),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_4),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_102),
.Y(n_138)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_94),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_23),
.B(n_35),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_98),
.Y(n_174)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

NAND2x1_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_4),
.Y(n_100)
);

HAxp5_ASAP7_75t_SL g137 ( 
.A(n_100),
.B(n_65),
.CON(n_137),
.SN(n_137)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_25),
.Y(n_102)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_25),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_108),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_29),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_23),
.B(n_5),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_27),
.B(n_5),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_27),
.B(n_38),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_115),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

BUFx4f_ASAP7_75t_SL g115 ( 
.A(n_29),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_20),
.Y(n_116)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx11_ASAP7_75t_SL g117 ( 
.A(n_29),
.Y(n_117)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_21),
.Y(n_160)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_36),
.Y(n_121)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_28),
.B(n_38),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_122),
.B(n_35),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_61),
.A2(n_46),
.B1(n_56),
.B2(n_57),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_128),
.A2(n_130),
.B1(n_149),
.B2(n_151),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_63),
.A2(n_56),
.B1(n_57),
.B2(n_41),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_137),
.A2(n_163),
.B(n_200),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_89),
.A2(n_57),
.B1(n_41),
.B2(n_24),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_140),
.A2(n_180),
.B1(n_189),
.B2(n_193),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_64),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_142),
.B(n_166),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_77),
.A2(n_41),
.B1(n_24),
.B2(n_40),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_105),
.A2(n_24),
.B1(n_48),
.B2(n_40),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_199),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_160),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_80),
.A2(n_48),
.B1(n_40),
.B2(n_100),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_162),
.B(n_163),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_68),
.B(n_55),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_106),
.A2(n_48),
.B1(n_55),
.B2(n_21),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_164),
.A2(n_165),
.B1(n_185),
.B2(n_188),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_114),
.A2(n_55),
.B1(n_21),
.B2(n_53),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_60),
.B(n_54),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_103),
.A2(n_54),
.B(n_53),
.C(n_51),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_171),
.B(n_82),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_179),
.A2(n_187),
.B1(n_117),
.B2(n_73),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_79),
.A2(n_121),
.B1(n_123),
.B2(n_74),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_62),
.A2(n_21),
.B1(n_55),
.B2(n_51),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_84),
.A2(n_58),
.B1(n_52),
.B2(n_45),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_62),
.A2(n_59),
.B1(n_45),
.B2(n_28),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_86),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_94),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_95),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_194),
.A2(n_193),
.B1(n_140),
.B2(n_166),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_115),
.B(n_10),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_66),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_115),
.B(n_11),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_69),
.B(n_29),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_202),
.B(n_203),
.Y(n_272)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_204),
.Y(n_285)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_206),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_87),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_208),
.B(n_213),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_184),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_209),
.B(n_244),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_135),
.B(n_12),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_211),
.B(n_182),
.Y(n_273)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_212),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_158),
.B(n_71),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_214),
.B(n_223),
.Y(n_296)
);

BUFx12_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_215),
.Y(n_310)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_216),
.Y(n_319)
);

OR2x2_ASAP7_75t_SL g218 ( 
.A(n_137),
.B(n_116),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_218),
.A2(n_259),
.B(n_213),
.Y(n_313)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_220),
.B(n_267),
.Y(n_276)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_222),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_147),
.B(n_82),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_125),
.Y(n_224)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_133),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_225),
.B(n_236),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_127),
.B(n_101),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_226),
.B(n_227),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_146),
.B(n_72),
.Y(n_227)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_187),
.A2(n_112),
.B1(n_104),
.B2(n_78),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g320 ( 
.A1(n_229),
.A2(n_247),
.B1(n_264),
.B2(n_202),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_230),
.A2(n_237),
.B1(n_258),
.B2(n_256),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_124),
.B(n_120),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_231),
.B(n_232),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_158),
.B(n_66),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_125),
.Y(n_233)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_233),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_126),
.B(n_120),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_234),
.Y(n_295)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_144),
.Y(n_235)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_235),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_158),
.B(n_13),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_154),
.B(n_13),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_238),
.Y(n_308)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_239),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_142),
.B(n_13),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_245),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_242),
.A2(n_143),
.B1(n_156),
.B2(n_152),
.Y(n_293)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_135),
.B(n_14),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_246),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_179),
.A2(n_16),
.B1(n_98),
.B2(n_176),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_184),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_262),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_155),
.B(n_98),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_253),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_148),
.A2(n_169),
.B1(n_144),
.B2(n_176),
.Y(n_250)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_150),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_178),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_135),
.B(n_138),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_256),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_150),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_255),
.A2(n_260),
.B1(n_266),
.B2(n_268),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_168),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_181),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_258),
.B(n_261),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_163),
.B(n_169),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_173),
.C(n_183),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_148),
.A2(n_172),
.B1(n_167),
.B2(n_161),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_190),
.B(n_170),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g262 ( 
.A(n_192),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_195),
.A2(n_171),
.B1(n_145),
.B2(n_175),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_183),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_265),
.B(n_270),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_200),
.A2(n_143),
.B1(n_181),
.B2(n_141),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_129),
.B(n_132),
.Y(n_267)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_194),
.A2(n_162),
.B1(n_175),
.B2(n_145),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_129),
.B(n_132),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_173),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_271),
.B(n_205),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_273),
.B(n_318),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_218),
.B(n_197),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_275),
.B(n_305),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_313),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_217),
.A2(n_156),
.B1(n_134),
.B2(n_152),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_286),
.A2(n_302),
.B1(n_303),
.B2(n_327),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_210),
.B(n_134),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_304),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_293),
.A2(n_252),
.B1(n_243),
.B2(n_246),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_220),
.A2(n_136),
.B1(n_141),
.B2(n_182),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_297),
.A2(n_320),
.B1(n_321),
.B2(n_248),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_242),
.A2(n_136),
.B1(n_139),
.B2(n_217),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_263),
.A2(n_139),
.B1(n_268),
.B2(n_210),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_211),
.B(n_257),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_225),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_254),
.A2(n_257),
.B(n_240),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_306),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_270),
.B(n_259),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_315),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_230),
.B(n_268),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_245),
.B(n_241),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_268),
.B(n_204),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_324),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_222),
.B(n_235),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_326),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_251),
.A2(n_244),
.B1(n_221),
.B2(n_219),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_253),
.B(n_233),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_262),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_328),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_329),
.B(n_340),
.Y(n_394)
);

OA22x2_ASAP7_75t_L g331 ( 
.A1(n_303),
.A2(n_239),
.B1(n_212),
.B2(n_206),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_331),
.A2(n_299),
.B(n_326),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_224),
.C(n_265),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_333),
.B(n_335),
.C(n_341),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_207),
.C(n_209),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_324),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_216),
.C(n_255),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_346),
.B1(n_367),
.B2(n_297),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_325),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_343),
.B(n_350),
.Y(n_397)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_345),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_216),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_348),
.B(n_349),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_280),
.B(n_216),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_279),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_351),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_262),
.C(n_271),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_354),
.C(n_326),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_290),
.B(n_262),
.C(n_271),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_356),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_276),
.B(n_271),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_276),
.B(n_304),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_368),
.Y(n_389)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_292),
.Y(n_359)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_228),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_362),
.Y(n_375)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_301),
.Y(n_361)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_279),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_301),
.Y(n_363)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_288),
.Y(n_364)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_215),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_366),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_279),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_302),
.A2(n_215),
.B1(n_315),
.B2(n_323),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_273),
.B(n_282),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_369),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_299),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_299),
.Y(n_390)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_298),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_371),
.B(n_278),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_355),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_373),
.B(n_382),
.Y(n_422)
);

OAI32xp33_ASAP7_75t_L g374 ( 
.A1(n_334),
.A2(n_296),
.A3(n_294),
.B1(n_275),
.B2(n_322),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_374),
.B(n_395),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_344),
.A2(n_317),
.B1(n_293),
.B2(n_306),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_377),
.A2(n_393),
.B1(n_396),
.B2(n_400),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_330),
.A2(n_313),
.B(n_289),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_379),
.A2(n_401),
.B(n_402),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_349),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_330),
.A2(n_272),
.B(n_295),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_383),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_336),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_391),
.C(n_403),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_388),
.A2(n_339),
.B1(n_340),
.B2(n_368),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_390),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_344),
.A2(n_296),
.B1(n_291),
.B2(n_308),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_334),
.A2(n_322),
.B1(n_308),
.B2(n_281),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_337),
.A2(n_367),
.B1(n_339),
.B2(n_356),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_329),
.A2(n_295),
.B(n_274),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_332),
.B(n_318),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_364),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_312),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_342),
.A2(n_307),
.B1(n_312),
.B2(n_283),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_406),
.A2(n_346),
.B1(n_363),
.B2(n_361),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_331),
.A2(n_338),
.B(n_352),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_393),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_408),
.A2(n_415),
.B1(n_421),
.B2(n_436),
.Y(n_440)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_381),
.Y(n_409)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_412),
.A2(n_419),
.B1(n_431),
.B2(n_433),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_401),
.A2(n_358),
.B1(n_341),
.B2(n_347),
.Y(n_415)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_416),
.Y(n_451)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_381),
.Y(n_417)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_377),
.A2(n_343),
.B1(n_354),
.B2(n_331),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_378),
.B(n_347),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_420),
.B(n_427),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_394),
.A2(n_333),
.B1(n_331),
.B2(n_335),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_336),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_438),
.C(n_376),
.Y(n_443)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_424),
.Y(n_453)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_425),
.Y(n_457)
);

NOR4xp25_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_350),
.C(n_362),
.D(n_366),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_430),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_378),
.B(n_370),
.Y(n_427)
);

BUFx5_ASAP7_75t_L g429 ( 
.A(n_399),
.Y(n_429)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_429),
.Y(n_458)
);

NOR4xp25_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_353),
.C(n_352),
.D(n_331),
.Y(n_430)
);

NOR3xp33_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_309),
.C(n_299),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_357),
.Y(n_432)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_373),
.B(n_345),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_390),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_434),
.A2(n_397),
.B(n_372),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_382),
.B(n_371),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_435),
.A2(n_395),
.B(n_405),
.Y(n_463)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_386),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_437),
.A2(n_392),
.B1(n_387),
.B2(n_386),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_376),
.B(n_359),
.Y(n_438)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_450),
.C(n_454),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_444),
.A2(n_445),
.B(n_448),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_416),
.A2(n_383),
.B(n_379),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_408),
.A2(n_407),
.B1(n_396),
.B2(n_393),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_447),
.A2(n_462),
.B1(n_422),
.B2(n_412),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_418),
.A2(n_375),
.B(n_380),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_391),
.C(n_400),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_413),
.B(n_372),
.C(n_403),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_407),
.C(n_402),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_456),
.C(n_459),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_407),
.C(n_374),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_421),
.B(n_387),
.C(n_398),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_410),
.A2(n_393),
.B1(n_406),
.B2(n_398),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_460),
.A2(n_434),
.B1(n_428),
.B2(n_433),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_415),
.B(n_392),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_424),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_418),
.A2(n_405),
.B1(n_404),
.B2(n_351),
.Y(n_462)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_463),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_414),
.B(n_369),
.C(n_399),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_464),
.B(n_427),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_466),
.B(n_475),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_464),
.Y(n_467)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_467),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_468),
.A2(n_478),
.B1(n_485),
.B2(n_486),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_428),
.Y(n_472)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_472),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_422),
.Y(n_474)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_411),
.Y(n_475)
);

XNOR2x1_ASAP7_75t_L g476 ( 
.A(n_439),
.B(n_410),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_476),
.B(n_477),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_411),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_460),
.A2(n_430),
.B1(n_419),
.B2(n_432),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_479),
.A2(n_457),
.B1(n_446),
.B2(n_458),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_442),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_482),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_459),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_448),
.B(n_435),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_488),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_450),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_487),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_441),
.A2(n_426),
.B1(n_436),
.B2(n_437),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_439),
.A2(n_409),
.B1(n_425),
.B2(n_417),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_447),
.A2(n_440),
.B1(n_444),
.B2(n_453),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_456),
.C(n_461),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_494),
.C(n_495),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_473),
.B(n_440),
.C(n_445),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_462),
.C(n_453),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_465),
.C(n_463),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_498),
.B(n_500),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_465),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_501),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_458),
.C(n_457),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_470),
.B(n_449),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_502),
.A2(n_468),
.B1(n_469),
.B2(n_474),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_470),
.A2(n_319),
.B(n_429),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_506),
.B(n_486),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_467),
.B(n_283),
.C(n_284),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_507),
.B(n_487),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_502),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_512),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_501),
.A2(n_485),
.B(n_478),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_510),
.A2(n_514),
.B(n_522),
.Y(n_529)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_493),
.Y(n_511)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_511),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_471),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_513),
.B(n_517),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_476),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_516),
.B(n_519),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_479),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_505),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_504),
.A2(n_469),
.B1(n_472),
.B2(n_307),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_489),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_507),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_503),
.A2(n_472),
.B(n_319),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_531),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_510),
.A2(n_497),
.B(n_511),
.Y(n_525)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_525),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_509),
.A2(n_494),
.B(n_498),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_534),
.Y(n_538)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_530),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_520),
.B(n_495),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_515),
.B(n_496),
.C(n_491),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_533),
.B(n_521),
.C(n_490),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_514),
.A2(n_505),
.B1(n_490),
.B2(n_499),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_525),
.A2(n_518),
.B1(n_508),
.B2(n_520),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_537),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_532),
.B(n_515),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_539),
.B(n_540),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_523),
.A2(n_522),
.B1(n_519),
.B2(n_521),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_541),
.B(n_544),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_516),
.Y(n_543)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_543),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_533),
.B(n_284),
.C(n_277),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_538),
.A2(n_529),
.B(n_528),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_548),
.A2(n_549),
.B(n_309),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_538),
.A2(n_536),
.B(n_535),
.Y(n_549)
);

AOI322xp5_ASAP7_75t_L g550 ( 
.A1(n_537),
.A2(n_526),
.A3(n_534),
.B1(n_524),
.B2(n_529),
.C1(n_532),
.C2(n_319),
.Y(n_550)
);

AOI322xp5_ASAP7_75t_L g552 ( 
.A1(n_550),
.A2(n_545),
.A3(n_310),
.B1(n_546),
.B2(n_277),
.C1(n_287),
.C2(n_551),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_552),
.A2(n_553),
.B(n_554),
.Y(n_556)
);

OAI321xp33_ASAP7_75t_L g553 ( 
.A1(n_545),
.A2(n_542),
.A3(n_543),
.B1(n_544),
.B2(n_539),
.C(n_540),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_547),
.A2(n_309),
.B(n_310),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_555),
.B(n_310),
.C(n_278),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_556),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_558),
.B(n_559),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_556),
.B(n_288),
.Y(n_559)
);


endmodule