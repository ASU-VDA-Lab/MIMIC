module fake_jpeg_24732_n_316 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_31),
.Y(n_53)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_52),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_31),
.Y(n_76)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_23),
.B1(n_30),
.B2(n_19),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_33),
.B1(n_31),
.B2(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_63),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_67),
.B1(n_20),
.B2(n_34),
.Y(n_108)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_29),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_30),
.B1(n_23),
.B2(n_33),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_35),
.B1(n_32),
.B2(n_28),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_75),
.Y(n_110)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_49),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_74),
.B(n_76),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_21),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_94),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_41),
.B(n_24),
.C(n_16),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_78),
.B(n_96),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_81),
.Y(n_121)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_95),
.B1(n_108),
.B2(n_20),
.Y(n_112)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_86),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_24),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_42),
.B1(n_33),
.B2(n_16),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_93),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_21),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_16),
.B(n_27),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_24),
.B1(n_27),
.B2(n_40),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_104),
.B1(n_107),
.B2(n_22),
.Y(n_113)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_101),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_0),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_77),
.Y(n_111)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_26),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_26),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_48),
.A2(n_27),
.B1(n_42),
.B2(n_34),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_62),
.A2(n_41),
.B1(n_26),
.B2(n_21),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_106),
.A2(n_103),
.B1(n_94),
.B2(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_111),
.B(n_113),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_112),
.A2(n_128),
.B1(n_22),
.B2(n_18),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_136),
.B1(n_71),
.B2(n_83),
.Y(n_144)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_127),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_106),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_36),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_88),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_22),
.B1(n_18),
.B2(n_17),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_134),
.Y(n_150)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_87),
.A2(n_26),
.B1(n_22),
.B2(n_18),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_108),
.A3(n_78),
.B1(n_100),
.B2(n_107),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_152),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_SL g179 ( 
.A1(n_142),
.A2(n_120),
.B(n_122),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_93),
.C(n_70),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_119),
.C(n_109),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_147),
.B1(n_151),
.B2(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_154),
.Y(n_191)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_80),
.B1(n_71),
.B2(n_79),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_113),
.B1(n_136),
.B2(n_125),
.Y(n_151)
);

AOI22x1_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_84),
.B1(n_80),
.B2(n_71),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_159),
.B1(n_162),
.B2(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_76),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_170),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_112),
.A2(n_86),
.B1(n_72),
.B2(n_98),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_101),
.B1(n_70),
.B2(n_92),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_158),
.A2(n_132),
.B1(n_130),
.B2(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_165),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_110),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

OAI22x1_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_90),
.B1(n_18),
.B2(n_17),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_109),
.B(n_10),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_119),
.A2(n_17),
.B1(n_69),
.B2(n_15),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_SL g168 ( 
.A(n_120),
.B(n_17),
.C(n_15),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_168),
.B(n_169),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_174),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_173),
.A2(n_181),
.B1(n_4),
.B2(n_5),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_135),
.C(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_175),
.B(n_177),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_158),
.C(n_154),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_179),
.A2(n_1),
.B(n_2),
.Y(n_213)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_180),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_122),
.B1(n_124),
.B2(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_182),
.B(n_197),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_117),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_185),
.B(n_195),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_126),
.C(n_117),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_124),
.B1(n_126),
.B2(n_105),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_196),
.B1(n_141),
.B2(n_146),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_148),
.B(n_14),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_140),
.A2(n_144),
.B1(n_142),
.B2(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_145),
.B(n_0),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_214),
.B1(n_222),
.B2(n_225),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_166),
.B(n_2),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_209),
.B(n_213),
.Y(n_234)
);

HAxp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_139),
.CON(n_209),
.SN(n_209)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_164),
.Y(n_217)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_1),
.B(n_3),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_1),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_14),
.B(n_13),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_4),
.B(n_5),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_223),
.B1(n_226),
.B2(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_183),
.B1(n_182),
.B2(n_178),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_174),
.C(n_199),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_233),
.C(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_216),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_202),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_244),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_247),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_172),
.C(n_190),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_183),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_243),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_173),
.C(n_171),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_175),
.B1(n_189),
.B2(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_177),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_212),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_SL g245 ( 
.A1(n_207),
.A2(n_178),
.B(n_186),
.C(n_6),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_214),
.B(n_227),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_197),
.B1(n_186),
.B2(n_184),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_241),
.B1(n_235),
.B2(n_238),
.Y(n_265)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_221),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_250),
.A2(n_230),
.B1(n_240),
.B2(n_245),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_217),
.B1(n_208),
.B2(n_215),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_254),
.B1(n_267),
.B2(n_249),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_216),
.B(n_219),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_264),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_213),
.B(n_225),
.Y(n_254)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_212),
.C(n_205),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_261),
.C(n_240),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_205),
.C(n_223),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_230),
.Y(n_262)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_211),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_236),
.A2(n_226),
.B1(n_211),
.B2(n_210),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_268),
.A2(n_279),
.B1(n_280),
.B2(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_252),
.C(n_265),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_260),
.C(n_257),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_274),
.C(n_263),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_243),
.C(n_203),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_245),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_276),
.B(n_258),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_245),
.C(n_12),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_250),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_281),
.B(n_251),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_292),
.B(n_276),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_263),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_268),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_286),
.C(n_270),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_255),
.C(n_253),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_291),
.C(n_272),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_290),
.B(n_275),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_259),
.C(n_267),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_259),
.B(n_264),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_294),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_269),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_282),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_299),
.Y(n_303)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_300),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_280),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_302),
.A2(n_304),
.B1(n_294),
.B2(n_297),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_298),
.B(n_296),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_279),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_309),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_305),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_306),
.C(n_301),
.Y(n_312)
);

AOI21x1_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_311),
.B(n_305),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_285),
.B1(n_284),
.B2(n_11),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_11),
.C(n_7),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_7),
.B1(n_8),
.B2(n_309),
.Y(n_316)
);


endmodule