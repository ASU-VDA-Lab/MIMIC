module fake_jpeg_11697_n_650 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_650);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_650;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_18),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_65),
.B(n_67),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_66),
.A2(n_33),
.B1(n_61),
.B2(n_37),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_8),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_68),
.B(n_84),
.Y(n_161)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_70),
.B(n_76),
.Y(n_143)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_75),
.B(n_104),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_78),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_79),
.B(n_82),
.Y(n_152)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_80),
.Y(n_180)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_83),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_7),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_85),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_90),
.Y(n_216)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_22),
.B(n_9),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_94),
.B(n_111),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_95),
.B(n_110),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_102),
.Y(n_197)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_26),
.B(n_9),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

BUFx24_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_9),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_113),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_25),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_26),
.B(n_9),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_48),
.B(n_6),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_23),
.Y(n_114)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_41),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_124),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_32),
.B(n_11),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_120),
.B(n_61),
.Y(n_172)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_121),
.Y(n_215)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_42),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_42),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_125),
.B(n_128),
.Y(n_202)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_126),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_23),
.Y(n_128)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_33),
.Y(n_129)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_147),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_167),
.A2(n_59),
.B1(n_47),
.B2(n_54),
.Y(n_264)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_172),
.B(n_177),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_75),
.B(n_57),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_173),
.B(n_176),
.Y(n_234)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_175),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_109),
.B(n_30),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_113),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_105),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_194),
.Y(n_230)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_63),
.Y(n_184)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_184),
.Y(n_263)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_74),
.Y(n_190)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_190),
.Y(n_276)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_64),
.Y(n_193)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_89),
.B(n_32),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_129),
.B(n_31),
.Y(n_195)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_195),
.B(n_57),
.Y(n_287)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_73),
.Y(n_196)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_196),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_107),
.B(n_51),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_198),
.B(n_203),
.Y(n_221)
);

HAxp5_ASAP7_75t_SL g199 ( 
.A(n_102),
.B(n_51),
.CON(n_199),
.SN(n_199)
);

NOR2x1_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_210),
.Y(n_233)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_76),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_82),
.B(n_54),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_205),
.B(n_207),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_81),
.B(n_126),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_92),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_128),
.B(n_49),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_78),
.Y(n_208)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_105),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_86),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_97),
.B(n_49),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_99),
.Y(n_211)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_85),
.Y(n_212)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_212),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_71),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_213),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_77),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_132),
.A2(n_62),
.B1(n_43),
.B2(n_80),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_217),
.Y(n_296)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

INVx6_ASAP7_75t_L g333 ( 
.A(n_218),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_150),
.B(n_27),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_219),
.B(n_222),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_181),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_223),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_144),
.A2(n_123),
.B1(n_127),
.B2(n_130),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_224),
.A2(n_226),
.B1(n_227),
.B2(n_254),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_143),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_225),
.B(n_236),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_161),
.A2(n_106),
.B1(n_118),
.B2(n_116),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_108),
.B1(n_115),
.B2(n_83),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_228),
.Y(n_304)
);

INVx6_ASAP7_75t_SL g229 ( 
.A(n_158),
.Y(n_229)
);

CKINVDCx6p67_ASAP7_75t_R g307 ( 
.A(n_229),
.Y(n_307)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_158),
.Y(n_231)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_235),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_173),
.B(n_53),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_135),
.A2(n_43),
.B1(n_72),
.B2(n_93),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_238),
.A2(n_268),
.B1(n_278),
.B2(n_291),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_103),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_239),
.B(n_241),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_240),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_176),
.B(n_27),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_140),
.B(n_168),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_242),
.B(n_243),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_137),
.B(n_53),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_152),
.B(n_121),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_246),
.B(n_255),
.Y(n_352)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_163),
.Y(n_248)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_248),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_277),
.Y(n_295)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_251),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_149),
.B(n_31),
.C(n_90),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_186),
.C(n_180),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_199),
.A2(n_100),
.B1(n_98),
.B2(n_96),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_183),
.B(n_38),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_256),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_191),
.B(n_38),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_257),
.B(n_261),
.Y(n_312)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_156),
.Y(n_259)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_259),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_146),
.B(n_37),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_136),
.Y(n_262)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_264),
.A2(n_270),
.B1(n_284),
.B2(n_286),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_213),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_265),
.B(n_201),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_157),
.Y(n_266)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_139),
.B(n_47),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_267),
.B(n_292),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_178),
.A2(n_87),
.B1(n_112),
.B2(n_30),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_162),
.A2(n_46),
.B1(n_60),
.B2(n_69),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_159),
.Y(n_271)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_159),
.Y(n_272)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_272),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_157),
.Y(n_273)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_273),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_155),
.A2(n_91),
.B1(n_60),
.B2(n_46),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_275),
.A2(n_280),
.B1(n_188),
.B2(n_145),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_169),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_178),
.A2(n_57),
.B1(n_56),
.B2(n_59),
.Y(n_278)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_179),
.Y(n_279)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_162),
.A2(n_60),
.B1(n_46),
.B2(n_101),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_206),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_281),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_179),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_189),
.A2(n_101),
.B1(n_57),
.B2(n_56),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_134),
.Y(n_285)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_155),
.A2(n_57),
.B1(n_56),
.B2(n_12),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_160),
.B(n_170),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_215),
.B(n_56),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_289),
.B(n_164),
.Y(n_309)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_186),
.Y(n_290)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_180),
.A2(n_56),
.B1(n_154),
.B2(n_214),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_141),
.B(n_0),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_294),
.B(n_298),
.C(n_305),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_234),
.B(n_197),
.Y(n_298)
);

OA22x2_ASAP7_75t_L g387 ( 
.A1(n_302),
.A2(n_319),
.B1(n_339),
.B2(n_341),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_234),
.B(n_142),
.C(n_148),
.Y(n_305)
);

A2O1A1O1Ixp25_ASAP7_75t_L g308 ( 
.A1(n_236),
.A2(n_197),
.B(n_215),
.C(n_147),
.D(n_164),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_308),
.B(n_342),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_314),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_230),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_281),
.A2(n_188),
.B1(n_145),
.B2(n_151),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_249),
.A2(n_164),
.B1(n_138),
.B2(n_131),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_321),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_323),
.B(n_335),
.Y(n_366)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_258),
.Y(n_325)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_328),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_287),
.A2(n_153),
.B(n_133),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_330),
.A2(n_237),
.B(n_276),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_249),
.A2(n_138),
.B1(n_131),
.B2(n_204),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_332),
.A2(n_245),
.B1(n_131),
.B2(n_272),
.Y(n_383)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_243),
.B(n_151),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_257),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_263),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_234),
.B(n_192),
.C(n_165),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_337),
.B(n_344),
.C(n_245),
.Y(n_384)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_247),
.Y(n_338)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_338),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_275),
.A2(n_189),
.B1(n_166),
.B2(n_192),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_250),
.A2(n_166),
.B1(n_165),
.B2(n_204),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_250),
.B(n_193),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_342),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_253),
.B(n_174),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_343),
.B(n_288),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_219),
.B(n_138),
.Y(n_344)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_247),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_350),
.B(n_351),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_354),
.B(n_370),
.Y(n_437)
);

INVx13_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

BUFx12f_ASAP7_75t_L g417 ( 
.A(n_357),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_322),
.A2(n_252),
.B1(n_261),
.B2(n_267),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_358),
.A2(n_376),
.B1(n_388),
.B2(n_398),
.Y(n_436)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_297),
.A2(n_264),
.B1(n_233),
.B2(n_286),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_360),
.A2(n_369),
.B1(n_295),
.B2(n_316),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_299),
.Y(n_362)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_362),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_317),
.B(n_292),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_364),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_241),
.Y(n_364)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_353),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_367),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_297),
.A2(n_233),
.B1(n_221),
.B2(n_218),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_296),
.A2(n_229),
.B1(n_231),
.B2(n_259),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_371),
.A2(n_374),
.B(n_399),
.Y(n_404)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_375),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_335),
.A2(n_220),
.B1(n_232),
.B2(n_279),
.Y(n_376)
);

CKINVDCx10_ASAP7_75t_R g378 ( 
.A(n_307),
.Y(n_378)
);

INVx3_ASAP7_75t_SL g415 ( 
.A(n_378),
.Y(n_415)
);

AND2x2_ASAP7_75t_SL g379 ( 
.A(n_298),
.B(n_232),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_397),
.Y(n_409)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_380),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_274),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_312),
.B(n_285),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_386),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_295),
.Y(n_422)
);

INVx11_ASAP7_75t_L g385 ( 
.A(n_307),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_312),
.B(n_274),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_335),
.A2(n_240),
.B1(n_256),
.B2(n_273),
.Y(n_388)
);

AND2x6_ASAP7_75t_L g389 ( 
.A(n_331),
.B(n_237),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_394),
.Y(n_412)
);

INVx13_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_391),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_244),
.C(n_228),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_396),
.C(n_345),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_296),
.A2(n_301),
.B1(n_316),
.B2(n_293),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g439 ( 
.A1(n_393),
.A2(n_304),
.B1(n_346),
.B2(n_327),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_335),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_300),
.B(n_337),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_313),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_305),
.B(n_282),
.C(n_266),
.Y(n_396)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_294),
.B(n_306),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_348),
.A2(n_271),
.B1(n_283),
.B2(n_269),
.Y(n_398)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_400),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_397),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_403),
.C(n_408),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_303),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_358),
.A2(n_330),
.B1(n_323),
.B2(n_349),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_405),
.A2(n_410),
.B1(n_416),
.B2(n_361),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_342),
.Y(n_408)
);

OAI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_388),
.A2(n_308),
.B1(n_329),
.B2(n_347),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_413),
.B(n_399),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_395),
.A2(n_333),
.B1(n_347),
.B2(n_346),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_385),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_421),
.B(n_428),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_425),
.C(n_433),
.Y(n_445)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_356),
.Y(n_424)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_424),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_295),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_386),
.Y(n_444)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_356),
.Y(n_427)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_378),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_366),
.B(n_333),
.Y(n_429)
);

OAI21xp33_ASAP7_75t_L g459 ( 
.A1(n_429),
.A2(n_431),
.B(n_394),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_366),
.A2(n_345),
.B(n_310),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_430),
.A2(n_439),
.B(n_367),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_366),
.B(n_311),
.Y(n_431)
);

MAJx2_ASAP7_75t_L g433 ( 
.A(n_384),
.B(n_320),
.C(n_318),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_355),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_354),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_435),
.B(n_392),
.C(n_396),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_369),
.A2(n_315),
.B1(n_327),
.B2(n_311),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_440),
.A2(n_376),
.B1(n_371),
.B2(n_398),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_417),
.Y(n_441)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_419),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_442),
.B(n_457),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_444),
.B(n_449),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_446),
.B(n_473),
.C(n_443),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_447),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_448),
.B(n_464),
.Y(n_487)
);

OAI22xp33_ASAP7_75t_SL g480 ( 
.A1(n_450),
.A2(n_476),
.B1(n_440),
.B2(n_413),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_431),
.A2(n_390),
.B(n_374),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_451),
.A2(n_404),
.B(n_429),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_412),
.B(n_389),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_452),
.A2(n_465),
.B(n_466),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_406),
.B(n_382),
.Y(n_455)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_455),
.Y(n_484)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_424),
.Y(n_456)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_456),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_429),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_418),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_468),
.Y(n_483)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_459),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_405),
.A2(n_379),
.B1(n_390),
.B2(n_361),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_460),
.A2(n_438),
.B1(n_423),
.B2(n_420),
.Y(n_504)
);

INVx13_ASAP7_75t_L g461 ( 
.A(n_417),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_461),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_406),
.B(n_363),
.Y(n_462)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_462),
.Y(n_495)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_427),
.Y(n_463)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_463),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_418),
.B(n_364),
.Y(n_464)
);

AOI32xp33_ASAP7_75t_L g466 ( 
.A1(n_411),
.A2(n_379),
.A3(n_365),
.B1(n_362),
.B2(n_355),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_426),
.B(n_379),
.Y(n_468)
);

A2O1A1Ixp33_ASAP7_75t_L g469 ( 
.A1(n_409),
.A2(n_359),
.B(n_372),
.C(n_377),
.Y(n_469)
);

O2A1O1Ixp33_ASAP7_75t_L g482 ( 
.A1(n_469),
.A2(n_409),
.B(n_404),
.C(n_430),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_416),
.B(n_368),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_471),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_437),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_403),
.B(n_372),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_472),
.B(n_475),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_402),
.B(n_359),
.C(n_377),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_431),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_436),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_414),
.B(n_368),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_407),
.A2(n_387),
.B1(n_362),
.B2(n_400),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g477 ( 
.A(n_422),
.B(n_380),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_477),
.A2(n_460),
.B(n_452),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_479),
.A2(n_488),
.B(n_500),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_480),
.A2(n_504),
.B1(n_449),
.B2(n_457),
.Y(n_524)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_482),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_447),
.A2(n_407),
.B(n_409),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_489),
.B(n_497),
.C(n_503),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_490),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_496),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_446),
.B(n_443),
.C(n_445),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_467),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_498),
.B(n_507),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_458),
.A2(n_435),
.B1(n_438),
.B2(n_433),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_499),
.A2(n_415),
.B1(n_401),
.B2(n_304),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_451),
.A2(n_425),
.B(n_408),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_444),
.B(n_432),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_501),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_448),
.B(n_432),
.Y(n_502)
);

OAI21xp33_ASAP7_75t_L g521 ( 
.A1(n_502),
.A2(n_506),
.B(n_470),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_445),
.B(n_473),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_471),
.B(n_414),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_464),
.B(n_420),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_472),
.B(n_320),
.C(n_326),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_509),
.C(n_453),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_468),
.B(n_375),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_499),
.B(n_462),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_512),
.B(n_529),
.Y(n_547)
);

NAND2x1_ASAP7_75t_SL g515 ( 
.A(n_494),
.B(n_474),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_515),
.A2(n_537),
.B(n_538),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_489),
.B(n_503),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_516),
.B(n_519),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_487),
.B(n_442),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_518),
.B(n_520),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_455),
.Y(n_520)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_521),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_524),
.A2(n_541),
.B1(n_493),
.B2(n_502),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_481),
.A2(n_450),
.B1(n_465),
.B2(n_466),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_525),
.A2(n_532),
.B1(n_504),
.B2(n_511),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_506),
.B(n_475),
.Y(n_526)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_526),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_497),
.B(n_463),
.Y(n_527)
);

CKINVDCx14_ASAP7_75t_R g548 ( 
.A(n_527),
.Y(n_548)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_528),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_483),
.B(n_477),
.Y(n_529)
);

XNOR2x1_ASAP7_75t_L g531 ( 
.A(n_509),
.B(n_469),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_531),
.B(n_536),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_481),
.A2(n_456),
.B1(n_454),
.B2(n_453),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_488),
.A2(n_479),
.B(n_494),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_533),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_454),
.C(n_401),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_540),
.C(n_508),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_478),
.A2(n_357),
.B(n_380),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_488),
.A2(n_461),
.B(n_357),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_478),
.A2(n_461),
.B(n_415),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_539),
.B(n_542),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_500),
.B(n_415),
.C(n_326),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_511),
.A2(n_441),
.B1(n_387),
.B2(n_340),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_482),
.A2(n_441),
.B(n_417),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_545),
.A2(n_566),
.B1(n_530),
.B2(n_536),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_525),
.A2(n_490),
.B1(n_484),
.B2(n_485),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_550),
.A2(n_567),
.B1(n_545),
.B2(n_566),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_516),
.B(n_514),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_551),
.B(n_564),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_523),
.A2(n_485),
.B1(n_495),
.B2(n_484),
.Y(n_556)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_556),
.Y(n_571)
);

XNOR2x1_ASAP7_75t_L g586 ( 
.A(n_558),
.B(n_560),
.Y(n_586)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_522),
.Y(n_559)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_559),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_523),
.A2(n_495),
.B1(n_483),
.B2(n_507),
.Y(n_561)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_561),
.Y(n_584)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_522),
.Y(n_562)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_562),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_524),
.A2(n_491),
.B1(n_501),
.B2(n_492),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_563),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_514),
.B(n_496),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_519),
.B(n_493),
.C(n_510),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_565),
.B(n_512),
.C(n_540),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_534),
.A2(n_482),
.B1(n_505),
.B2(n_491),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_532),
.A2(n_505),
.B1(n_510),
.B2(n_492),
.Y(n_567)
);

INVx6_ASAP7_75t_L g568 ( 
.A(n_548),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_568),
.B(n_579),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_570),
.A2(n_582),
.B1(n_587),
.B2(n_417),
.Y(n_599)
);

BUFx12_ASAP7_75t_L g572 ( 
.A(n_557),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_572),
.B(n_574),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_544),
.B(n_542),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_564),
.A2(n_537),
.B(n_539),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_575),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_552),
.A2(n_535),
.B1(n_541),
.B2(n_517),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_577),
.B(n_583),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_544),
.B(n_538),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_578),
.B(n_387),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_553),
.B(n_513),
.C(n_526),
.Y(n_579)
);

NOR3xp33_ASAP7_75t_SL g580 ( 
.A(n_554),
.B(n_530),
.C(n_529),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_580),
.A2(n_547),
.B1(n_515),
.B2(n_549),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_557),
.A2(n_533),
.B(n_513),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_581),
.A2(n_543),
.B(n_549),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_567),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_585),
.B(n_223),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_550),
.A2(n_517),
.B1(n_531),
.B2(n_515),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_589),
.A2(n_595),
.B(n_606),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_586),
.B(n_551),
.C(n_546),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_590),
.B(n_592),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_576),
.A2(n_543),
.B1(n_560),
.B2(n_558),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_591),
.A2(n_596),
.B1(n_587),
.B2(n_578),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_586),
.B(n_546),
.C(n_565),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_594),
.A2(n_597),
.B1(n_589),
.B2(n_595),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_SL g595 ( 
.A1(n_574),
.A2(n_547),
.B(n_528),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_576),
.A2(n_555),
.B1(n_486),
.B2(n_387),
.Y(n_596)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_583),
.B(n_391),
.Y(n_598)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_598),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_599),
.B(n_601),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_569),
.B(n_340),
.C(n_391),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_600),
.B(n_603),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_584),
.A2(n_315),
.B1(n_169),
.B2(n_185),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_605),
.B(n_568),
.Y(n_608)
);

MAJx2_ASAP7_75t_L g606 ( 
.A(n_574),
.B(n_277),
.C(n_251),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_592),
.B(n_571),
.C(n_582),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_607),
.B(n_608),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_602),
.B(n_578),
.C(n_581),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_610),
.B(n_612),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_611),
.B(n_620),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_590),
.B(n_588),
.C(n_573),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_572),
.C(n_580),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_613),
.B(n_612),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g615 ( 
.A1(n_593),
.A2(n_572),
.B1(n_201),
.B2(n_185),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_615),
.A2(n_617),
.B1(n_603),
.B2(n_260),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_596),
.A2(n_283),
.B1(n_269),
.B2(n_260),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_610),
.A2(n_604),
.B(n_597),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_622),
.A2(n_629),
.B(n_630),
.Y(n_638)
);

OAI21xp33_ASAP7_75t_L g623 ( 
.A1(n_614),
.A2(n_599),
.B(n_601),
.Y(n_623)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_623),
.Y(n_636)
);

MAJx2_ASAP7_75t_L g633 ( 
.A(n_626),
.B(n_631),
.C(n_609),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_627),
.B(n_628),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_616),
.B(n_600),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_613),
.A2(n_606),
.B(n_5),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_607),
.B(n_5),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_611),
.B(n_0),
.C(n_1),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_621),
.B(n_609),
.C(n_618),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_632),
.B(n_634),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_633),
.A2(n_624),
.B1(n_631),
.B2(n_13),
.Y(n_640)
);

AOI322xp5_ASAP7_75t_L g634 ( 
.A1(n_623),
.A2(n_619),
.A3(n_617),
.B1(n_13),
.B2(n_15),
.C1(n_4),
.C2(n_17),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_625),
.A2(n_4),
.B(n_14),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_637),
.B(n_624),
.C(n_17),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_640),
.B(n_641),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_635),
.Y(n_642)
);

AOI322xp5_ASAP7_75t_L g643 ( 
.A1(n_642),
.A2(n_635),
.A3(n_636),
.B1(n_638),
.B2(n_17),
.C1(n_3),
.C2(n_2),
.Y(n_643)
);

OA21x2_ASAP7_75t_L g645 ( 
.A1(n_643),
.A2(n_639),
.B(n_1),
.Y(n_645)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_645),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g646 ( 
.A1(n_644),
.A2(n_0),
.B(n_2),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_647),
.A2(n_646),
.B(n_2),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_SL g649 ( 
.A1(n_648),
.A2(n_2),
.B(n_3),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_649),
.A2(n_2),
.B(n_3),
.Y(n_650)
);


endmodule