module fake_jpeg_27319_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_23),
.B(n_24),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_9),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_9),
.C(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_14),
.B(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_13),
.B1(n_16),
.B2(n_21),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_24),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_16),
.B1(n_21),
.B2(n_11),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_39),
.B1(n_17),
.B2(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_20),
.B1(n_22),
.B2(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_31),
.B(n_33),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_11),
.B(n_18),
.Y(n_48)
);

A2O1A1O1Ixp25_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_31),
.B(n_32),
.C(n_22),
.D(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_31),
.B1(n_39),
.B2(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_22),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_26),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_55),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_38),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_50),
.B(n_41),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_59),
.B1(n_62),
.B2(n_33),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_37),
.B1(n_33),
.B2(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_69),
.Y(n_75)
);

XNOR2x1_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_52),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_72),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_71),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_52),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_53),
.B(n_61),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_61),
.C(n_49),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_20),
.B(n_19),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_82),
.B1(n_43),
.B2(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_12),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_60),
.C(n_55),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_22),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_37),
.B1(n_42),
.B2(n_44),
.Y(n_82)
);

A2O1A1O1Ixp25_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_67),
.B(n_69),
.C(n_66),
.D(n_22),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_88),
.A3(n_76),
.B1(n_40),
.B2(n_81),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_1),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_19),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_87),
.A2(n_78),
.B1(n_40),
.B2(n_19),
.Y(n_91)
);

AOI211xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_91),
.B(n_40),
.C(n_3),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_79),
.C(n_75),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_92),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

OAI31xp33_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_90),
.A3(n_6),
.B(n_4),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_91),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

AOI31xp67_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_97),
.A3(n_3),
.B(n_5),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_2),
.B(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_100),
.Y(n_104)
);


endmodule