module fake_jpeg_445_n_542 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_542);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_6),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_50),
.B(n_59),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_21),
.B(n_6),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_63),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_79),
.Y(n_113)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

INVx11_ASAP7_75t_SL g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_13),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_82),
.B(n_13),
.Y(n_126)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_42),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_92),
.Y(n_114)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_36),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_96),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_46),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

NAND2x1_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_28),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_101),
.B(n_116),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_44),
.B1(n_34),
.B2(n_41),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_107),
.A2(n_86),
.B1(n_91),
.B2(n_39),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_51),
.A2(n_39),
.B1(n_35),
.B2(n_27),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_119),
.A2(n_30),
.B1(n_24),
.B2(n_31),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_54),
.B(n_45),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_144),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_67),
.A2(n_18),
.B1(n_43),
.B2(n_31),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_124),
.A2(n_87),
.B1(n_52),
.B2(n_28),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_126),
.B(n_9),
.Y(n_202)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_75),
.B(n_0),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_35),
.B(n_76),
.C(n_24),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_135),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_71),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_69),
.B(n_33),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_88),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_33),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_158),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_53),
.B(n_18),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_153),
.B(n_154),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_56),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_53),
.B(n_47),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_155),
.B(n_161),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_70),
.B(n_41),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_66),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_168),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_72),
.B1(n_68),
.B2(n_74),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_170),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_245)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_171),
.Y(n_243)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_179),
.Y(n_222)
);

CKINVDCx9p33_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

BUFx24_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_102),
.Y(n_179)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_135),
.A2(n_58),
.B1(n_60),
.B2(n_65),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_137),
.A2(n_77),
.B1(n_47),
.B2(n_30),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_188),
.B(n_190),
.Y(n_249)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_120),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_48),
.B1(n_81),
.B2(n_84),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_121),
.B(n_99),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_208),
.Y(n_246)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_106),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_194),
.B(n_196),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_158),
.B(n_34),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_108),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_125),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_198),
.B(n_200),
.Y(n_221)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_206),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_125),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_137),
.A2(n_43),
.B1(n_34),
.B2(n_55),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_139),
.B1(n_143),
.B2(n_130),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_202),
.B(n_203),
.Y(n_250)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_144),
.A2(n_80),
.B1(n_95),
.B2(n_89),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_205),
.A2(n_207),
.B1(n_34),
.B2(n_130),
.Y(n_219)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_211),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_133),
.B(n_34),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_210),
.B(n_115),
.Y(n_239)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_129),
.C(n_160),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_214),
.B(n_227),
.C(n_166),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_219),
.A2(n_242),
.B1(n_170),
.B2(n_207),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_157),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_184),
.B(n_162),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_237),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_184),
.B(n_113),
.CI(n_125),
.CON(n_231),
.SN(n_231)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_231),
.B(n_210),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_236),
.A2(n_132),
.B1(n_173),
.B2(n_199),
.Y(n_267)
);

AO22x2_ASAP7_75t_L g237 ( 
.A1(n_174),
.A2(n_140),
.B1(n_136),
.B2(n_151),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_195),
.A2(n_109),
.B1(n_147),
.B2(n_151),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_197),
.A2(n_136),
.B(n_146),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_258),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_192),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_252),
.B(n_263),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_195),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_255),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_254),
.B(n_256),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_213),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_212),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_249),
.Y(n_258)
);

AO21x2_ASAP7_75t_L g302 ( 
.A1(n_259),
.A2(n_219),
.B(n_242),
.Y(n_302)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_181),
.Y(n_263)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_191),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_264),
.B(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_176),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_217),
.Y(n_266)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_267),
.A2(n_236),
.B(n_233),
.Y(n_287)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_271),
.B(n_190),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_277),
.Y(n_310)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_216),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_275),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_222),
.A2(n_193),
.B1(n_208),
.B2(n_203),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_234),
.B1(n_241),
.B2(n_245),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_249),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_217),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_281),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_250),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_280),
.B(n_243),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_179),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_249),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_172),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_285),
.B(n_304),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_287),
.A2(n_295),
.B(n_301),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_292),
.A2(n_282),
.B1(n_277),
.B2(n_265),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_276),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_294),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_278),
.A2(n_230),
.B1(n_233),
.B2(n_222),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_268),
.A2(n_222),
.B1(n_235),
.B2(n_239),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_297),
.A2(n_305),
.B1(n_309),
.B2(n_311),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_268),
.A2(n_248),
.B(n_237),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_302),
.A2(n_305),
.B1(n_301),
.B2(n_309),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_254),
.A2(n_231),
.B(n_237),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_268),
.A2(n_237),
.B(n_247),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_268),
.A2(n_237),
.B1(n_234),
.B2(n_238),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_307),
.B(n_280),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_259),
.A2(n_240),
.B1(n_215),
.B2(n_232),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_255),
.A2(n_240),
.B1(n_215),
.B2(n_232),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_257),
.A2(n_168),
.B(n_244),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_281),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_258),
.A2(n_244),
.B1(n_165),
.B2(n_204),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_313),
.A2(n_275),
.B1(n_273),
.B2(n_270),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_271),
.C(n_253),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_316),
.B(n_320),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_349),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_299),
.B(n_252),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_288),
.B(n_271),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_321),
.B(n_302),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_310),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_334),
.B1(n_335),
.B2(n_338),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_285),
.B(n_262),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_323),
.B(n_330),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_324),
.A2(n_329),
.B1(n_341),
.B2(n_342),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_SL g325 ( 
.A1(n_304),
.A2(n_264),
.B(n_267),
.C(n_275),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_339),
.Y(n_353)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_326),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_336),
.C(n_298),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_294),
.A2(n_264),
.B1(n_279),
.B2(n_266),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_256),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_263),
.Y(n_333)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_261),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_229),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_337),
.B(n_322),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_310),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_299),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_340),
.B(n_343),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_302),
.A2(n_260),
.B1(n_274),
.B2(n_272),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_291),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_298),
.B(n_274),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_345),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_292),
.A2(n_302),
.B1(n_303),
.B2(n_284),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_302),
.A2(n_272),
.B1(n_269),
.B2(n_220),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_290),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_364),
.C(n_319),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_284),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_361),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_317),
.A2(n_287),
.B1(n_283),
.B2(n_295),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_358),
.A2(n_368),
.B1(n_325),
.B2(n_335),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_316),
.B(n_283),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_360),
.B(n_374),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_297),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_312),
.C(n_311),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_329),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_365),
.B(n_366),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_344),
.Y(n_366)
);

AND2x4_ASAP7_75t_SL g369 ( 
.A(n_318),
.B(n_313),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_369),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_339),
.Y(n_370)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_302),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_380),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_320),
.B(n_229),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_223),
.Y(n_375)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_375),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_376),
.Y(n_386)
);

AOI322xp5_ASAP7_75t_SL g377 ( 
.A1(n_338),
.A2(n_290),
.A3(n_270),
.B1(n_273),
.B2(n_216),
.C1(n_293),
.C2(n_289),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_383),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_308),
.Y(n_378)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_378),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_347),
.A2(n_293),
.B(n_308),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_379),
.A2(n_162),
.B(n_118),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_317),
.B(n_300),
.Y(n_381)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_381),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_334),
.B(n_300),
.Y(n_382)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_382),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_326),
.B(n_182),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_398),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_361),
.B(n_345),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_405),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_319),
.C(n_347),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_399),
.C(n_413),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_362),
.A2(n_346),
.B1(n_325),
.B2(n_341),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_395),
.A2(n_131),
.B1(n_159),
.B2(n_156),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_350),
.A2(n_325),
.B1(n_327),
.B2(n_342),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_396),
.A2(n_407),
.B1(n_362),
.B2(n_408),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_357),
.B(n_331),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_343),
.C(n_340),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_178),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_403),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_358),
.B(n_325),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_350),
.A2(n_177),
.B(n_206),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_406),
.A2(n_408),
.B(n_139),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_367),
.A2(n_167),
.B1(n_185),
.B2(n_142),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_189),
.Y(n_409)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_409),
.Y(n_416)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_410),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_209),
.Y(n_411)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_411),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_364),
.B(n_226),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_369),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_359),
.B(n_188),
.C(n_169),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_359),
.B(n_128),
.C(n_115),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_379),
.C(n_378),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_415),
.A2(n_427),
.B1(n_428),
.B2(n_435),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_396),
.A2(n_367),
.B1(n_365),
.B2(n_350),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_418),
.A2(n_419),
.B1(n_426),
.B2(n_431),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_384),
.A2(n_355),
.B1(n_353),
.B2(n_373),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_433),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_404),
.A2(n_353),
.B1(n_373),
.B2(n_368),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_371),
.C(n_354),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_432),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_401),
.A2(n_356),
.B1(n_363),
.B2(n_352),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_391),
.B(n_382),
.C(n_369),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_128),
.C(n_110),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_434),
.B(n_143),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_436),
.A2(n_407),
.B1(n_406),
.B2(n_390),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_226),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_402),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_118),
.Y(n_438)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_399),
.C(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_387),
.Y(n_439)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_439),
.Y(n_450)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_393),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_110),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_392),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_441),
.B(n_398),
.Y(n_444)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_460),
.Y(n_466)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_444),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_445),
.A2(n_418),
.B1(n_421),
.B2(n_416),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_446),
.B(n_451),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_419),
.A2(n_405),
.B(n_402),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_448),
.A2(n_455),
.B(n_433),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_395),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_417),
.A2(n_385),
.B1(n_397),
.B2(n_413),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_452),
.B(n_458),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_422),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_462),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_422),
.A2(n_414),
.B(n_211),
.Y(n_455)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_456),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_424),
.B(n_437),
.C(n_423),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_420),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_459),
.B(n_461),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_438),
.B(n_117),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_426),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_417),
.A2(n_142),
.B1(n_156),
.B2(n_159),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_463),
.A2(n_132),
.B1(n_109),
.B2(n_111),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_424),
.B(n_432),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_122),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_482),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_469),
.A2(n_471),
.B1(n_127),
.B2(n_100),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_453),
.C(n_464),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_470),
.B(n_479),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_457),
.A2(n_436),
.B1(n_425),
.B2(n_434),
.Y(n_471)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_450),
.Y(n_473)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_473),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_475),
.B(n_97),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_122),
.C(n_111),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_147),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_484),
.Y(n_495)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_450),
.Y(n_481)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_481),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_131),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_449),
.Y(n_483)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_483),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_442),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_488),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_468),
.A2(n_448),
.B(n_442),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_486),
.A2(n_497),
.B1(n_473),
.B2(n_479),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_451),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_469),
.A2(n_443),
.B(n_460),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_490),
.A2(n_500),
.B(n_17),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_478),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_499),
.Y(n_510)
);

OAI21xp33_ASAP7_75t_L g493 ( 
.A1(n_466),
.A2(n_9),
.B(n_10),
.Y(n_493)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_493),
.Y(n_509)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_494),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_466),
.A2(n_127),
.B(n_97),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_498),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_7),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_471),
.A2(n_46),
.B(n_17),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_474),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_503),
.B(n_506),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_474),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_505),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_487),
.B(n_472),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_494),
.A2(n_496),
.B1(n_489),
.B2(n_501),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_507),
.A2(n_10),
.B(n_9),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_495),
.B(n_472),
.Y(n_508)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_508),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_482),
.C(n_16),
.Y(n_511)
);

AOI31xp33_ASAP7_75t_L g517 ( 
.A1(n_511),
.A2(n_493),
.A3(n_497),
.B(n_7),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_512),
.A2(n_5),
.B(n_1),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_490),
.B(n_16),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_509),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_517),
.A2(n_518),
.B1(n_521),
.B2(n_525),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_502),
.B(n_5),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_519),
.B(n_4),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_505),
.B(n_46),
.C(n_5),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_504),
.Y(n_527)
);

AOI21x1_ASAP7_75t_L g524 ( 
.A1(n_513),
.A2(n_10),
.B(n_8),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_524),
.A2(n_509),
.B(n_510),
.Y(n_528)
);

AO21x1_ASAP7_75t_L g526 ( 
.A1(n_516),
.A2(n_522),
.B(n_523),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_526),
.A2(n_529),
.B(n_530),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_528),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_523),
.A2(n_514),
.B(n_511),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_0),
.Y(n_530)
);

NOR3xp33_ASAP7_75t_SL g533 ( 
.A(n_532),
.B(n_0),
.C(n_1),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_533),
.B(n_535),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_526),
.A2(n_0),
.B(n_1),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_534),
.B(n_531),
.C(n_1),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_536),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_537),
.C(n_2),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_541)
);

NAND3xp33_ASAP7_75t_SL g542 ( 
.A(n_541),
.B(n_3),
.C(n_4),
.Y(n_542)
);


endmodule