module fake_ibex_882_n_3243 (n_151, n_85, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_13, n_122, n_523, n_116, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_355, n_474, n_594, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_536, n_352, n_290, n_558, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_267, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3243);

input n_151;
input n_85;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_594;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_536;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_267;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3243;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2498;
wire n_1802;
wire n_2235;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_930;
wire n_1044;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3168;
wire n_667;
wire n_884;
wire n_2396;
wire n_3135;
wire n_850;
wire n_3175;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_3192;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_3242;
wire n_1654;
wire n_2995;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_2373;
wire n_630;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_2987;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3203;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_3117;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3091;
wire n_3006;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3055;
wire n_1633;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_3214;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3003;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_2252;
wire n_1982;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_607;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_615;
wire n_2905;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1539;
wire n_712;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3167;
wire n_997;
wire n_2308;
wire n_3238;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_634;
wire n_991;
wire n_1331;
wire n_1223;
wire n_961;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_2862;
wire n_3100;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_1952;
wire n_785;
wire n_2180;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_604;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_768;
wire n_839;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2251;
wire n_722;
wire n_2012;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1871;
wire n_1642;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_2818;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2675;
wire n_2417;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_885;
wire n_1530;
wire n_3215;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_1256;
wire n_2798;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3109;
wire n_1961;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_3104;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_682;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_3230;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_1532;
wire n_791;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_1488;
wire n_849;
wire n_980;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3207;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_3124;
wire n_999;
wire n_2634;
wire n_2982;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_635;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_783;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2618;
wire n_2303;
wire n_2653;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3114;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2302;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_2066;
wire n_1719;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_866;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_3195;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_2282;
wire n_970;
wire n_2673;
wire n_2430;
wire n_921;
wire n_2676;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_1506;

INVx1_ASAP7_75t_L g599 ( 
.A(n_209),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_186),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_225),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_145),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_531),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_264),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_376),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_270),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_41),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_304),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_525),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_546),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_275),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_512),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_239),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_77),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_156),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_297),
.Y(n_616)
);

CKINVDCx16_ASAP7_75t_R g617 ( 
.A(n_407),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_192),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_41),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_310),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_67),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_43),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_340),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_298),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_518),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_47),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_174),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_517),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_145),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_554),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_580),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_286),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_153),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_475),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_470),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_59),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_590),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_576),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_414),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_246),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_1),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_505),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_252),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_163),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_83),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_407),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_237),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_401),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_176),
.Y(n_649)
);

CKINVDCx16_ASAP7_75t_R g650 ( 
.A(n_208),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_289),
.Y(n_651)
);

INVxp33_ASAP7_75t_R g652 ( 
.A(n_548),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_542),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_474),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_387),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_506),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_545),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_343),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_31),
.Y(n_659)
);

CKINVDCx14_ASAP7_75t_R g660 ( 
.A(n_355),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_514),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_241),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_541),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_116),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_21),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_589),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_444),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_345),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_491),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_47),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_195),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_189),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_585),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_520),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_372),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_483),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_235),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_248),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_91),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_586),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_367),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_400),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_328),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_261),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_56),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_320),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_521),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_451),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_411),
.Y(n_689)
);

BUFx10_ASAP7_75t_L g690 ( 
.A(n_89),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_398),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_551),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_7),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_184),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_234),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_294),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_348),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_116),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_20),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_318),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_592),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_396),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_507),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_562),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_435),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_169),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_467),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_335),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_148),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_273),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_217),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_504),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_49),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_530),
.Y(n_714)
);

CKINVDCx14_ASAP7_75t_R g715 ( 
.A(n_410),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_495),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_187),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_394),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_415),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_28),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_394),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_117),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_60),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_225),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_28),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_282),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_11),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_202),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_104),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_410),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_10),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_199),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_267),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_428),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_111),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_56),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_91),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_367),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_472),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_34),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_359),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_575),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_125),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_238),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_131),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_257),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_11),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_579),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_120),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_527),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_502),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_351),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_42),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_82),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_44),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_560),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_138),
.Y(n_757)
);

INVx1_ASAP7_75t_SL g758 ( 
.A(n_362),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_236),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_425),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_88),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_265),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_123),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_478),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_205),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_258),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_365),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_473),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_468),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_154),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_240),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_203),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_101),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_50),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_182),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_44),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_29),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_264),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_564),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_133),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_14),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_529),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_398),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_295),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_533),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_23),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_226),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_289),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_125),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_164),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_78),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_572),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_6),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_370),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_209),
.Y(n_795)
);

BUFx10_ASAP7_75t_L g796 ( 
.A(n_559),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_567),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_233),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_189),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_306),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_318),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_390),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_497),
.Y(n_803)
);

BUFx10_ASAP7_75t_L g804 ( 
.A(n_565),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_2),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_231),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_255),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_200),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_261),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_247),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_183),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_124),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_503),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_26),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_115),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_532),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_131),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_210),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_496),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_385),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_45),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_199),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_427),
.Y(n_823)
);

CKINVDCx14_ASAP7_75t_R g824 ( 
.A(n_509),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_487),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_301),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_246),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_31),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_64),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_411),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_516),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_435),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_561),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_239),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_12),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_10),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_340),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_347),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_232),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_342),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_51),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_224),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_138),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_183),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_124),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_218),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_372),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_24),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_445),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_544),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_33),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_320),
.Y(n_852)
);

CKINVDCx14_ASAP7_75t_R g853 ( 
.A(n_2),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_373),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_381),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_238),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_185),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_129),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_260),
.Y(n_859)
);

BUFx10_ASAP7_75t_L g860 ( 
.A(n_74),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_418),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_389),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_494),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_354),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_262),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_292),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_266),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_101),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_176),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_587),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_194),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_237),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_62),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_19),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_94),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_309),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_457),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_13),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_357),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_345),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_216),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_78),
.Y(n_882)
);

BUFx8_ASAP7_75t_SL g883 ( 
.A(n_158),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_110),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_388),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_284),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_595),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_54),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_14),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_353),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_390),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_378),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_308),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_537),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_85),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_36),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_121),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_383),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_207),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_463),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_391),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_4),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_194),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_227),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_593),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_439),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_132),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_13),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_492),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_354),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_400),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_248),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_479),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_383),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_143),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_326),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_388),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_193),
.Y(n_918)
);

BUFx8_ASAP7_75t_SL g919 ( 
.A(n_353),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_180),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_108),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_449),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_12),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_70),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_179),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_279),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_534),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_113),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_17),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_76),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_130),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_574),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_276),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_196),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_375),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_103),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_332),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_540),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_323),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_149),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_182),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_393),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_283),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_59),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_432),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_443),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_302),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_489),
.Y(n_948)
);

CKINVDCx16_ASAP7_75t_R g949 ( 
.A(n_256),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_404),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_207),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_144),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_566),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_215),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_376),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_493),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_71),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_198),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_485),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_569),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_549),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_528),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_260),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_202),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_543),
.Y(n_965)
);

BUFx10_ASAP7_75t_L g966 ( 
.A(n_387),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_563),
.Y(n_967)
);

CKINVDCx12_ASAP7_75t_R g968 ( 
.A(n_379),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_290),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_16),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_4),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_584),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_342),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_448),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_430),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_386),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_153),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_137),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_39),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_107),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_226),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_61),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_88),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_333),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_397),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_344),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_539),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_100),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_171),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_82),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_309),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_612),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_617),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_702),
.Y(n_994)
);

CKINVDCx16_ASAP7_75t_R g995 ( 
.A(n_650),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_702),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_628),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_638),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_767),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_680),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_767),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_692),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_703),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_714),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_769),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_823),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_655),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_823),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_828),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_828),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_851),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_660),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_668),
.B(n_0),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_851),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_809),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_949),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_874),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_638),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_779),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_715),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_853),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_874),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_681),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_813),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_929),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_929),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_883),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_782),
.B(n_0),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_619),
.Y(n_1029)
);

INVxp33_ASAP7_75t_SL g1030 ( 
.A(n_720),
.Y(n_1030)
);

INVxp33_ASAP7_75t_SL g1031 ( 
.A(n_778),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_919),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_968),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_706),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_706),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_968),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_601),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_709),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_709),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_732),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_602),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_639),
.Y(n_1042)
);

INVxp33_ASAP7_75t_SL g1043 ( 
.A(n_937),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_782),
.B(n_1),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_604),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_991),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_732),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_643),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_733),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_654),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_819),
.B(n_3),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_733),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_606),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_607),
.Y(n_1054)
);

INVxp67_ASAP7_75t_SL g1055 ( 
.A(n_735),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_611),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_670),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_819),
.B(n_3),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_735),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_613),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_787),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_814),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_814),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_882),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_882),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_925),
.Y(n_1066)
);

INVxp67_ASAP7_75t_SL g1067 ( 
.A(n_925),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_626),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_683),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_806),
.Y(n_1070)
);

INVxp33_ASAP7_75t_SL g1071 ( 
.A(n_615),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_626),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_629),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_614),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_629),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_700),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_632),
.Y(n_1077)
);

CKINVDCx16_ASAP7_75t_R g1078 ( 
.A(n_608),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_616),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_620),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_726),
.Y(n_1081)
);

CKINVDCx14_ASAP7_75t_R g1082 ( 
.A(n_824),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_788),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_654),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_632),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_821),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_603),
.B(n_5),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_820),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_848),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_645),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_645),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_682),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_866),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_880),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_682),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_896),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_771),
.Y(n_1097)
);

INVxp33_ASAP7_75t_SL g1098 ( 
.A(n_621),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_771),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_836),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_836),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_837),
.Y(n_1102)
);

NAND2xp33_ASAP7_75t_R g1103 ( 
.A(n_627),
.B(n_440),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_R g1104 ( 
.A(n_610),
.B(n_441),
.Y(n_1104)
);

CKINVDCx16_ASAP7_75t_R g1105 ( 
.A(n_608),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_837),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_881),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_603),
.B(n_5),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_881),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_903),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_609),
.B(n_6),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_636),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_608),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_640),
.Y(n_1114)
);

INVxp67_ASAP7_75t_SL g1115 ( 
.A(n_886),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_886),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_944),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_641),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_649),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_977),
.Y(n_1120)
);

OR2x6_ASAP7_75t_L g1121 ( 
.A(n_1012),
.B(n_652),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1030),
.A2(n_600),
.B1(n_605),
.B2(n_599),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1011),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1014),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1017),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_992),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1023),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1022),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1074),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1025),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_997),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1026),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1059),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1034),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1035),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_1029),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1000),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1074),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1074),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1002),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1003),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1004),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1074),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1058),
.B(n_803),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1021),
.B(n_690),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1038),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1005),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1019),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_1082),
.B(n_651),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1050),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1039),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_998),
.B(n_803),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1040),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1024),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1029),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1071),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1050),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1047),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1084),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1078),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_R g1161 ( 
.A(n_1020),
.B(n_658),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1084),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1071),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1098),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1098),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_993),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1070),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_998),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_1042),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1018),
.Y(n_1170)
);

AND3x2_ASAP7_75t_L g1171 ( 
.A(n_1113),
.B(n_852),
.C(n_979),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1030),
.A2(n_600),
.B1(n_605),
.B2(n_599),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1086),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1037),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1018),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1068),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1072),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_993),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_994),
.B(n_996),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1049),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1073),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1007),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1055),
.B(n_978),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1041),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1105),
.B(n_690),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1007),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_999),
.B(n_622),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1075),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1052),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1015),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1096),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1045),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1062),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1077),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1063),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1001),
.B(n_622),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1061),
.B(n_982),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1064),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1015),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1016),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1065),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1067),
.B(n_983),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1066),
.Y(n_1203)
);

AND3x2_ASAP7_75t_L g1204 ( 
.A(n_1006),
.B(n_676),
.C(n_635),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1028),
.B(n_609),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1046),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1085),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_L g1208 ( 
.A(n_1033),
.B(n_625),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1016),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1027),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_995),
.B(n_1008),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1032),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1109),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1042),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1115),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1120),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1090),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1009),
.B(n_690),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1053),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1091),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1092),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1010),
.B(n_860),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1095),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1048),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1097),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1099),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_1054),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1100),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1048),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1101),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1102),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1031),
.B(n_631),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1106),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1107),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_1057),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1031),
.B(n_631),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_1036),
.B(n_1116),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1044),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1057),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1056),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1069),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1013),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1051),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1069),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1076),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_R g1246 ( 
.A(n_1020),
.B(n_664),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1087),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1108),
.A2(n_661),
.B(n_642),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1076),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1111),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1043),
.B(n_988),
.Y(n_1251)
);

BUFx8_ASAP7_75t_L g1252 ( 
.A(n_1043),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1060),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1079),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1080),
.B(n_623),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1112),
.B(n_860),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1104),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1114),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1118),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1119),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1103),
.Y(n_1261)
);

NOR2x1_ASAP7_75t_L g1262 ( 
.A(n_1081),
.B(n_642),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1081),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1083),
.B(n_989),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1083),
.B(n_860),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1088),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1088),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1089),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1089),
.B(n_671),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1093),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1093),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1094),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1094),
.Y(n_1273)
);

NAND2xp33_ASAP7_75t_SL g1274 ( 
.A(n_1110),
.B(n_672),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1110),
.Y(n_1275)
);

INVx4_ASAP7_75t_L g1276 ( 
.A(n_1117),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1117),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1011),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1011),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_992),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1055),
.B(n_973),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1011),
.B(n_661),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_1029),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1011),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1058),
.B(n_688),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_992),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_994),
.B(n_623),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_992),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1011),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1023),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_992),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_992),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1012),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1012),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_992),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1011),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1023),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1011),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_992),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_992),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1055),
.B(n_975),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1011),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1011),
.B(n_688),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1074),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1074),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_998),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1012),
.B(n_966),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1055),
.B(n_984),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1012),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1011),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1011),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_994),
.B(n_624),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_992),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1074),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_992),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1011),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1011),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1058),
.B(n_701),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_992),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1074),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_992),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_992),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_992),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1011),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1023),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1058),
.A2(n_750),
.B(n_701),
.Y(n_1326)
);

BUFx8_ASAP7_75t_L g1327 ( 
.A(n_1012),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_992),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1055),
.B(n_675),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1029),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_R g1331 ( 
.A(n_1082),
.B(n_679),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_998),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1123),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1123),
.Y(n_1334)
);

OR2x6_ASAP7_75t_L g1335 ( 
.A(n_1160),
.B(n_624),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1168),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1128),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1174),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1250),
.A2(n_633),
.B1(n_647),
.B2(n_646),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1290),
.B(n_1242),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1128),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1168),
.Y(n_1342)
);

NAND3xp33_ASAP7_75t_L g1343 ( 
.A(n_1232),
.B(n_685),
.C(n_684),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1168),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1132),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1132),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1238),
.B(n_687),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1278),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1243),
.B(n_750),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1278),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1247),
.B(n_687),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1237),
.B(n_633),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1252),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1213),
.B(n_1215),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1168),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1332),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1290),
.B(n_687),
.Y(n_1357)
);

NOR2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1156),
.B(n_686),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1250),
.A2(n_647),
.B1(n_648),
.B2(n_646),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1316),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1332),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1316),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1218),
.B(n_648),
.Y(n_1363)
);

AO22x2_ASAP7_75t_L g1364 ( 
.A1(n_1122),
.A2(n_1172),
.B1(n_1261),
.B2(n_1196),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1176),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1216),
.B(n_1329),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1191),
.B(n_796),
.Y(n_1367)
);

INVx4_ASAP7_75t_SL g1368 ( 
.A(n_1150),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1176),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1124),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1176),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1176),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1177),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1175),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1232),
.B(n_756),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1236),
.B(n_785),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1326),
.A2(n_665),
.B1(n_677),
.B2(n_662),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1175),
.Y(n_1378)
);

INVx5_ASAP7_75t_L g1379 ( 
.A(n_1150),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1236),
.B(n_785),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1326),
.B(n_792),
.Y(n_1381)
);

INVxp33_ASAP7_75t_L g1382 ( 
.A(n_1127),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1150),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1183),
.B(n_796),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1326),
.B(n_792),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1127),
.B(n_618),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1191),
.B(n_796),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1187),
.A2(n_665),
.B1(n_677),
.B2(n_662),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1150),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1297),
.B(n_966),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1309),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1197),
.B(n_1202),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1177),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1125),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1297),
.B(n_966),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1187),
.B(n_804),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1130),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1279),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1325),
.B(n_705),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1162),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1162),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1253),
.Y(n_1402)
);

INVx3_ASAP7_75t_SL g1403 ( 
.A(n_1163),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_1325),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1248),
.B(n_816),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1285),
.B(n_816),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1284),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1196),
.B(n_804),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1167),
.B(n_691),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1162),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1253),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1285),
.B(n_831),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1289),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1222),
.B(n_678),
.Y(n_1414)
);

BUFx4f_ASAP7_75t_L g1415 ( 
.A(n_1179),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1184),
.Y(n_1416)
);

AND3x4_ASAP7_75t_L g1417 ( 
.A(n_1275),
.B(n_985),
.C(n_977),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1296),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1287),
.A2(n_689),
.B1(n_708),
.B2(n_678),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1206),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1177),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1298),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1167),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1173),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1302),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1281),
.B(n_804),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1173),
.B(n_693),
.Y(n_1427)
);

AND2x6_ASAP7_75t_L g1428 ( 
.A(n_1261),
.B(n_974),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1177),
.Y(n_1429)
);

AND2x6_ASAP7_75t_L g1430 ( 
.A(n_1185),
.B(n_1258),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1258),
.B(n_689),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1293),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1194),
.Y(n_1433)
);

INVx5_ASAP7_75t_L g1434 ( 
.A(n_1162),
.Y(n_1434)
);

AND2x6_ASAP7_75t_L g1435 ( 
.A(n_1259),
.B(n_974),
.Y(n_1435)
);

NAND2xp33_ASAP7_75t_L g1436 ( 
.A(n_1257),
.B(n_630),
.Y(n_1436)
);

INVx4_ASAP7_75t_SL g1437 ( 
.A(n_1194),
.Y(n_1437)
);

BUFx10_ASAP7_75t_L g1438 ( 
.A(n_1164),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1219),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1194),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1301),
.B(n_1308),
.Y(n_1441)
);

AND2x6_ASAP7_75t_L g1442 ( 
.A(n_1260),
.B(n_831),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1294),
.B(n_695),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1170),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1287),
.B(n_634),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1312),
.B(n_637),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1318),
.B(n_1205),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1310),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1318),
.B(n_712),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1240),
.B(n_696),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1211),
.B(n_697),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1145),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1192),
.B(n_698),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1307),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1264),
.B(n_758),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1194),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1252),
.Y(n_1457)
);

INVxp67_ASAP7_75t_SL g1458 ( 
.A(n_1233),
.Y(n_1458)
);

INVx4_ASAP7_75t_SL g1459 ( 
.A(n_1225),
.Y(n_1459)
);

OR2x6_ASAP7_75t_L g1460 ( 
.A(n_1121),
.B(n_708),
.Y(n_1460)
);

AND2x6_ASAP7_75t_L g1461 ( 
.A(n_1254),
.B(n_850),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1205),
.B(n_1144),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1312),
.B(n_653),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1311),
.Y(n_1464)
);

INVx4_ASAP7_75t_L g1465 ( 
.A(n_1233),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1144),
.B(n_905),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1306),
.Y(n_1467)
);

INVx4_ASAP7_75t_L g1468 ( 
.A(n_1225),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1225),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1255),
.B(n_656),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1317),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1225),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1324),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1226),
.Y(n_1474)
);

AND2x6_ASAP7_75t_L g1475 ( 
.A(n_1255),
.B(n_850),
.Y(n_1475)
);

BUFx10_ASAP7_75t_L g1476 ( 
.A(n_1165),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1192),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1226),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1327),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1195),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1327),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1198),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1133),
.B(n_710),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1227),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1226),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1134),
.B(n_863),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1226),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1227),
.B(n_699),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1135),
.B(n_863),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1146),
.B(n_900),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1210),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1212),
.Y(n_1492)
);

NAND2x1p5_ASAP7_75t_L g1493 ( 
.A(n_1256),
.B(n_981),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1161),
.Y(n_1494)
);

BUFx10_ASAP7_75t_L g1495 ( 
.A(n_1204),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1204),
.B(n_710),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1251),
.B(n_657),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1151),
.B(n_900),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1149),
.B(n_711),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1157),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1269),
.B(n_775),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1217),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1220),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1159),
.Y(n_1504)
);

OR2x6_ASAP7_75t_L g1505 ( 
.A(n_1121),
.B(n_717),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1153),
.B(n_909),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1158),
.B(n_909),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1159),
.Y(n_1508)
);

AND2x6_ASAP7_75t_L g1509 ( 
.A(n_1282),
.B(n_927),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1180),
.B(n_927),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1214),
.Y(n_1511)
);

BUFx10_ASAP7_75t_L g1512 ( 
.A(n_1171),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1181),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1189),
.B(n_663),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1221),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1188),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1188),
.A2(n_717),
.B1(n_721),
.B2(n_718),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1207),
.Y(n_1518)
);

NOR2x1p5_ASAP7_75t_L g1519 ( 
.A(n_1276),
.B(n_713),
.Y(n_1519)
);

AND2x6_ASAP7_75t_L g1520 ( 
.A(n_1282),
.B(n_825),
.Y(n_1520)
);

INVx4_ASAP7_75t_L g1521 ( 
.A(n_1171),
.Y(n_1521)
);

BUFx4f_ASAP7_75t_L g1522 ( 
.A(n_1121),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1303),
.B(n_666),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1223),
.Y(n_1524)
);

NAND2xp33_ASAP7_75t_L g1525 ( 
.A(n_1149),
.B(n_667),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1331),
.B(n_719),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1207),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1193),
.B(n_718),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1201),
.B(n_669),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1303),
.B(n_673),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1265),
.Y(n_1531)
);

AND2x6_ASAP7_75t_L g1532 ( 
.A(n_1203),
.B(n_825),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1262),
.B(n_721),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1208),
.B(n_674),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1228),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1224),
.Y(n_1536)
);

INVxp33_ASAP7_75t_L g1537 ( 
.A(n_1161),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1230),
.B(n_723),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1234),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1231),
.B(n_704),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1231),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1126),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_1136),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1331),
.B(n_729),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1152),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1152),
.B(n_707),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1139),
.Y(n_1547)
);

INVx6_ASAP7_75t_L g1548 ( 
.A(n_1129),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1129),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1129),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1246),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1266),
.B(n_716),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1129),
.Y(n_1553)
);

AND2x6_ASAP7_75t_L g1554 ( 
.A(n_1263),
.B(n_723),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1139),
.B(n_739),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1246),
.B(n_731),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1304),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1304),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1131),
.B(n_742),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1138),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1266),
.B(n_748),
.Y(n_1561)
);

BUFx2_ASAP7_75t_L g1562 ( 
.A(n_1276),
.Y(n_1562)
);

INVx5_ASAP7_75t_L g1563 ( 
.A(n_1138),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1138),
.B(n_751),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1272),
.B(n_764),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1138),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1143),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1274),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1143),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1271),
.B(n_724),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1137),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1143),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1143),
.Y(n_1573)
);

AND2x2_ASAP7_75t_SL g1574 ( 
.A(n_1263),
.B(n_724),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1305),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1140),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1141),
.B(n_734),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1305),
.Y(n_1578)
);

BUFx4f_ASAP7_75t_L g1579 ( 
.A(n_1263),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1271),
.B(n_725),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1305),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1142),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1147),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1314),
.B(n_768),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1314),
.Y(n_1585)
);

CKINVDCx16_ASAP7_75t_R g1586 ( 
.A(n_1155),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1272),
.A2(n_725),
.B1(n_728),
.B2(n_727),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1273),
.B(n_797),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1148),
.B(n_737),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1314),
.B(n_833),
.Y(n_1590)
);

NAND2x1p5_ASAP7_75t_L g1591 ( 
.A(n_1263),
.B(n_963),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1229),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1275),
.B(n_727),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1154),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1239),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1314),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1273),
.B(n_849),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1267),
.A2(n_728),
.B1(n_736),
.B2(n_730),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1320),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1320),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1320),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1320),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1270),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1280),
.B(n_870),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1270),
.B(n_730),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1286),
.B(n_877),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1288),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1291),
.B(n_887),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1292),
.Y(n_1609)
);

XNOR2x2_ASAP7_75t_L g1610 ( 
.A(n_1169),
.B(n_777),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1295),
.B(n_894),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1299),
.B(n_906),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1300),
.B(n_913),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1366),
.B(n_738),
.Y(n_1614)
);

OR2x6_ASAP7_75t_L g1615 ( 
.A(n_1460),
.B(n_1270),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1341),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1382),
.B(n_1166),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1364),
.A2(n_694),
.B1(n_741),
.B2(n_736),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1423),
.B(n_922),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1423),
.A2(n_1313),
.B1(n_1319),
.B2(n_1315),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1465),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1366),
.B(n_1392),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1424),
.B(n_1452),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1424),
.B(n_932),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1341),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1364),
.A2(n_743),
.B1(n_747),
.B2(n_741),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1336),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1392),
.B(n_740),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1458),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1454),
.B(n_1178),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1391),
.B(n_1404),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1391),
.B(n_938),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1493),
.B(n_1182),
.Y(n_1633)
);

NAND2x1p5_ASAP7_75t_L g1634 ( 
.A(n_1402),
.B(n_743),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1404),
.B(n_946),
.Y(n_1635)
);

NAND2x1p5_ASAP7_75t_L g1636 ( 
.A(n_1402),
.B(n_747),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1451),
.A2(n_1390),
.B1(n_1395),
.B2(n_1441),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1447),
.B(n_744),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1411),
.B(n_948),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1458),
.A2(n_1322),
.B1(n_1323),
.B2(n_1321),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1364),
.A2(n_757),
.B1(n_759),
.B2(n_752),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1411),
.B(n_953),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1447),
.B(n_745),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1493),
.B(n_1186),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1415),
.B(n_956),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1432),
.B(n_1241),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1336),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1462),
.B(n_746),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1370),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1415),
.B(n_1190),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1462),
.B(n_1394),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1484),
.B(n_959),
.Y(n_1652)
);

INVx8_ASAP7_75t_L g1653 ( 
.A(n_1335),
.Y(n_1653)
);

AND2x6_ASAP7_75t_SL g1654 ( 
.A(n_1460),
.B(n_1235),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1335),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1465),
.B(n_1477),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1432),
.B(n_1328),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1542),
.B(n_1199),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1538),
.B(n_749),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1488),
.B(n_960),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1338),
.B(n_961),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1340),
.B(n_1200),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1475),
.A2(n_753),
.B1(n_755),
.B2(n_754),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1513),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1416),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1353),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1542),
.B(n_1277),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1420),
.B(n_962),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1538),
.B(n_760),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1513),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1475),
.A2(n_765),
.B1(n_770),
.B2(n_763),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1527),
.Y(n_1672)
);

NAND3xp33_ASAP7_75t_SL g1673 ( 
.A(n_1511),
.B(n_1209),
.C(n_1245),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1333),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1397),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1439),
.Y(n_1676)
);

O2A1O1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1598),
.A2(n_1531),
.B(n_1375),
.C(n_1380),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1398),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1479),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1335),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1528),
.B(n_1431),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1528),
.B(n_773),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1336),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1407),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1453),
.B(n_987),
.Y(n_1685)
);

AND2x6_ASAP7_75t_L g1686 ( 
.A(n_1381),
.B(n_752),
.Y(n_1686)
);

AND2x6_ASAP7_75t_SL g1687 ( 
.A(n_1460),
.B(n_1244),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1334),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1413),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1470),
.B(n_1277),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1533),
.A2(n_759),
.B1(n_761),
.B2(n_757),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1533),
.B(n_965),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1418),
.B(n_774),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1455),
.B(n_1277),
.Y(n_1694)
);

INVx2_ASAP7_75t_SL g1695 ( 
.A(n_1579),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1422),
.B(n_776),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1425),
.B(n_780),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1579),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1556),
.B(n_967),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1448),
.B(n_786),
.Y(n_1700)
);

AO22x1_ASAP7_75t_L g1701 ( 
.A1(n_1417),
.A2(n_1403),
.B1(n_1594),
.B2(n_1583),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1464),
.B(n_790),
.Y(n_1702)
);

BUFx8_ASAP7_75t_L g1703 ( 
.A(n_1457),
.Y(n_1703)
);

A2O1A1Ixp33_ASAP7_75t_SL g1704 ( 
.A1(n_1347),
.A2(n_762),
.B(n_766),
.C(n_761),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1337),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1471),
.B(n_793),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1473),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1468),
.Y(n_1708)
);

NOR3x1_ASAP7_75t_L g1709 ( 
.A(n_1571),
.B(n_1283),
.C(n_1249),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1501),
.B(n_1277),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1431),
.B(n_794),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1509),
.A2(n_766),
.B1(n_781),
.B2(n_762),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1598),
.A2(n_783),
.B(n_784),
.C(n_781),
.Y(n_1713)
);

AND2x6_ASAP7_75t_L g1714 ( 
.A(n_1381),
.B(n_783),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1409),
.B(n_972),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1355),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1475),
.A2(n_798),
.B1(n_800),
.B2(n_799),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1427),
.B(n_1268),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1603),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1354),
.B(n_802),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1509),
.B(n_805),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1349),
.A2(n_789),
.B(n_784),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1509),
.B(n_807),
.Y(n_1723)
);

NOR3x1_ASAP7_75t_L g1724 ( 
.A(n_1576),
.B(n_1330),
.C(n_801),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1509),
.B(n_808),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1386),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1475),
.A2(n_801),
.B1(n_812),
.B2(n_789),
.Y(n_1727)
);

NOR3xp33_ASAP7_75t_L g1728 ( 
.A(n_1586),
.B(n_795),
.C(n_810),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1363),
.A2(n_815),
.B1(n_818),
.B2(n_811),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1363),
.B(n_822),
.Y(n_1730)
);

INVxp67_ASAP7_75t_L g1731 ( 
.A(n_1399),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1502),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1483),
.A2(n_817),
.B1(n_829),
.B2(n_812),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1450),
.B(n_826),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1414),
.B(n_827),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1414),
.B(n_830),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1345),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1375),
.A2(n_829),
.B1(n_832),
.B2(n_817),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1376),
.B(n_834),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1346),
.Y(n_1740)
);

A2O1A1Ixp33_ASAP7_75t_L g1741 ( 
.A1(n_1405),
.A2(n_838),
.B(n_839),
.C(n_832),
.Y(n_1741)
);

O2A1O1Ixp5_ASAP7_75t_L g1742 ( 
.A1(n_1376),
.A2(n_839),
.B(n_841),
.C(n_838),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1403),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1503),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1468),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1515),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1483),
.A2(n_844),
.B1(n_846),
.B2(n_841),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1519),
.B(n_1352),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1521),
.B(n_835),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1380),
.B(n_840),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1524),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1348),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1562),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1535),
.Y(n_1754)
);

A2O1A1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1405),
.A2(n_846),
.B(n_847),
.C(n_844),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1350),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1443),
.B(n_842),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1539),
.B(n_843),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1388),
.B(n_845),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1438),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1388),
.B(n_854),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1357),
.B(n_855),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1419),
.B(n_857),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1367),
.B(n_858),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1521),
.B(n_862),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_1582),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1481),
.Y(n_1767)
);

NAND2x1p5_ASAP7_75t_L g1768 ( 
.A(n_1500),
.B(n_847),
.Y(n_1768)
);

BUFx12f_ASAP7_75t_L g1769 ( 
.A(n_1438),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1480),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1419),
.B(n_864),
.Y(n_1771)
);

NOR3xp33_ASAP7_75t_L g1772 ( 
.A(n_1343),
.B(n_868),
.C(n_867),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1435),
.B(n_869),
.Y(n_1773)
);

AND2x6_ASAP7_75t_L g1774 ( 
.A(n_1385),
.B(n_856),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1435),
.B(n_871),
.Y(n_1775)
);

OAI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1505),
.A2(n_1522),
.B1(n_1594),
.B2(n_1583),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1435),
.B(n_873),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1360),
.Y(n_1778)
);

INVx2_ASAP7_75t_SL g1779 ( 
.A(n_1476),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1355),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1482),
.Y(n_1781)
);

O2A1O1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1385),
.A2(n_861),
.B(n_872),
.C(n_859),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1387),
.B(n_1445),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1476),
.Y(n_1784)
);

NOR2x1p5_ASAP7_75t_L g1785 ( 
.A(n_1491),
.B(n_954),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1435),
.B(n_875),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1514),
.B(n_878),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1514),
.B(n_879),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_SL g1789 ( 
.A1(n_1543),
.A2(n_885),
.B1(n_888),
.B2(n_884),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1591),
.Y(n_1790)
);

O2A1O1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1406),
.A2(n_1412),
.B(n_1510),
.C(n_1490),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1442),
.B(n_889),
.Y(n_1792)
);

XOR2xp5_ASAP7_75t_L g1793 ( 
.A(n_1536),
.B(n_891),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1442),
.A2(n_876),
.B1(n_890),
.B2(n_872),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1377),
.A2(n_1412),
.B1(n_1406),
.B2(n_1359),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1362),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1516),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1446),
.B(n_893),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1377),
.B(n_895),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1605),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1478),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1463),
.B(n_897),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1355),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1442),
.B(n_898),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1505),
.B(n_1492),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1339),
.A2(n_890),
.B1(n_892),
.B2(n_876),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1518),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_SL g1808 ( 
.A1(n_1522),
.A2(n_899),
.B1(n_902),
.B2(n_901),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1396),
.B(n_904),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1408),
.B(n_908),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1540),
.A2(n_907),
.B(n_892),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1541),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1605),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1374),
.Y(n_1814)
);

BUFx6f_ASAP7_75t_L g1815 ( 
.A(n_1365),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1591),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1442),
.B(n_910),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1378),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_SL g1819 ( 
.A(n_1592),
.B(n_971),
.C(n_912),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1529),
.B(n_911),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1444),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1512),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1499),
.B(n_914),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1529),
.B(n_915),
.Y(n_1824)
);

NAND2x1p5_ASAP7_75t_L g1825 ( 
.A(n_1603),
.B(n_907),
.Y(n_1825)
);

NOR3x1_ASAP7_75t_L g1826 ( 
.A(n_1494),
.B(n_921),
.C(n_920),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1512),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1551),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1365),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1486),
.B(n_1489),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1486),
.B(n_916),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1489),
.B(n_917),
.Y(n_1832)
);

OAI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1587),
.A2(n_924),
.B1(n_926),
.B2(n_923),
.C(n_918),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1540),
.B(n_928),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1498),
.B(n_930),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1498),
.B(n_931),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1505),
.A2(n_935),
.B1(n_936),
.B2(n_933),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1430),
.A2(n_940),
.B1(n_941),
.B2(n_939),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1506),
.B(n_1507),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1430),
.A2(n_1351),
.B1(n_1347),
.B2(n_1570),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1467),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1365),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1506),
.B(n_942),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1507),
.B(n_943),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1339),
.B(n_1359),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1587),
.A2(n_921),
.B1(n_934),
.B2(n_920),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1526),
.B(n_945),
.Y(n_1847)
);

A2O1A1Ixp33_ASAP7_75t_SL g1848 ( 
.A1(n_1351),
.A2(n_951),
.B(n_955),
.C(n_934),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1461),
.B(n_947),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1461),
.B(n_950),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1461),
.B(n_952),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1430),
.A2(n_958),
.B1(n_964),
.B2(n_957),
.Y(n_1852)
);

BUFx3_ASAP7_75t_L g1853 ( 
.A(n_1603),
.Y(n_1853)
);

A2O1A1Ixp33_ASAP7_75t_L g1854 ( 
.A1(n_1449),
.A2(n_955),
.B(n_963),
.C(n_951),
.Y(n_1854)
);

NAND2xp33_ASAP7_75t_L g1855 ( 
.A(n_1532),
.B(n_969),
.Y(n_1855)
);

NAND2xp33_ASAP7_75t_L g1856 ( 
.A(n_1532),
.B(n_614),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1430),
.A2(n_976),
.B1(n_980),
.B2(n_970),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1593),
.Y(n_1858)
);

NAND2xp33_ASAP7_75t_SL g1859 ( 
.A(n_1537),
.B(n_1544),
.Y(n_1859)
);

NAND2xp33_ASAP7_75t_L g1860 ( 
.A(n_1532),
.B(n_1428),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1577),
.B(n_970),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1570),
.A2(n_980),
.B1(n_981),
.B2(n_976),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1504),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1595),
.B(n_986),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1508),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1461),
.B(n_986),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1490),
.B(n_990),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1371),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1495),
.B(n_614),
.Y(n_1869)
);

AO22x1_ASAP7_75t_L g1870 ( 
.A1(n_1554),
.A2(n_644),
.B1(n_659),
.B2(n_614),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1589),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1371),
.Y(n_1872)
);

O2A1O1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1510),
.A2(n_644),
.B(n_659),
.C(n_614),
.Y(n_1873)
);

OR2x6_ASAP7_75t_L g1874 ( 
.A(n_1358),
.B(n_865),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1449),
.A2(n_1574),
.B1(n_1466),
.B2(n_1517),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1496),
.A2(n_1428),
.B1(n_1520),
.B2(n_1352),
.Y(n_1876)
);

AND2x6_ASAP7_75t_SL g1877 ( 
.A(n_1607),
.B(n_8),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1428),
.B(n_644),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1428),
.B(n_644),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1466),
.B(n_1384),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1384),
.B(n_1426),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1495),
.B(n_644),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1371),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1426),
.B(n_659),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1523),
.B(n_659),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1530),
.B(n_659),
.Y(n_1886)
);

NAND2xp33_ASAP7_75t_L g1887 ( 
.A(n_1532),
.B(n_722),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1545),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1580),
.A2(n_772),
.B1(n_791),
.B2(n_722),
.Y(n_1889)
);

A2O1A1Ixp33_ASAP7_75t_SL g1890 ( 
.A1(n_1534),
.A2(n_772),
.B(n_791),
.C(n_722),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1554),
.Y(n_1891)
);

NAND2x1p5_ASAP7_75t_L g1892 ( 
.A(n_1379),
.B(n_1434),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1373),
.Y(n_1893)
);

A2O1A1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1552),
.A2(n_772),
.B(n_791),
.C(n_722),
.Y(n_1894)
);

BUFx6f_ASAP7_75t_L g1895 ( 
.A(n_1373),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1520),
.B(n_722),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1496),
.A2(n_791),
.B1(n_865),
.B2(n_772),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1373),
.Y(n_1898)
);

AO22x1_ASAP7_75t_L g1899 ( 
.A1(n_1554),
.A2(n_791),
.B1(n_865),
.B2(n_772),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1593),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1604),
.B(n_8),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1568),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1580),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1393),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1520),
.A2(n_1552),
.B1(n_1588),
.B2(n_1561),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1612),
.B(n_865),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1520),
.B(n_865),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1561),
.A2(n_16),
.B1(n_9),
.B2(n_15),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1517),
.A2(n_17),
.B1(n_9),
.B2(n_15),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1588),
.B(n_18),
.Y(n_1910)
);

BUFx2_ASAP7_75t_L g1911 ( 
.A(n_1610),
.Y(n_1911)
);

INVxp67_ASAP7_75t_L g1912 ( 
.A(n_1612),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1604),
.B(n_18),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1597),
.B(n_19),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1546),
.B(n_20),
.Y(n_1915)
);

NOR2xp67_ASAP7_75t_L g1916 ( 
.A(n_1609),
.B(n_21),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1597),
.B(n_22),
.Y(n_1917)
);

AND2x6_ASAP7_75t_SL g1918 ( 
.A(n_1608),
.B(n_22),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_SL g1919 ( 
.A(n_1608),
.B(n_23),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1555),
.A2(n_446),
.B(n_442),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1565),
.B(n_24),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1611),
.B(n_25),
.Y(n_1922)
);

AOI22xp33_ASAP7_75t_L g1923 ( 
.A1(n_1356),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1546),
.B(n_29),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1497),
.B(n_30),
.Y(n_1925)
);

CKINVDCx20_ASAP7_75t_R g1926 ( 
.A(n_1611),
.Y(n_1926)
);

O2A1O1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1436),
.A2(n_33),
.B(n_30),
.C(n_32),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1525),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1393),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1393),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1649),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1622),
.B(n_1559),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1655),
.B(n_1606),
.Y(n_1933)
);

INVx1_ASAP7_75t_SL g1934 ( 
.A(n_1766),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1622),
.B(n_1613),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1825),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1675),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1678),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1684),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1825),
.Y(n_1940)
);

O2A1O1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1677),
.A2(n_1555),
.B(n_1361),
.C(n_1564),
.Y(n_1941)
);

BUFx3_ASAP7_75t_L g1942 ( 
.A(n_1769),
.Y(n_1942)
);

NAND3xp33_ASAP7_75t_SL g1943 ( 
.A(n_1905),
.B(n_1584),
.C(n_1564),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1689),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1628),
.B(n_1379),
.Y(n_1945)
);

BUFx2_ASAP7_75t_L g1946 ( 
.A(n_1653),
.Y(n_1946)
);

HB1xp67_ASAP7_75t_L g1947 ( 
.A(n_1653),
.Y(n_1947)
);

INVx5_ASAP7_75t_L g1948 ( 
.A(n_1653),
.Y(n_1948)
);

BUFx2_ASAP7_75t_L g1949 ( 
.A(n_1655),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1892),
.Y(n_1950)
);

NOR2xp67_ASAP7_75t_L g1951 ( 
.A(n_1673),
.B(n_35),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1707),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1731),
.B(n_1584),
.Y(n_1953)
);

INVx5_ASAP7_75t_L g1954 ( 
.A(n_1627),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1743),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1703),
.Y(n_1956)
);

OR2x6_ASAP7_75t_L g1957 ( 
.A(n_1701),
.B(n_1680),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1815),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_R g1959 ( 
.A(n_1666),
.B(n_1434),
.Y(n_1959)
);

INVx3_ASAP7_75t_L g1960 ( 
.A(n_1892),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1815),
.Y(n_1961)
);

BUFx6f_ASAP7_75t_L g1962 ( 
.A(n_1829),
.Y(n_1962)
);

OR2x4_ASAP7_75t_L g1963 ( 
.A(n_1633),
.B(n_1590),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1732),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1726),
.B(n_1437),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1753),
.B(n_1437),
.Y(n_1966)
);

INVxp67_ASAP7_75t_SL g1967 ( 
.A(n_1681),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1646),
.B(n_1590),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1845),
.B(n_1434),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_1665),
.Y(n_1970)
);

BUFx3_ASAP7_75t_L g1971 ( 
.A(n_1703),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1744),
.Y(n_1972)
);

INVx4_ASAP7_75t_L g1973 ( 
.A(n_1679),
.Y(n_1973)
);

INVx3_ASAP7_75t_L g1974 ( 
.A(n_1621),
.Y(n_1974)
);

NOR3xp33_ASAP7_75t_SL g1975 ( 
.A(n_1776),
.B(n_1558),
.C(n_1547),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1746),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1654),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1829),
.B(n_1883),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1657),
.B(n_1369),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1687),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1767),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1845),
.B(n_1369),
.Y(n_1982)
);

CKINVDCx14_ASAP7_75t_R g1983 ( 
.A(n_1837),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1637),
.B(n_1372),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1623),
.A2(n_1926),
.B1(n_1718),
.B2(n_1617),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1751),
.Y(n_1986)
);

BUFx4f_ASAP7_75t_L g1987 ( 
.A(n_1615),
.Y(n_1987)
);

NAND3xp33_ASAP7_75t_SL g1988 ( 
.A(n_1911),
.B(n_1344),
.C(n_1342),
.Y(n_1988)
);

NOR3xp33_ASAP7_75t_SL g1989 ( 
.A(n_1819),
.B(n_1566),
.C(n_1560),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1676),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1614),
.B(n_1372),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1754),
.Y(n_1992)
);

NAND3xp33_ASAP7_75t_SL g1993 ( 
.A(n_1927),
.B(n_1472),
.C(n_1469),
.Y(n_1993)
);

A2O1A1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1791),
.A2(n_1433),
.B(n_1456),
.C(n_1429),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1634),
.Y(n_1995)
);

AND2x4_ASAP7_75t_L g1996 ( 
.A(n_1822),
.B(n_1437),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1634),
.Y(n_1997)
);

NAND2x2_ASAP7_75t_L g1998 ( 
.A(n_1785),
.B(n_1760),
.Y(n_1998)
);

INVxp67_ASAP7_75t_SL g1999 ( 
.A(n_1790),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1674),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1830),
.B(n_1433),
.Y(n_2001)
);

NAND2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1876),
.B(n_1421),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1830),
.B(n_1456),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_R g2004 ( 
.A(n_1860),
.B(n_36),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1881),
.B(n_1474),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1839),
.B(n_1485),
.Y(n_2006)
);

OR2x2_ASAP7_75t_L g2007 ( 
.A(n_1620),
.B(n_37),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1903),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1789),
.Y(n_2009)
);

NOR3xp33_ASAP7_75t_SL g2010 ( 
.A(n_1859),
.B(n_1578),
.C(n_1572),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1829),
.Y(n_2011)
);

INVxp67_ASAP7_75t_L g2012 ( 
.A(n_1631),
.Y(n_2012)
);

A2O1A1Ixp33_ASAP7_75t_L g2013 ( 
.A1(n_1839),
.A2(n_1487),
.B(n_1383),
.C(n_1400),
.Y(n_2013)
);

AOI22xp33_ASAP7_75t_L g2014 ( 
.A1(n_1875),
.A2(n_1440),
.B1(n_1459),
.B2(n_1389),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1900),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1688),
.Y(n_2016)
);

BUFx3_ASAP7_75t_L g2017 ( 
.A(n_1779),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_1827),
.B(n_1459),
.Y(n_2018)
);

BUFx2_ASAP7_75t_L g2019 ( 
.A(n_1636),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1705),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1737),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1757),
.B(n_1368),
.Y(n_2022)
);

AND2x4_ASAP7_75t_L g2023 ( 
.A(n_1784),
.B(n_1368),
.Y(n_2023)
);

AOI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1644),
.A2(n_1440),
.B1(n_1401),
.B2(n_1410),
.Y(n_2024)
);

INVx3_ASAP7_75t_L g2025 ( 
.A(n_1621),
.Y(n_2025)
);

BUFx6f_ASAP7_75t_L g2026 ( 
.A(n_1883),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1770),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_R g2028 ( 
.A(n_1856),
.B(n_37),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1880),
.B(n_1440),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1781),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1748),
.Y(n_2031)
);

BUFx10_ASAP7_75t_L g2032 ( 
.A(n_1615),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1636),
.Y(n_2033)
);

INVx5_ASAP7_75t_L g2034 ( 
.A(n_1627),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1880),
.B(n_1368),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1748),
.B(n_1563),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1691),
.B(n_38),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1881),
.B(n_1861),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1888),
.Y(n_2039)
);

INVx4_ASAP7_75t_L g2040 ( 
.A(n_1615),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1866),
.Y(n_2041)
);

NOR2x1p5_ASAP7_75t_L g2042 ( 
.A(n_1805),
.B(n_39),
.Y(n_2042)
);

OR2x2_ASAP7_75t_SL g2043 ( 
.A(n_1864),
.B(n_40),
.Y(n_2043)
);

INVx3_ASAP7_75t_L g2044 ( 
.A(n_1708),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1858),
.B(n_40),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1740),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1795),
.A2(n_1557),
.B1(n_1563),
.B2(n_1548),
.Y(n_2047)
);

BUFx3_ASAP7_75t_L g2048 ( 
.A(n_1768),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1871),
.A2(n_1550),
.B1(n_1575),
.B2(n_1569),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_1656),
.B(n_1563),
.Y(n_2050)
);

NOR3xp33_ASAP7_75t_SL g2051 ( 
.A(n_1902),
.B(n_1599),
.C(n_1581),
.Y(n_2051)
);

A2O1A1Ixp33_ASAP7_75t_L g2052 ( 
.A1(n_1651),
.A2(n_1550),
.B(n_1575),
.C(n_1569),
.Y(n_2052)
);

INVx6_ASAP7_75t_L g2053 ( 
.A(n_1719),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1752),
.Y(n_2054)
);

AND2x4_ASAP7_75t_L g2055 ( 
.A(n_1912),
.B(n_1563),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1651),
.B(n_42),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_R g2057 ( 
.A(n_1887),
.B(n_43),
.Y(n_2057)
);

INVx3_ASAP7_75t_L g2058 ( 
.A(n_1708),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1866),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1756),
.Y(n_2060)
);

NAND2xp33_ASAP7_75t_R g2061 ( 
.A(n_1891),
.B(n_45),
.Y(n_2061)
);

BUFx6f_ASAP7_75t_L g2062 ( 
.A(n_1883),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1778),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1895),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1796),
.Y(n_2065)
);

CKINVDCx11_ASAP7_75t_R g2066 ( 
.A(n_1874),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1694),
.B(n_46),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1640),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_1840),
.B(n_1693),
.Y(n_2069)
);

AND2x6_ASAP7_75t_L g2070 ( 
.A(n_1816),
.B(n_1585),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1854),
.B(n_46),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1693),
.B(n_48),
.Y(n_2072)
);

BUFx3_ASAP7_75t_L g2073 ( 
.A(n_1768),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1710),
.B(n_48),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1800),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_1658),
.B(n_1585),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1638),
.B(n_49),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1638),
.B(n_50),
.Y(n_2078)
);

INVx4_ASAP7_75t_L g2079 ( 
.A(n_1874),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1797),
.Y(n_2080)
);

OAI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_1919),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_2081)
);

NOR3xp33_ASAP7_75t_SL g2082 ( 
.A(n_1650),
.B(n_1602),
.C(n_1600),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_1745),
.Y(n_2083)
);

INVx1_ASAP7_75t_SL g2084 ( 
.A(n_1793),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1643),
.B(n_52),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1895),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1826),
.B(n_53),
.Y(n_2087)
);

BUFx6f_ASAP7_75t_L g2088 ( 
.A(n_1895),
.Y(n_2088)
);

INVxp67_ASAP7_75t_L g2089 ( 
.A(n_1686),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_1667),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_R g2091 ( 
.A(n_1855),
.B(n_54),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_R g2092 ( 
.A(n_1695),
.B(n_55),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1627),
.B(n_1549),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1807),
.Y(n_2094)
);

INVxp67_ASAP7_75t_L g2095 ( 
.A(n_1686),
.Y(n_2095)
);

AND2x6_ASAP7_75t_L g2096 ( 
.A(n_1629),
.B(n_1549),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_1922),
.B(n_55),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1647),
.B(n_1549),
.Y(n_2098)
);

OR2x2_ASAP7_75t_SL g2099 ( 
.A(n_1709),
.B(n_57),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_R g2100 ( 
.A(n_1698),
.B(n_57),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1643),
.B(n_58),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1648),
.B(n_58),
.Y(n_2102)
);

HB1xp67_ASAP7_75t_L g2103 ( 
.A(n_1686),
.Y(n_2103)
);

AOI21x1_ASAP7_75t_L g2104 ( 
.A1(n_1896),
.A2(n_1596),
.B(n_1573),
.Y(n_2104)
);

INVx1_ASAP7_75t_SL g2105 ( 
.A(n_1828),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1812),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1749),
.B(n_60),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1765),
.B(n_61),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1813),
.Y(n_2109)
);

NAND3xp33_ASAP7_75t_SL g2110 ( 
.A(n_1908),
.B(n_1601),
.C(n_63),
.Y(n_2110)
);

BUFx8_ASAP7_75t_L g2111 ( 
.A(n_1906),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_1730),
.B(n_63),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_1735),
.B(n_64),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_1736),
.B(n_65),
.Y(n_2114)
);

BUFx2_ASAP7_75t_L g2115 ( 
.A(n_1874),
.Y(n_2115)
);

BUFx6f_ASAP7_75t_L g2116 ( 
.A(n_1647),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1867),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1814),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1818),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1867),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1647),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1821),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1696),
.B(n_65),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1696),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1683),
.B(n_1553),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1841),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_1877),
.Y(n_2127)
);

BUFx6f_ASAP7_75t_L g2128 ( 
.A(n_1683),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1683),
.B(n_1780),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_1686),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_R g2131 ( 
.A(n_1853),
.B(n_66),
.Y(n_2131)
);

AOI22xp5_ASAP7_75t_SL g2132 ( 
.A1(n_1630),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_2132)
);

NOR2xp33_ASAP7_75t_L g2133 ( 
.A(n_1697),
.B(n_68),
.Y(n_2133)
);

BUFx6f_ASAP7_75t_L g2134 ( 
.A(n_1716),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1716),
.B(n_1553),
.Y(n_2135)
);

AND2x4_ASAP7_75t_SL g2136 ( 
.A(n_1728),
.B(n_1663),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_1745),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1918),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_SL g2139 ( 
.A(n_1716),
.B(n_1567),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1780),
.B(n_1567),
.Y(n_2140)
);

INVx2_ASAP7_75t_SL g2141 ( 
.A(n_1661),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1697),
.B(n_69),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1700),
.B(n_69),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1700),
.B(n_70),
.Y(n_2144)
);

OAI22xp33_ASAP7_75t_L g2145 ( 
.A1(n_1928),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1702),
.B(n_72),
.Y(n_2146)
);

NOR2xp67_ASAP7_75t_L g2147 ( 
.A(n_1729),
.B(n_1833),
.Y(n_2147)
);

INVx5_ASAP7_75t_L g2148 ( 
.A(n_1780),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_1808),
.Y(n_2149)
);

NOR3xp33_ASAP7_75t_SL g2150 ( 
.A(n_1909),
.B(n_73),
.C(n_74),
.Y(n_2150)
);

BUFx6f_ASAP7_75t_L g2151 ( 
.A(n_1803),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_1801),
.Y(n_2152)
);

BUFx12f_ASAP7_75t_SL g2153 ( 
.A(n_1724),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1863),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1702),
.Y(n_2155)
);

INVx3_ASAP7_75t_L g2156 ( 
.A(n_1664),
.Y(n_2156)
);

INVx5_ASAP7_75t_L g2157 ( 
.A(n_1803),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1706),
.B(n_75),
.Y(n_2158)
);

INVx8_ASAP7_75t_L g2159 ( 
.A(n_1714),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1706),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_R g2161 ( 
.A(n_1714),
.B(n_75),
.Y(n_2161)
);

NOR2xp33_ASAP7_75t_L g2162 ( 
.A(n_1692),
.B(n_76),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_1787),
.B(n_77),
.Y(n_2163)
);

INVx3_ASAP7_75t_L g2164 ( 
.A(n_1664),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_1788),
.B(n_79),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1865),
.Y(n_2166)
);

BUFx4f_ASAP7_75t_SL g2167 ( 
.A(n_1869),
.Y(n_2167)
);

INVx3_ASAP7_75t_L g2168 ( 
.A(n_1616),
.Y(n_2168)
);

INVx6_ASAP7_75t_L g2169 ( 
.A(n_1714),
.Y(n_2169)
);

NAND3xp33_ASAP7_75t_SL g2170 ( 
.A(n_1618),
.B(n_79),
.C(n_80),
.Y(n_2170)
);

BUFx2_ASAP7_75t_L g2171 ( 
.A(n_1714),
.Y(n_2171)
);

BUFx3_ASAP7_75t_L g2172 ( 
.A(n_1774),
.Y(n_2172)
);

BUFx12f_ASAP7_75t_L g2173 ( 
.A(n_1774),
.Y(n_2173)
);

NOR3xp33_ASAP7_75t_SL g2174 ( 
.A(n_1901),
.B(n_80),
.C(n_81),
.Y(n_2174)
);

NOR3xp33_ASAP7_75t_SL g2175 ( 
.A(n_1913),
.B(n_81),
.C(n_83),
.Y(n_2175)
);

BUFx3_ASAP7_75t_L g2176 ( 
.A(n_1774),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1823),
.B(n_84),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1670),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1672),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1711),
.Y(n_2180)
);

OR2x2_ASAP7_75t_L g2181 ( 
.A(n_1659),
.B(n_84),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1758),
.Y(n_2182)
);

INVx5_ASAP7_75t_L g2183 ( 
.A(n_1774),
.Y(n_2183)
);

AND2x4_ASAP7_75t_SL g2184 ( 
.A(n_1671),
.B(n_85),
.Y(n_2184)
);

INVx2_ASAP7_75t_SL g2185 ( 
.A(n_1668),
.Y(n_2185)
);

INVx3_ASAP7_75t_L g2186 ( 
.A(n_1625),
.Y(n_2186)
);

AND3x1_ASAP7_75t_L g2187 ( 
.A(n_1662),
.B(n_86),
.C(n_87),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1925),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_1847),
.B(n_87),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_1820),
.B(n_89),
.Y(n_2190)
);

AOI22xp33_ASAP7_75t_SL g2191 ( 
.A1(n_1774),
.A2(n_93),
.B1(n_90),
.B2(n_92),
.Y(n_2191)
);

AND2x4_ASAP7_75t_L g2192 ( 
.A(n_1824),
.B(n_90),
.Y(n_2192)
);

INVx4_ASAP7_75t_L g2193 ( 
.A(n_1930),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1925),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1733),
.B(n_93),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1747),
.B(n_94),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1862),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_1690),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1842),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1742),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1626),
.B(n_1548),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_1759),
.B(n_95),
.Y(n_2202)
);

NOR3xp33_ASAP7_75t_SL g2203 ( 
.A(n_1734),
.B(n_95),
.C(n_96),
.Y(n_2203)
);

INVx2_ASAP7_75t_SL g2204 ( 
.A(n_1619),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1739),
.B(n_96),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1717),
.Y(n_2206)
);

INVx1_ASAP7_75t_SL g2207 ( 
.A(n_1849),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1641),
.B(n_97),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_1761),
.B(n_97),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_1750),
.B(n_98),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1831),
.B(n_1832),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1889),
.Y(n_2212)
);

INVx3_ASAP7_75t_L g2213 ( 
.A(n_1868),
.Y(n_2213)
);

NOR2x1_ASAP7_75t_L g2214 ( 
.A(n_1699),
.B(n_98),
.Y(n_2214)
);

AND2x6_ASAP7_75t_L g2215 ( 
.A(n_1896),
.B(n_447),
.Y(n_2215)
);

INVx3_ASAP7_75t_L g2216 ( 
.A(n_1872),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_1763),
.B(n_1771),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1669),
.B(n_99),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1907),
.Y(n_2219)
);

NOR3xp33_ASAP7_75t_SL g2220 ( 
.A(n_1741),
.B(n_102),
.C(n_103),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1907),
.Y(n_2221)
);

INVx5_ASAP7_75t_L g2222 ( 
.A(n_1893),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_R g2223 ( 
.A(n_1727),
.B(n_102),
.Y(n_2223)
);

BUFx3_ASAP7_75t_L g2224 ( 
.A(n_1783),
.Y(n_2224)
);

INVx2_ASAP7_75t_SL g2225 ( 
.A(n_1624),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_1849),
.Y(n_2226)
);

HB1xp67_ASAP7_75t_L g2227 ( 
.A(n_1870),
.Y(n_2227)
);

BUFx2_ASAP7_75t_L g2228 ( 
.A(n_1804),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1898),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1915),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1924),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1904),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1806),
.Y(n_2233)
);

BUFx3_ASAP7_75t_L g2234 ( 
.A(n_1850),
.Y(n_2234)
);

BUFx10_ASAP7_75t_L g2235 ( 
.A(n_1809),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1682),
.Y(n_2236)
);

AOI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_1772),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_2237)
);

AND2x4_ASAP7_75t_L g2238 ( 
.A(n_1834),
.B(n_105),
.Y(n_2238)
);

NAND2x2_ASAP7_75t_L g2239 ( 
.A(n_1835),
.B(n_106),
.Y(n_2239)
);

BUFx3_ASAP7_75t_L g2240 ( 
.A(n_1850),
.Y(n_2240)
);

NOR3xp33_ASAP7_75t_SL g2241 ( 
.A(n_1755),
.B(n_108),
.C(n_109),
.Y(n_2241)
);

OR2x4_ASAP7_75t_L g2242 ( 
.A(n_1798),
.B(n_109),
.Y(n_2242)
);

NOR3xp33_ASAP7_75t_SL g2243 ( 
.A(n_1846),
.B(n_110),
.C(n_111),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1929),
.Y(n_2244)
);

A2O1A1Ixp33_ASAP7_75t_L g2245 ( 
.A1(n_1782),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1835),
.B(n_1836),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_R g2247 ( 
.A(n_1804),
.B(n_112),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1799),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1836),
.B(n_114),
.Y(n_2249)
);

BUFx8_ASAP7_75t_L g2250 ( 
.A(n_1916),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1799),
.Y(n_2251)
);

INVxp67_ASAP7_75t_SL g2252 ( 
.A(n_1899),
.Y(n_2252)
);

NAND2xp33_ASAP7_75t_R g2253 ( 
.A(n_1817),
.B(n_115),
.Y(n_2253)
);

INVx5_ASAP7_75t_L g2254 ( 
.A(n_1794),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1843),
.B(n_1844),
.Y(n_2255)
);

NOR3xp33_ASAP7_75t_SL g2256 ( 
.A(n_1738),
.B(n_117),
.C(n_118),
.Y(n_2256)
);

OAI22xp33_ASAP7_75t_L g2257 ( 
.A1(n_1910),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_2257)
);

HB1xp67_ASAP7_75t_L g2258 ( 
.A(n_1878),
.Y(n_2258)
);

HB1xp67_ASAP7_75t_L g2259 ( 
.A(n_1879),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1713),
.Y(n_2260)
);

AND2x4_ASAP7_75t_L g2261 ( 
.A(n_1660),
.B(n_119),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1910),
.Y(n_2262)
);

INVx2_ASAP7_75t_SL g2263 ( 
.A(n_1645),
.Y(n_2263)
);

BUFx3_ASAP7_75t_L g2264 ( 
.A(n_1851),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_L g2265 ( 
.A(n_1843),
.B(n_121),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_1844),
.B(n_122),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_1720),
.B(n_122),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_1879),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1715),
.B(n_123),
.Y(n_2269)
);

AO22x1_ASAP7_75t_L g2270 ( 
.A1(n_1817),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_2270)
);

NAND2xp33_ASAP7_75t_SL g2271 ( 
.A(n_1914),
.B(n_1917),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_1882),
.Y(n_2272)
);

NAND3xp33_ASAP7_75t_SL g2273 ( 
.A(n_1704),
.B(n_126),
.C(n_127),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1914),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_1712),
.B(n_128),
.Y(n_2275)
);

BUFx3_ASAP7_75t_L g2276 ( 
.A(n_1851),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1722),
.B(n_129),
.Y(n_2277)
);

NAND3xp33_ASAP7_75t_L g2278 ( 
.A(n_1894),
.B(n_130),
.C(n_132),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1811),
.B(n_133),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1857),
.B(n_134),
.Y(n_2280)
);

BUFx3_ASAP7_75t_L g2281 ( 
.A(n_1810),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1635),
.B(n_1838),
.Y(n_2282)
);

INVx3_ASAP7_75t_L g2283 ( 
.A(n_1917),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_1852),
.B(n_134),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1884),
.Y(n_2285)
);

NOR3xp33_ASAP7_75t_SL g2286 ( 
.A(n_1685),
.B(n_135),
.C(n_136),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_1802),
.B(n_135),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_1920),
.B(n_450),
.Y(n_2288)
);

INVx5_ASAP7_75t_L g2289 ( 
.A(n_1848),
.Y(n_2289)
);

OAI21xp33_ASAP7_75t_L g2290 ( 
.A1(n_1921),
.A2(n_136),
.B(n_137),
.Y(n_2290)
);

NAND2xp33_ASAP7_75t_SL g2291 ( 
.A(n_1921),
.B(n_139),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1762),
.B(n_139),
.Y(n_2292)
);

OR2x6_ASAP7_75t_L g2293 ( 
.A(n_1652),
.B(n_140),
.Y(n_2293)
);

INVx5_ASAP7_75t_L g2294 ( 
.A(n_1897),
.Y(n_2294)
);

AOI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_1764),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_1721),
.B(n_141),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1723),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_R g2298 ( 
.A(n_1773),
.B(n_143),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1885),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_1775),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1725),
.Y(n_2301)
);

BUFx2_ASAP7_75t_L g2302 ( 
.A(n_1934),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2117),
.B(n_1777),
.Y(n_2303)
);

OAI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2246),
.A2(n_1886),
.B(n_1885),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2120),
.B(n_1786),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1952),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2048),
.B(n_1632),
.Y(n_2307)
);

INVx4_ASAP7_75t_L g2308 ( 
.A(n_1948),
.Y(n_2308)
);

OAI21x1_ASAP7_75t_L g2309 ( 
.A1(n_2104),
.A2(n_1886),
.B(n_1873),
.Y(n_2309)
);

OAI21xp5_ASAP7_75t_L g2310 ( 
.A1(n_2246),
.A2(n_2255),
.B(n_2211),
.Y(n_2310)
);

OAI21x1_ASAP7_75t_L g2311 ( 
.A1(n_1978),
.A2(n_1642),
.B(n_1639),
.Y(n_2311)
);

OAI21xp5_ASAP7_75t_L g2312 ( 
.A1(n_1941),
.A2(n_1923),
.B(n_1792),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2038),
.B(n_1890),
.Y(n_2313)
);

INVx3_ASAP7_75t_L g2314 ( 
.A(n_1950),
.Y(n_2314)
);

A2O1A1Ixp33_ASAP7_75t_L g2315 ( 
.A1(n_2069),
.A2(n_147),
.B(n_144),
.C(n_146),
.Y(n_2315)
);

OAI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_1941),
.A2(n_146),
.B(n_147),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1964),
.Y(n_2317)
);

OAI21x1_ASAP7_75t_L g2318 ( 
.A1(n_2129),
.A2(n_453),
.B(n_452),
.Y(n_2318)
);

NAND2x1p5_ASAP7_75t_L g2319 ( 
.A(n_1948),
.B(n_148),
.Y(n_2319)
);

OAI21x1_ASAP7_75t_L g2320 ( 
.A1(n_2129),
.A2(n_455),
.B(n_454),
.Y(n_2320)
);

AOI21xp5_ASAP7_75t_L g2321 ( 
.A1(n_2271),
.A2(n_458),
.B(n_456),
.Y(n_2321)
);

AOI31xp67_ASAP7_75t_L g2322 ( 
.A1(n_2288),
.A2(n_598),
.A3(n_460),
.B(n_461),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2069),
.B(n_2260),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2248),
.B(n_149),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2251),
.B(n_150),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2124),
.B(n_150),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_SL g2327 ( 
.A(n_1987),
.B(n_151),
.Y(n_2327)
);

OAI21x1_ASAP7_75t_L g2328 ( 
.A1(n_2093),
.A2(n_462),
.B(n_459),
.Y(n_2328)
);

NOR4xp25_ASAP7_75t_L g2329 ( 
.A(n_2170),
.B(n_154),
.C(n_151),
.D(n_152),
.Y(n_2329)
);

OAI21x1_ASAP7_75t_L g2330 ( 
.A1(n_2093),
.A2(n_2125),
.B(n_2098),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2073),
.B(n_1999),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_L g2332 ( 
.A(n_1985),
.B(n_152),
.Y(n_2332)
);

AOI221x1_ASAP7_75t_L g2333 ( 
.A1(n_2271),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.C(n_158),
.Y(n_2333)
);

AND2x4_ASAP7_75t_L g2334 ( 
.A(n_1948),
.B(n_155),
.Y(n_2334)
);

OAI21x1_ASAP7_75t_L g2335 ( 
.A1(n_2098),
.A2(n_465),
.B(n_464),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_1987),
.B(n_157),
.Y(n_2336)
);

NAND3xp33_ASAP7_75t_SL g2337 ( 
.A(n_2131),
.B(n_159),
.C(n_160),
.Y(n_2337)
);

A2O1A1Ixp33_ASAP7_75t_L g2338 ( 
.A1(n_2265),
.A2(n_2217),
.B(n_2072),
.C(n_2133),
.Y(n_2338)
);

OAI21x1_ASAP7_75t_L g2339 ( 
.A1(n_2125),
.A2(n_2139),
.B(n_2135),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2155),
.B(n_159),
.Y(n_2340)
);

INVxp67_ASAP7_75t_SL g2341 ( 
.A(n_1995),
.Y(n_2341)
);

HB1xp67_ASAP7_75t_L g2342 ( 
.A(n_1995),
.Y(n_2342)
);

AOI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_2013),
.A2(n_469),
.B(n_466),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2160),
.B(n_160),
.Y(n_2344)
);

CKINVDCx16_ASAP7_75t_R g2345 ( 
.A(n_1971),
.Y(n_2345)
);

OAI21x1_ASAP7_75t_L g2346 ( 
.A1(n_2135),
.A2(n_476),
.B(n_471),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_1999),
.B(n_161),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2233),
.B(n_161),
.Y(n_2348)
);

A2O1A1Ixp33_ASAP7_75t_L g2349 ( 
.A1(n_2265),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_2349)
);

BUFx3_ASAP7_75t_L g2350 ( 
.A(n_1942),
.Y(n_2350)
);

NAND2xp33_ASAP7_75t_L g2351 ( 
.A(n_2028),
.B(n_162),
.Y(n_2351)
);

AO21x2_ASAP7_75t_L g2352 ( 
.A1(n_1994),
.A2(n_480),
.B(n_477),
.Y(n_2352)
);

OAI21xp33_ASAP7_75t_L g2353 ( 
.A1(n_2223),
.A2(n_165),
.B(n_166),
.Y(n_2353)
);

BUFx2_ASAP7_75t_SL g2354 ( 
.A(n_1948),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_1950),
.Y(n_2355)
);

OAI21x1_ASAP7_75t_L g2356 ( 
.A1(n_2139),
.A2(n_482),
.B(n_481),
.Y(n_2356)
);

OAI21x1_ASAP7_75t_L g2357 ( 
.A1(n_2140),
.A2(n_486),
.B(n_484),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2197),
.B(n_165),
.Y(n_2358)
);

OAI21x1_ASAP7_75t_L g2359 ( 
.A1(n_2140),
.A2(n_490),
.B(n_488),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2091),
.B(n_166),
.Y(n_2360)
);

A2O1A1Ixp33_ASAP7_75t_L g2361 ( 
.A1(n_2217),
.A2(n_169),
.B(n_167),
.C(n_168),
.Y(n_2361)
);

BUFx2_ASAP7_75t_SL g2362 ( 
.A(n_1973),
.Y(n_2362)
);

NOR2x1_ASAP7_75t_R g2363 ( 
.A(n_1956),
.B(n_167),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2182),
.B(n_168),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2262),
.B(n_170),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2013),
.A2(n_1994),
.B(n_2288),
.Y(n_2366)
);

AOI21xp33_ASAP7_75t_L g2367 ( 
.A1(n_2274),
.A2(n_170),
.B(n_171),
.Y(n_2367)
);

NAND3xp33_ASAP7_75t_L g2368 ( 
.A(n_2174),
.B(n_172),
.C(n_173),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_1977),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1972),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2188),
.B(n_175),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_1976),
.Y(n_2372)
);

OA22x2_ASAP7_75t_L g2373 ( 
.A1(n_1957),
.A2(n_178),
.B1(n_175),
.B2(n_177),
.Y(n_2373)
);

OAI21xp5_ASAP7_75t_L g2374 ( 
.A1(n_1969),
.A2(n_177),
.B(n_178),
.Y(n_2374)
);

AOI21x1_ASAP7_75t_L g2375 ( 
.A1(n_2227),
.A2(n_499),
.B(n_498),
.Y(n_2375)
);

INVx3_ASAP7_75t_SL g2376 ( 
.A(n_1981),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2194),
.B(n_179),
.Y(n_2377)
);

OAI21x1_ASAP7_75t_L g2378 ( 
.A1(n_2047),
.A2(n_501),
.B(n_500),
.Y(n_2378)
);

NAND3xp33_ASAP7_75t_L g2379 ( 
.A(n_2174),
.B(n_180),
.C(n_181),
.Y(n_2379)
);

BUFx2_ASAP7_75t_L g2380 ( 
.A(n_2161),
.Y(n_2380)
);

AO31x2_ASAP7_75t_L g2381 ( 
.A1(n_2052),
.A2(n_2285),
.A3(n_2299),
.B(n_2200),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_SL g2382 ( 
.A1(n_2252),
.A2(n_510),
.B(n_508),
.Y(n_2382)
);

INVx3_ASAP7_75t_L g2383 ( 
.A(n_1960),
.Y(n_2383)
);

OAI21x1_ASAP7_75t_L g2384 ( 
.A1(n_2047),
.A2(n_513),
.B(n_511),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_1931),
.B(n_181),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_1943),
.A2(n_519),
.B(n_515),
.Y(n_2386)
);

O2A1O1Ixp5_ASAP7_75t_L g2387 ( 
.A1(n_2002),
.A2(n_523),
.B(n_524),
.C(n_522),
.Y(n_2387)
);

AOI21x1_ASAP7_75t_L g2388 ( 
.A1(n_2227),
.A2(n_535),
.B(n_526),
.Y(n_2388)
);

AOI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_1943),
.A2(n_538),
.B(n_536),
.Y(n_2389)
);

HB1xp67_ASAP7_75t_L g2390 ( 
.A(n_1997),
.Y(n_2390)
);

AOI22xp5_ASAP7_75t_L g2391 ( 
.A1(n_2147),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_L g2392 ( 
.A(n_2206),
.B(n_187),
.Y(n_2392)
);

AO21x1_ASAP7_75t_L g2393 ( 
.A1(n_2291),
.A2(n_188),
.B(n_190),
.Y(n_2393)
);

OA22x2_ASAP7_75t_L g2394 ( 
.A1(n_1957),
.A2(n_191),
.B1(n_188),
.B2(n_190),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_2136),
.B(n_191),
.Y(n_2395)
);

OAI21x1_ASAP7_75t_SL g2396 ( 
.A1(n_2079),
.A2(n_192),
.B(n_193),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_1937),
.B(n_195),
.Y(n_2397)
);

BUFx8_ASAP7_75t_L g2398 ( 
.A(n_1946),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1938),
.B(n_196),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_1963),
.B(n_197),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_1939),
.B(n_197),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_1980),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1944),
.Y(n_2403)
);

INVx3_ASAP7_75t_L g2404 ( 
.A(n_1960),
.Y(n_2404)
);

INVx2_ASAP7_75t_SL g2405 ( 
.A(n_1959),
.Y(n_2405)
);

OA21x2_ASAP7_75t_L g2406 ( 
.A1(n_2014),
.A2(n_550),
.B(n_547),
.Y(n_2406)
);

A2O1A1Ixp33_ASAP7_75t_L g2407 ( 
.A1(n_2072),
.A2(n_201),
.B(n_198),
.C(n_200),
.Y(n_2407)
);

NOR2xp67_ASAP7_75t_L g2408 ( 
.A(n_1973),
.B(n_201),
.Y(n_2408)
);

AOI21xp5_ASAP7_75t_L g2409 ( 
.A1(n_2029),
.A2(n_553),
.B(n_552),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2019),
.B(n_203),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_1986),
.B(n_204),
.Y(n_2411)
);

AO21x1_ASAP7_75t_L g2412 ( 
.A1(n_2291),
.A2(n_204),
.B(n_205),
.Y(n_2412)
);

CKINVDCx20_ASAP7_75t_R g2413 ( 
.A(n_2066),
.Y(n_2413)
);

AOI21xp5_ASAP7_75t_L g2414 ( 
.A1(n_2035),
.A2(n_556),
.B(n_555),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_1992),
.B(n_2041),
.Y(n_2415)
);

OA22x2_ASAP7_75t_L g2416 ( 
.A1(n_1957),
.A2(n_210),
.B1(n_206),
.B2(n_208),
.Y(n_2416)
);

OAI221xp5_ASAP7_75t_L g2417 ( 
.A1(n_2236),
.A2(n_206),
.B1(n_211),
.B2(n_212),
.C(n_213),
.Y(n_2417)
);

AO31x2_ASAP7_75t_L g2418 ( 
.A1(n_2245),
.A2(n_213),
.A3(n_211),
.B(n_212),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_1963),
.B(n_214),
.Y(n_2419)
);

BUFx2_ASAP7_75t_L g2420 ( 
.A(n_2161),
.Y(n_2420)
);

AOI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_1982),
.A2(n_558),
.B(n_557),
.Y(n_2421)
);

INVx3_ASAP7_75t_L g2422 ( 
.A(n_2159),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2059),
.B(n_214),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_1967),
.B(n_215),
.Y(n_2424)
);

AO31x2_ASAP7_75t_L g2425 ( 
.A1(n_2245),
.A2(n_218),
.A3(n_216),
.B(n_217),
.Y(n_2425)
);

OAI21xp33_ASAP7_75t_L g2426 ( 
.A1(n_2223),
.A2(n_219),
.B(n_220),
.Y(n_2426)
);

OAI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_1967),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_2427)
);

OR2x6_ASAP7_75t_L g2428 ( 
.A(n_2159),
.B(n_221),
.Y(n_2428)
);

OAI21xp5_ASAP7_75t_L g2429 ( 
.A1(n_2005),
.A2(n_222),
.B(n_223),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_1932),
.B(n_222),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_1935),
.B(n_223),
.Y(n_2431)
);

NAND3x1_ASAP7_75t_L g2432 ( 
.A(n_2087),
.B(n_224),
.C(n_227),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2105),
.B(n_228),
.Y(n_2433)
);

A2O1A1Ixp33_ASAP7_75t_L g2434 ( 
.A1(n_2133),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_1947),
.B(n_229),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_1947),
.B(n_230),
.Y(n_2436)
);

OAI21x1_ASAP7_75t_L g2437 ( 
.A1(n_2219),
.A2(n_570),
.B(n_568),
.Y(n_2437)
);

INVx3_ASAP7_75t_L g2438 ( 
.A(n_2159),
.Y(n_2438)
);

BUFx2_ASAP7_75t_L g2439 ( 
.A(n_1959),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2084),
.B(n_231),
.Y(n_2440)
);

O2A1O1Ixp5_ASAP7_75t_L g2441 ( 
.A1(n_2002),
.A2(n_573),
.B(n_577),
.C(n_571),
.Y(n_2441)
);

AOI21xp5_ASAP7_75t_L g2442 ( 
.A1(n_2283),
.A2(n_2006),
.B(n_1945),
.Y(n_2442)
);

INVx3_ASAP7_75t_L g2443 ( 
.A(n_2173),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_1958),
.Y(n_2444)
);

NAND3x1_ASAP7_75t_L g2445 ( 
.A(n_2099),
.B(n_2295),
.C(n_2153),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2027),
.B(n_232),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2030),
.B(n_233),
.Y(n_2447)
);

AOI21x1_ASAP7_75t_L g2448 ( 
.A1(n_2103),
.A2(n_2130),
.B(n_2171),
.Y(n_2448)
);

OA21x2_ASAP7_75t_L g2449 ( 
.A1(n_2290),
.A2(n_581),
.B(n_578),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2166),
.Y(n_2450)
);

OAI21x1_ASAP7_75t_L g2451 ( 
.A1(n_2221),
.A2(n_583),
.B(n_582),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_1997),
.B(n_234),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2180),
.B(n_235),
.Y(n_2453)
);

AOI21xp5_ASAP7_75t_L g2454 ( 
.A1(n_1991),
.A2(n_591),
.B(n_588),
.Y(n_2454)
);

BUFx8_ASAP7_75t_L g2455 ( 
.A(n_1970),
.Y(n_2455)
);

INVx2_ASAP7_75t_SL g2456 ( 
.A(n_2017),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_SL g2457 ( 
.A(n_2057),
.B(n_236),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2039),
.B(n_240),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2266),
.B(n_241),
.Y(n_2459)
);

AOI21x1_ASAP7_75t_L g2460 ( 
.A1(n_2103),
.A2(n_596),
.B(n_594),
.Y(n_2460)
);

BUFx10_ASAP7_75t_L g2461 ( 
.A(n_2036),
.Y(n_2461)
);

OAI21x1_ASAP7_75t_L g2462 ( 
.A1(n_1988),
.A2(n_597),
.B(n_242),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_L g2463 ( 
.A(n_2224),
.B(n_242),
.Y(n_2463)
);

BUFx6f_ASAP7_75t_L g2464 ( 
.A(n_1958),
.Y(n_2464)
);

OAI21x1_ASAP7_75t_L g2465 ( 
.A1(n_1988),
.A2(n_243),
.B(n_244),
.Y(n_2465)
);

OAI21xp5_ASAP7_75t_L g2466 ( 
.A1(n_2005),
.A2(n_245),
.B(n_247),
.Y(n_2466)
);

AOI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_2001),
.A2(n_245),
.B(n_249),
.Y(n_2467)
);

AOI211x1_ASAP7_75t_L g2468 ( 
.A1(n_2145),
.A2(n_2081),
.B(n_2257),
.C(n_2270),
.Y(n_2468)
);

NAND3xp33_ASAP7_75t_L g2469 ( 
.A(n_2175),
.B(n_249),
.C(n_250),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_2003),
.A2(n_250),
.B(n_251),
.Y(n_2470)
);

INVxp67_ASAP7_75t_L g2471 ( 
.A(n_2253),
.Y(n_2471)
);

OAI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2056),
.A2(n_251),
.B(n_252),
.Y(n_2472)
);

OAI22xp5_ASAP7_75t_L g2473 ( 
.A1(n_2254),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_2473)
);

CKINVDCx8_ASAP7_75t_R g2474 ( 
.A(n_2127),
.Y(n_2474)
);

AOI21xp5_ASAP7_75t_L g2475 ( 
.A1(n_1993),
.A2(n_253),
.B(n_254),
.Y(n_2475)
);

INVxp67_ASAP7_75t_SL g2476 ( 
.A(n_2111),
.Y(n_2476)
);

AND2x4_ASAP7_75t_L g2477 ( 
.A(n_2033),
.B(n_256),
.Y(n_2477)
);

OAI21x1_ASAP7_75t_L g2478 ( 
.A1(n_2268),
.A2(n_257),
.B(n_258),
.Y(n_2478)
);

OAI22xp5_ASAP7_75t_L g2479 ( 
.A1(n_2254),
.A2(n_259),
.B1(n_262),
.B2(n_263),
.Y(n_2479)
);

BUFx6f_ASAP7_75t_L g2480 ( 
.A(n_1958),
.Y(n_2480)
);

AO31x2_ASAP7_75t_L g2481 ( 
.A1(n_2212),
.A2(n_259),
.A3(n_263),
.B(n_265),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2057),
.B(n_266),
.Y(n_2482)
);

OAI21x1_ASAP7_75t_L g2483 ( 
.A1(n_2199),
.A2(n_267),
.B(n_268),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2301),
.B(n_268),
.Y(n_2484)
);

AOI211x1_ASAP7_75t_L g2485 ( 
.A1(n_2145),
.A2(n_269),
.B(n_270),
.C(n_271),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2053),
.Y(n_2486)
);

OAI21x1_ASAP7_75t_SL g2487 ( 
.A1(n_2079),
.A2(n_269),
.B(n_271),
.Y(n_2487)
);

OAI21xp5_ASAP7_75t_L g2488 ( 
.A1(n_2202),
.A2(n_272),
.B(n_273),
.Y(n_2488)
);

OAI21xp5_ASAP7_75t_SL g2489 ( 
.A1(n_2191),
.A2(n_272),
.B(n_274),
.Y(n_2489)
);

OAI21xp5_ASAP7_75t_L g2490 ( 
.A1(n_2202),
.A2(n_275),
.B(n_276),
.Y(n_2490)
);

AO21x1_ASAP7_75t_L g2491 ( 
.A1(n_2257),
.A2(n_277),
.B(n_278),
.Y(n_2491)
);

AO31x2_ASAP7_75t_L g2492 ( 
.A1(n_2209),
.A2(n_279),
.A3(n_280),
.B(n_281),
.Y(n_2492)
);

AO31x2_ASAP7_75t_L g2493 ( 
.A1(n_2209),
.A2(n_280),
.A3(n_281),
.B(n_282),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_SL g2494 ( 
.A(n_2004),
.B(n_283),
.Y(n_2494)
);

AO31x2_ASAP7_75t_L g2495 ( 
.A1(n_2077),
.A2(n_284),
.A3(n_285),
.B(n_286),
.Y(n_2495)
);

OAI21x1_ASAP7_75t_L g2496 ( 
.A1(n_2213),
.A2(n_2216),
.B(n_1993),
.Y(n_2496)
);

OAI21xp5_ASAP7_75t_L g2497 ( 
.A1(n_2277),
.A2(n_285),
.B(n_287),
.Y(n_2497)
);

A2O1A1Ixp33_ASAP7_75t_L g2498 ( 
.A1(n_2150),
.A2(n_287),
.B(n_288),
.C(n_290),
.Y(n_2498)
);

BUFx2_ASAP7_75t_L g2499 ( 
.A(n_2131),
.Y(n_2499)
);

OAI21xp33_ASAP7_75t_L g2500 ( 
.A1(n_2150),
.A2(n_291),
.B(n_292),
.Y(n_2500)
);

AO21x2_ASAP7_75t_L g2501 ( 
.A1(n_2110),
.A2(n_293),
.B(n_294),
.Y(n_2501)
);

O2A1O1Ixp5_ASAP7_75t_L g2502 ( 
.A1(n_2201),
.A2(n_293),
.B(n_295),
.C(n_296),
.Y(n_2502)
);

AOI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_2078),
.A2(n_296),
.B(n_297),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2000),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2016),
.Y(n_2505)
);

AOI21xp5_ASAP7_75t_L g2506 ( 
.A1(n_2085),
.A2(n_298),
.B(n_299),
.Y(n_2506)
);

AO21x1_ASAP7_75t_L g2507 ( 
.A1(n_2081),
.A2(n_299),
.B(n_300),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2101),
.A2(n_300),
.B(n_301),
.Y(n_2508)
);

AOI21xp5_ASAP7_75t_L g2509 ( 
.A1(n_2102),
.A2(n_302),
.B(n_303),
.Y(n_2509)
);

OAI21x1_ASAP7_75t_L g2510 ( 
.A1(n_2216),
.A2(n_303),
.B(n_304),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2297),
.B(n_305),
.Y(n_2511)
);

INVx2_ASAP7_75t_SL g2512 ( 
.A(n_1998),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2020),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2021),
.Y(n_2514)
);

AO31x2_ASAP7_75t_L g2515 ( 
.A1(n_2249),
.A2(n_305),
.A3(n_306),
.B(n_307),
.Y(n_2515)
);

OAI21x1_ASAP7_75t_L g2516 ( 
.A1(n_1936),
.A2(n_307),
.B(n_308),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2046),
.Y(n_2517)
);

INVxp67_ASAP7_75t_SL g2518 ( 
.A(n_2111),
.Y(n_2518)
);

OAI21x1_ASAP7_75t_L g2519 ( 
.A1(n_1940),
.A2(n_311),
.B(n_312),
.Y(n_2519)
);

OAI21xp5_ASAP7_75t_L g2520 ( 
.A1(n_2279),
.A2(n_312),
.B(n_313),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2205),
.B(n_314),
.Y(n_2521)
);

OAI22xp5_ASAP7_75t_L g2522 ( 
.A1(n_2254),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_2522)
);

OAI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_1984),
.A2(n_315),
.B(n_316),
.Y(n_2523)
);

AOI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_2252),
.A2(n_317),
.B(n_319),
.Y(n_2524)
);

OAI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2254),
.A2(n_319),
.B1(n_321),
.B2(n_322),
.Y(n_2525)
);

OAI21x1_ASAP7_75t_L g2526 ( 
.A1(n_2229),
.A2(n_321),
.B(n_323),
.Y(n_2526)
);

AOI21xp5_ASAP7_75t_L g2527 ( 
.A1(n_2282),
.A2(n_324),
.B(n_325),
.Y(n_2527)
);

NAND3xp33_ASAP7_75t_L g2528 ( 
.A(n_2175),
.B(n_326),
.C(n_327),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2004),
.B(n_327),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2210),
.B(n_328),
.Y(n_2530)
);

OAI21x1_ASAP7_75t_L g2531 ( 
.A1(n_2232),
.A2(n_2244),
.B(n_2164),
.Y(n_2531)
);

AOI21x1_ASAP7_75t_L g2532 ( 
.A1(n_2130),
.A2(n_329),
.B(n_330),
.Y(n_2532)
);

OAI21xp5_ASAP7_75t_L g2533 ( 
.A1(n_2071),
.A2(n_2110),
.B(n_2123),
.Y(n_2533)
);

OAI21x1_ASAP7_75t_L g2534 ( 
.A1(n_2156),
.A2(n_329),
.B(n_330),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2054),
.Y(n_2535)
);

AOI21xp5_ASAP7_75t_L g2536 ( 
.A1(n_2142),
.A2(n_331),
.B(n_332),
.Y(n_2536)
);

CKINVDCx5p33_ASAP7_75t_R g2537 ( 
.A(n_2066),
.Y(n_2537)
);

AO32x2_ASAP7_75t_L g2538 ( 
.A1(n_2040),
.A2(n_331),
.A3(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_2538)
);

BUFx6f_ASAP7_75t_SL g2539 ( 
.A(n_2293),
.Y(n_2539)
);

BUFx12f_ASAP7_75t_L g2540 ( 
.A(n_2138),
.Y(n_2540)
);

NOR2xp33_ASAP7_75t_L g2541 ( 
.A(n_2068),
.B(n_334),
.Y(n_2541)
);

AOI21x1_ASAP7_75t_SL g2542 ( 
.A1(n_2292),
.A2(n_336),
.B(n_337),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2060),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2042),
.B(n_336),
.Y(n_2544)
);

OAI21x1_ASAP7_75t_L g2545 ( 
.A1(n_2156),
.A2(n_337),
.B(n_338),
.Y(n_2545)
);

OAI21x1_ASAP7_75t_L g2546 ( 
.A1(n_2164),
.A2(n_338),
.B(n_339),
.Y(n_2546)
);

AOI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_2149),
.A2(n_339),
.B1(n_341),
.B2(n_343),
.Y(n_2547)
);

OAI21x1_ASAP7_75t_L g2548 ( 
.A1(n_1974),
.A2(n_341),
.B(n_344),
.Y(n_2548)
);

BUFx6f_ASAP7_75t_L g2549 ( 
.A(n_1958),
.Y(n_2549)
);

BUFx2_ASAP7_75t_L g2550 ( 
.A(n_1955),
.Y(n_2550)
);

AOI21xp5_ASAP7_75t_L g2551 ( 
.A1(n_2143),
.A2(n_346),
.B(n_348),
.Y(n_2551)
);

OAI21x1_ASAP7_75t_L g2552 ( 
.A1(n_2025),
.A2(n_349),
.B(n_350),
.Y(n_2552)
);

OAI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2239),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_2553)
);

AO32x2_ASAP7_75t_L g2554 ( 
.A1(n_2040),
.A2(n_352),
.A3(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_2053),
.Y(n_2555)
);

INVx5_ASAP7_75t_L g2556 ( 
.A(n_2096),
.Y(n_2556)
);

AOI21xp5_ASAP7_75t_L g2557 ( 
.A1(n_2144),
.A2(n_358),
.B(n_359),
.Y(n_2557)
);

NAND2x1p5_ASAP7_75t_L g2558 ( 
.A(n_2183),
.B(n_360),
.Y(n_2558)
);

OAI21x1_ASAP7_75t_L g2559 ( 
.A1(n_2025),
.A2(n_2186),
.B(n_2168),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2063),
.B(n_361),
.Y(n_2560)
);

AOI21xp5_ASAP7_75t_L g2561 ( 
.A1(n_2146),
.A2(n_361),
.B(n_362),
.Y(n_2561)
);

OAI21xp5_ASAP7_75t_L g2562 ( 
.A1(n_2158),
.A2(n_363),
.B(n_364),
.Y(n_2562)
);

NAND2xp33_ASAP7_75t_SL g2563 ( 
.A(n_2247),
.B(n_363),
.Y(n_2563)
);

BUFx2_ASAP7_75t_L g2564 ( 
.A(n_2092),
.Y(n_2564)
);

AOI22xp33_ASAP7_75t_L g2565 ( 
.A1(n_2097),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_2565)
);

OA22x2_ASAP7_75t_L g2566 ( 
.A1(n_2293),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2065),
.B(n_369),
.Y(n_2567)
);

OAI21x1_ASAP7_75t_L g2568 ( 
.A1(n_2186),
.A2(n_371),
.B(n_373),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2207),
.B(n_371),
.Y(n_2569)
);

AOI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2258),
.A2(n_374),
.B(n_375),
.Y(n_2570)
);

OAI21xp5_ASAP7_75t_L g2571 ( 
.A1(n_2208),
.A2(n_374),
.B(n_377),
.Y(n_2571)
);

OAI21x1_ASAP7_75t_L g2572 ( 
.A1(n_2201),
.A2(n_377),
.B(n_378),
.Y(n_2572)
);

O2A1O1Ixp5_ASAP7_75t_L g2573 ( 
.A1(n_2296),
.A2(n_379),
.B(n_380),
.C(n_381),
.Y(n_2573)
);

OAI21x1_ASAP7_75t_L g2574 ( 
.A1(n_2044),
.A2(n_380),
.B(n_382),
.Y(n_2574)
);

AOI21xp5_ASAP7_75t_L g2575 ( 
.A1(n_2258),
.A2(n_382),
.B(n_384),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_1983),
.Y(n_2576)
);

OA21x2_ASAP7_75t_L g2577 ( 
.A1(n_2278),
.A2(n_384),
.B(n_385),
.Y(n_2577)
);

HB1xp67_ASAP7_75t_L g2578 ( 
.A(n_1979),
.Y(n_2578)
);

OAI21x1_ASAP7_75t_L g2579 ( 
.A1(n_2058),
.A2(n_391),
.B(n_392),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_1968),
.B(n_1953),
.Y(n_2580)
);

OAI21x1_ASAP7_75t_L g2581 ( 
.A1(n_2058),
.A2(n_392),
.B(n_393),
.Y(n_2581)
);

OAI21x1_ASAP7_75t_L g2582 ( 
.A1(n_2330),
.A2(n_2152),
.B(n_2083),
.Y(n_2582)
);

AOI221xp5_ASAP7_75t_L g2583 ( 
.A1(n_2310),
.A2(n_2187),
.B1(n_2162),
.B2(n_2269),
.C(n_2170),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2539),
.B(n_2009),
.Y(n_2584)
);

AOI22xp33_ASAP7_75t_L g2585 ( 
.A1(n_2539),
.A2(n_2239),
.B1(n_2165),
.B2(n_2190),
.Y(n_2585)
);

OAI21xp5_ASAP7_75t_L g2586 ( 
.A1(n_2338),
.A2(n_2243),
.B(n_2256),
.Y(n_2586)
);

OAI21x1_ASAP7_75t_L g2587 ( 
.A1(n_2339),
.A2(n_2152),
.B(n_2083),
.Y(n_2587)
);

OAI21xp5_ASAP7_75t_L g2588 ( 
.A1(n_2316),
.A2(n_2243),
.B(n_2256),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2403),
.Y(n_2589)
);

BUFx3_ASAP7_75t_L g2590 ( 
.A(n_2350),
.Y(n_2590)
);

OAI21x1_ASAP7_75t_L g2591 ( 
.A1(n_2496),
.A2(n_2259),
.B(n_2094),
.Y(n_2591)
);

OR2x6_ASAP7_75t_L g2592 ( 
.A(n_2428),
.B(n_2169),
.Y(n_2592)
);

NOR2xp67_ASAP7_75t_L g2593 ( 
.A(n_2556),
.B(n_2183),
.Y(n_2593)
);

AOI21xp5_ASAP7_75t_L g2594 ( 
.A1(n_2366),
.A2(n_2259),
.B(n_1962),
.Y(n_2594)
);

HB1xp67_ASAP7_75t_L g2595 ( 
.A(n_2331),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2323),
.B(n_1975),
.Y(n_2596)
);

AO21x2_ASAP7_75t_L g2597 ( 
.A1(n_2316),
.A2(n_2273),
.B(n_1975),
.Y(n_2597)
);

O2A1O1Ixp33_ASAP7_75t_L g2598 ( 
.A1(n_2310),
.A2(n_2007),
.B(n_2162),
.C(n_2293),
.Y(n_2598)
);

OAI21x1_ASAP7_75t_L g2599 ( 
.A1(n_2531),
.A2(n_2106),
.B(n_2080),
.Y(n_2599)
);

OAI21x1_ASAP7_75t_L g2600 ( 
.A1(n_2309),
.A2(n_2119),
.B(n_2118),
.Y(n_2600)
);

INVx6_ASAP7_75t_L g2601 ( 
.A(n_2398),
.Y(n_2601)
);

O2A1O1Ixp33_ASAP7_75t_SL g2602 ( 
.A1(n_2489),
.A2(n_2089),
.B(n_2095),
.C(n_2273),
.Y(n_2602)
);

INVx3_ASAP7_75t_SL g2603 ( 
.A(n_2345),
.Y(n_2603)
);

OA21x2_ASAP7_75t_L g2604 ( 
.A1(n_2462),
.A2(n_2010),
.B(n_2089),
.Y(n_2604)
);

OAI21x1_ASAP7_75t_L g2605 ( 
.A1(n_2559),
.A2(n_2179),
.B(n_2178),
.Y(n_2605)
);

NAND2x1p5_ASAP7_75t_L g2606 ( 
.A(n_2308),
.B(n_1949),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2323),
.B(n_2230),
.Y(n_2607)
);

NOR2x1_ASAP7_75t_SL g2608 ( 
.A(n_2354),
.B(n_2183),
.Y(n_2608)
);

OAI21xp33_ASAP7_75t_SL g2609 ( 
.A1(n_2566),
.A2(n_2095),
.B(n_2237),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2342),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2450),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2372),
.Y(n_2612)
);

OR2x2_ASAP7_75t_L g2613 ( 
.A(n_2580),
.B(n_2043),
.Y(n_2613)
);

OAI21xp5_ASAP7_75t_L g2614 ( 
.A1(n_2533),
.A2(n_2275),
.B(n_2267),
.Y(n_2614)
);

BUFx10_ASAP7_75t_L g2615 ( 
.A(n_2334),
.Y(n_2615)
);

AOI22xp5_ASAP7_75t_L g2616 ( 
.A1(n_2351),
.A2(n_2253),
.B1(n_2061),
.B2(n_2097),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2415),
.B(n_2231),
.Y(n_2617)
);

OAI211xp5_ASAP7_75t_L g2618 ( 
.A1(n_2489),
.A2(n_2092),
.B(n_2100),
.C(n_1951),
.Y(n_2618)
);

BUFx2_ASAP7_75t_L g2619 ( 
.A(n_2455),
.Y(n_2619)
);

O2A1O1Ixp33_ASAP7_75t_L g2620 ( 
.A1(n_2498),
.A2(n_2269),
.B(n_2181),
.C(n_2112),
.Y(n_2620)
);

OAI22xp33_ASAP7_75t_L g2621 ( 
.A1(n_2327),
.A2(n_2061),
.B1(n_2242),
.B2(n_1998),
.Y(n_2621)
);

OAI21x1_ASAP7_75t_L g2622 ( 
.A1(n_2437),
.A2(n_2126),
.B(n_2122),
.Y(n_2622)
);

OAI21x1_ASAP7_75t_SL g2623 ( 
.A1(n_2553),
.A2(n_2214),
.B(n_2284),
.Y(n_2623)
);

AO31x2_ASAP7_75t_L g2624 ( 
.A1(n_2333),
.A2(n_2193),
.A3(n_2280),
.B(n_2154),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_2413),
.Y(n_2625)
);

O2A1O1Ixp33_ASAP7_75t_L g2626 ( 
.A1(n_2553),
.A2(n_2114),
.B(n_2113),
.C(n_2037),
.Y(n_2626)
);

OR2x2_ASAP7_75t_L g2627 ( 
.A(n_2302),
.B(n_2226),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2452),
.B(n_2132),
.Y(n_2628)
);

CKINVDCx11_ASAP7_75t_R g2629 ( 
.A(n_2474),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2306),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2415),
.B(n_2533),
.Y(n_2631)
);

OAI21x1_ASAP7_75t_L g2632 ( 
.A1(n_2451),
.A2(n_2300),
.B(n_2024),
.Y(n_2632)
);

OAI21x1_ASAP7_75t_L g2633 ( 
.A1(n_2442),
.A2(n_2300),
.B(n_2049),
.Y(n_2633)
);

AOI22x1_ASAP7_75t_L g2634 ( 
.A1(n_2362),
.A2(n_2115),
.B1(n_2177),
.B2(n_2189),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2317),
.Y(n_2635)
);

OA21x2_ASAP7_75t_L g2636 ( 
.A1(n_2465),
.A2(n_2010),
.B(n_2082),
.Y(n_2636)
);

OAI221xp5_ASAP7_75t_L g2637 ( 
.A1(n_2332),
.A2(n_2426),
.B1(n_2353),
.B2(n_2500),
.C(n_2329),
.Y(n_2637)
);

AOI22xp33_ASAP7_75t_L g2638 ( 
.A1(n_2563),
.A2(n_2190),
.B1(n_2192),
.B2(n_2165),
.Y(n_2638)
);

OAI21x1_ASAP7_75t_L g2639 ( 
.A1(n_2328),
.A2(n_2109),
.B(n_2075),
.Y(n_2639)
);

OAI21x1_ASAP7_75t_L g2640 ( 
.A1(n_2335),
.A2(n_2022),
.B(n_2067),
.Y(n_2640)
);

OR2x6_ASAP7_75t_L g2641 ( 
.A(n_2428),
.B(n_2380),
.Y(n_2641)
);

OAI221xp5_ASAP7_75t_L g2642 ( 
.A1(n_2329),
.A2(n_2241),
.B1(n_2220),
.B2(n_2191),
.C(n_2203),
.Y(n_2642)
);

BUFx2_ASAP7_75t_L g2643 ( 
.A(n_2398),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2370),
.Y(n_2644)
);

OAI21x1_ASAP7_75t_L g2645 ( 
.A1(n_2346),
.A2(n_2357),
.B(n_2356),
.Y(n_2645)
);

AND2x4_ASAP7_75t_L g2646 ( 
.A(n_2308),
.B(n_2183),
.Y(n_2646)
);

BUFx3_ASAP7_75t_L g2647 ( 
.A(n_2376),
.Y(n_2647)
);

AOI21x1_ASAP7_75t_L g2648 ( 
.A1(n_2448),
.A2(n_2074),
.B(n_2228),
.Y(n_2648)
);

AO21x2_ASAP7_75t_L g2649 ( 
.A1(n_2312),
.A2(n_2082),
.B(n_2220),
.Y(n_2649)
);

OA21x2_ASAP7_75t_L g2650 ( 
.A1(n_2475),
.A2(n_2012),
.B(n_2241),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2471),
.B(n_2281),
.Y(n_2651)
);

OR2x2_ASAP7_75t_L g2652 ( 
.A(n_2390),
.B(n_2341),
.Y(n_2652)
);

OAI21x1_ASAP7_75t_L g2653 ( 
.A1(n_2359),
.A2(n_2015),
.B(n_2008),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2348),
.B(n_2012),
.Y(n_2654)
);

NAND2x1p5_ASAP7_75t_L g2655 ( 
.A(n_2439),
.B(n_1990),
.Y(n_2655)
);

AO21x2_ASAP7_75t_L g2656 ( 
.A1(n_2312),
.A2(n_2051),
.B(n_1989),
.Y(n_2656)
);

OR2x6_ASAP7_75t_L g2657 ( 
.A(n_2428),
.B(n_2169),
.Y(n_2657)
);

OR2x2_ASAP7_75t_L g2658 ( 
.A(n_2550),
.B(n_2163),
.Y(n_2658)
);

INVx3_ASAP7_75t_L g2659 ( 
.A(n_2556),
.Y(n_2659)
);

AND2x4_ASAP7_75t_L g2660 ( 
.A(n_2314),
.B(n_2172),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2348),
.B(n_2234),
.Y(n_2661)
);

NAND2x1p5_ASAP7_75t_L g2662 ( 
.A(n_2334),
.B(n_1954),
.Y(n_2662)
);

OAI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2468),
.A2(n_2169),
.B1(n_2242),
.B2(n_2294),
.Y(n_2663)
);

INVx3_ASAP7_75t_L g2664 ( 
.A(n_2556),
.Y(n_2664)
);

OAI21xp5_ASAP7_75t_L g2665 ( 
.A1(n_2304),
.A2(n_2196),
.B(n_2195),
.Y(n_2665)
);

NOR2xp33_ASAP7_75t_L g2666 ( 
.A(n_2564),
.B(n_2031),
.Y(n_2666)
);

BUFx6f_ASAP7_75t_L g2667 ( 
.A(n_2444),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2543),
.Y(n_2668)
);

AOI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2327),
.A2(n_2163),
.B1(n_2192),
.B2(n_2238),
.Y(n_2669)
);

A2O1A1Ixp33_ASAP7_75t_L g2670 ( 
.A1(n_2429),
.A2(n_2286),
.B(n_2203),
.C(n_2184),
.Y(n_2670)
);

BUFx2_ASAP7_75t_R g2671 ( 
.A(n_2576),
.Y(n_2671)
);

NOR2xp67_ASAP7_75t_L g2672 ( 
.A(n_2556),
.B(n_1954),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2385),
.Y(n_2673)
);

OAI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2420),
.A2(n_2294),
.B1(n_2176),
.B2(n_2286),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2385),
.Y(n_2675)
);

BUFx2_ASAP7_75t_L g2676 ( 
.A(n_2476),
.Y(n_2676)
);

NAND2xp33_ASAP7_75t_L g2677 ( 
.A(n_2405),
.B(n_2247),
.Y(n_2677)
);

AOI22xp33_ASAP7_75t_L g2678 ( 
.A1(n_2337),
.A2(n_2499),
.B1(n_2566),
.B2(n_2238),
.Y(n_2678)
);

OA21x2_ASAP7_75t_L g2679 ( 
.A1(n_2313),
.A2(n_2051),
.B(n_1989),
.Y(n_2679)
);

BUFx3_ASAP7_75t_L g2680 ( 
.A(n_2456),
.Y(n_2680)
);

AOI22xp33_ASAP7_75t_L g2681 ( 
.A1(n_2368),
.A2(n_2261),
.B1(n_2107),
.B2(n_2108),
.Y(n_2681)
);

AO32x2_ASAP7_75t_L g2682 ( 
.A1(n_2473),
.A2(n_2204),
.A3(n_2225),
.B1(n_2090),
.B2(n_2185),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2504),
.Y(n_2683)
);

INVx2_ASAP7_75t_SL g2684 ( 
.A(n_2461),
.Y(n_2684)
);

AOI22xp33_ASAP7_75t_L g2685 ( 
.A1(n_2379),
.A2(n_2261),
.B1(n_2287),
.B2(n_2240),
.Y(n_2685)
);

BUFx3_ASAP7_75t_L g2686 ( 
.A(n_2537),
.Y(n_2686)
);

A2O1A1Ixp33_ASAP7_75t_L g2687 ( 
.A1(n_2429),
.A2(n_2264),
.B(n_2276),
.C(n_2218),
.Y(n_2687)
);

AO21x2_ASAP7_75t_L g2688 ( 
.A1(n_2313),
.A2(n_2298),
.B(n_2100),
.Y(n_2688)
);

OAI21x1_ASAP7_75t_SL g2689 ( 
.A1(n_2466),
.A2(n_2141),
.B(n_2250),
.Y(n_2689)
);

AND2x4_ASAP7_75t_L g2690 ( 
.A(n_2314),
.B(n_1954),
.Y(n_2690)
);

BUFx3_ASAP7_75t_L g2691 ( 
.A(n_2461),
.Y(n_2691)
);

AOI21x1_ASAP7_75t_L g2692 ( 
.A1(n_2375),
.A2(n_2388),
.B(n_2449),
.Y(n_2692)
);

OAI221xp5_ASAP7_75t_L g2693 ( 
.A1(n_2488),
.A2(n_2198),
.B1(n_2263),
.B2(n_2045),
.C(n_1965),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2347),
.B(n_2036),
.Y(n_2694)
);

OAI21x1_ASAP7_75t_L g2695 ( 
.A1(n_2318),
.A2(n_2088),
.B(n_1962),
.Y(n_2695)
);

OAI21x1_ASAP7_75t_L g2696 ( 
.A1(n_2320),
.A2(n_2088),
.B(n_2011),
.Y(n_2696)
);

OAI21x1_ASAP7_75t_L g2697 ( 
.A1(n_2378),
.A2(n_2088),
.B(n_2011),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2410),
.B(n_2298),
.Y(n_2698)
);

A2O1A1Ixp33_ASAP7_75t_L g2699 ( 
.A1(n_2466),
.A2(n_2055),
.B(n_2294),
.C(n_2289),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_SL g2700 ( 
.A(n_2558),
.B(n_2294),
.Y(n_2700)
);

AND2x4_ASAP7_75t_L g2701 ( 
.A(n_2355),
.B(n_1954),
.Y(n_2701)
);

AOI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2445),
.A2(n_1933),
.B1(n_2055),
.B2(n_2167),
.Y(n_2702)
);

OAI21x1_ASAP7_75t_L g2703 ( 
.A1(n_2384),
.A2(n_2088),
.B(n_1961),
.Y(n_2703)
);

OAI21x1_ASAP7_75t_L g2704 ( 
.A1(n_2542),
.A2(n_2441),
.B(n_2387),
.Y(n_2704)
);

OAI21x1_ASAP7_75t_L g2705 ( 
.A1(n_2460),
.A2(n_2086),
.B(n_1961),
.Y(n_2705)
);

OAI21x1_ASAP7_75t_SL g2706 ( 
.A1(n_2491),
.A2(n_2250),
.B(n_2193),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2505),
.Y(n_2707)
);

AOI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2321),
.A2(n_2134),
.B(n_2064),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2477),
.B(n_2235),
.Y(n_2709)
);

NOR2xp67_ASAP7_75t_L g2710 ( 
.A(n_2473),
.B(n_2034),
.Y(n_2710)
);

AOI21xp5_ASAP7_75t_L g2711 ( 
.A1(n_2343),
.A2(n_2424),
.B(n_2389),
.Y(n_2711)
);

NOR2x1p5_ASAP7_75t_L g2712 ( 
.A(n_2518),
.B(n_1933),
.Y(n_2712)
);

OR2x2_ASAP7_75t_L g2713 ( 
.A(n_2578),
.B(n_2137),
.Y(n_2713)
);

OAI21x1_ASAP7_75t_SL g2714 ( 
.A1(n_2396),
.A2(n_2096),
.B(n_2215),
.Y(n_2714)
);

OAI21x1_ASAP7_75t_L g2715 ( 
.A1(n_2386),
.A2(n_1961),
.B(n_2011),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2513),
.Y(n_2716)
);

BUFx2_ASAP7_75t_L g2717 ( 
.A(n_2355),
.Y(n_2717)
);

INVx2_ASAP7_75t_SL g2718 ( 
.A(n_2443),
.Y(n_2718)
);

OAI21xp5_ASAP7_75t_L g2719 ( 
.A1(n_2358),
.A2(n_2289),
.B(n_2215),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2397),
.Y(n_2720)
);

INVx2_ASAP7_75t_SL g2721 ( 
.A(n_2443),
.Y(n_2721)
);

BUFx2_ASAP7_75t_L g2722 ( 
.A(n_2319),
.Y(n_2722)
);

AOI21xp5_ASAP7_75t_L g2723 ( 
.A1(n_2424),
.A2(n_2086),
.B(n_2026),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2397),
.Y(n_2724)
);

AOI22xp33_ASAP7_75t_L g2725 ( 
.A1(n_2469),
.A2(n_2289),
.B1(n_2235),
.B2(n_2167),
.Y(n_2725)
);

AND2x2_ASAP7_75t_L g2726 ( 
.A(n_2477),
.B(n_1966),
.Y(n_2726)
);

OA21x2_ASAP7_75t_L g2727 ( 
.A1(n_2478),
.A2(n_2050),
.B(n_2076),
.Y(n_2727)
);

AOI22xp33_ASAP7_75t_L g2728 ( 
.A1(n_2528),
.A2(n_2289),
.B1(n_2032),
.B2(n_2076),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2433),
.B(n_2435),
.Y(n_2729)
);

AOI22xp5_ASAP7_75t_L g2730 ( 
.A1(n_2427),
.A2(n_1966),
.B1(n_2096),
.B2(n_2032),
.Y(n_2730)
);

AOI21xp5_ASAP7_75t_L g2731 ( 
.A1(n_2421),
.A2(n_2128),
.B(n_2064),
.Y(n_2731)
);

OAI21x1_ASAP7_75t_L g2732 ( 
.A1(n_2311),
.A2(n_2572),
.B(n_2526),
.Y(n_2732)
);

BUFx2_ASAP7_75t_R g2733 ( 
.A(n_2369),
.Y(n_2733)
);

OA21x2_ASAP7_75t_L g2734 ( 
.A1(n_2483),
.A2(n_2050),
.B(n_2215),
.Y(n_2734)
);

AOI22xp5_ASAP7_75t_L g2735 ( 
.A1(n_2427),
.A2(n_2479),
.B1(n_2525),
.B2(n_2522),
.Y(n_2735)
);

OR2x2_ASAP7_75t_L g2736 ( 
.A(n_2569),
.B(n_2023),
.Y(n_2736)
);

OAI22xp5_ASAP7_75t_L g2737 ( 
.A1(n_2479),
.A2(n_2148),
.B1(n_2034),
.B2(n_2157),
.Y(n_2737)
);

OAI21x1_ASAP7_75t_SL g2738 ( 
.A1(n_2487),
.A2(n_2096),
.B(n_2215),
.Y(n_2738)
);

AOI221xp5_ASAP7_75t_L g2739 ( 
.A1(n_2485),
.A2(n_2023),
.B1(n_1996),
.B2(n_2018),
.C(n_2272),
.Y(n_2739)
);

A2O1A1Ixp33_ASAP7_75t_L g2740 ( 
.A1(n_2488),
.A2(n_1996),
.B(n_2018),
.C(n_2034),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2514),
.Y(n_2741)
);

OAI21xp5_ASAP7_75t_L g2742 ( 
.A1(n_2358),
.A2(n_2215),
.B(n_2096),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2399),
.Y(n_2743)
);

INVx2_ASAP7_75t_SL g2744 ( 
.A(n_2512),
.Y(n_2744)
);

OAI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_2522),
.A2(n_2148),
.B1(n_2157),
.B2(n_2053),
.Y(n_2745)
);

OR2x6_ASAP7_75t_L g2746 ( 
.A(n_2319),
.B(n_2128),
.Y(n_2746)
);

OAI21x1_ASAP7_75t_L g2747 ( 
.A1(n_2510),
.A2(n_2449),
.B(n_2409),
.Y(n_2747)
);

BUFx5_ASAP7_75t_L g2748 ( 
.A(n_2444),
.Y(n_2748)
);

OAI22xp5_ASAP7_75t_SL g2749 ( 
.A1(n_2392),
.A2(n_2541),
.B1(n_2395),
.B2(n_2525),
.Y(n_2749)
);

AO21x2_ASAP7_75t_L g2750 ( 
.A1(n_2352),
.A2(n_2134),
.B(n_2064),
.Y(n_2750)
);

OR2x6_ASAP7_75t_L g2751 ( 
.A(n_2558),
.B(n_2134),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2436),
.B(n_395),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2422),
.B(n_2148),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2453),
.B(n_2544),
.Y(n_2754)
);

AOI22x1_ASAP7_75t_L g2755 ( 
.A1(n_2527),
.A2(n_2272),
.B1(n_2121),
.B2(n_2151),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2517),
.Y(n_2756)
);

A2O1A1Ixp33_ASAP7_75t_L g2757 ( 
.A1(n_2490),
.A2(n_2523),
.B(n_2472),
.C(n_2562),
.Y(n_2757)
);

OAI221xp5_ASAP7_75t_L g2758 ( 
.A1(n_2490),
.A2(n_2157),
.B1(n_2222),
.B2(n_2151),
.C(n_2116),
.Y(n_2758)
);

OAI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2494),
.A2(n_2151),
.B1(n_2062),
.B2(n_2222),
.Y(n_2759)
);

BUFx6f_ASAP7_75t_L g2760 ( 
.A(n_2444),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2399),
.Y(n_2761)
);

AOI22xp33_ASAP7_75t_L g2762 ( 
.A1(n_2373),
.A2(n_2070),
.B1(n_2222),
.B2(n_2062),
.Y(n_2762)
);

AO21x2_ASAP7_75t_L g2763 ( 
.A1(n_2352),
.A2(n_2070),
.B(n_396),
.Y(n_2763)
);

AO21x1_ASAP7_75t_L g2764 ( 
.A1(n_2457),
.A2(n_395),
.B(n_397),
.Y(n_2764)
);

BUFx6f_ASAP7_75t_L g2765 ( 
.A(n_2464),
.Y(n_2765)
);

AOI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2406),
.A2(n_2070),
.B(n_401),
.Y(n_2766)
);

OAI21x1_ASAP7_75t_L g2767 ( 
.A1(n_2568),
.A2(n_2070),
.B(n_402),
.Y(n_2767)
);

AOI21x1_ASAP7_75t_L g2768 ( 
.A1(n_2406),
.A2(n_399),
.B(n_402),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_2540),
.Y(n_2769)
);

OAI22xp5_ASAP7_75t_L g2770 ( 
.A1(n_2529),
.A2(n_399),
.B1(n_403),
.B2(n_404),
.Y(n_2770)
);

OAI21x1_ASAP7_75t_L g2771 ( 
.A1(n_2414),
.A2(n_403),
.B(n_405),
.Y(n_2771)
);

CKINVDCx20_ASAP7_75t_R g2772 ( 
.A(n_2402),
.Y(n_2772)
);

BUFx12f_ASAP7_75t_L g2773 ( 
.A(n_2629),
.Y(n_2773)
);

AOI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2700),
.A2(n_2382),
.B(n_2365),
.Y(n_2774)
);

INVx4_ASAP7_75t_L g2775 ( 
.A(n_2601),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2589),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2595),
.B(n_2400),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2611),
.B(n_2419),
.Y(n_2778)
);

INVx6_ASAP7_75t_L g2779 ( 
.A(n_2601),
.Y(n_2779)
);

OR2x2_ASAP7_75t_L g2780 ( 
.A(n_2652),
.B(n_2610),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2630),
.Y(n_2781)
);

OR2x2_ASAP7_75t_L g2782 ( 
.A(n_2627),
.B(n_2569),
.Y(n_2782)
);

INVx4_ASAP7_75t_L g2783 ( 
.A(n_2603),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2635),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2644),
.B(n_2401),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_SL g2786 ( 
.A(n_2616),
.B(n_2507),
.Y(n_2786)
);

OAI22xp5_ASAP7_75t_L g2787 ( 
.A1(n_2616),
.A2(n_2394),
.B1(n_2373),
.B2(n_2416),
.Y(n_2787)
);

OR2x2_ASAP7_75t_L g2788 ( 
.A(n_2613),
.B(n_2729),
.Y(n_2788)
);

INVx4_ASAP7_75t_L g2789 ( 
.A(n_2590),
.Y(n_2789)
);

OAI22xp33_ASAP7_75t_L g2790 ( 
.A1(n_2669),
.A2(n_2394),
.B1(n_2416),
.B2(n_2547),
.Y(n_2790)
);

CKINVDCx20_ASAP7_75t_R g2791 ( 
.A(n_2772),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2668),
.B(n_2673),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2675),
.B(n_2401),
.Y(n_2793)
);

INVx3_ASAP7_75t_L g2794 ( 
.A(n_2646),
.Y(n_2794)
);

O2A1O1Ixp33_ASAP7_75t_L g2795 ( 
.A1(n_2670),
.A2(n_2360),
.B(n_2336),
.C(n_2407),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2612),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2720),
.B(n_2411),
.Y(n_2797)
);

AOI22xp33_ASAP7_75t_SL g2798 ( 
.A1(n_2749),
.A2(n_2501),
.B1(n_2523),
.B2(n_2520),
.Y(n_2798)
);

OAI22xp33_ASAP7_75t_L g2799 ( 
.A1(n_2669),
.A2(n_2482),
.B1(n_2408),
.B2(n_2391),
.Y(n_2799)
);

AOI22xp33_ASAP7_75t_L g2800 ( 
.A1(n_2749),
.A2(n_2463),
.B1(n_2417),
.B2(n_2412),
.Y(n_2800)
);

INVx2_ASAP7_75t_SL g2801 ( 
.A(n_2643),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2724),
.B(n_2411),
.Y(n_2802)
);

NAND2xp33_ASAP7_75t_R g2803 ( 
.A(n_2619),
.B(n_2438),
.Y(n_2803)
);

AOI22xp33_ASAP7_75t_L g2804 ( 
.A1(n_2693),
.A2(n_2393),
.B1(n_2565),
.B2(n_2520),
.Y(n_2804)
);

OAI21xp5_ASAP7_75t_L g2805 ( 
.A1(n_2586),
.A2(n_2757),
.B(n_2588),
.Y(n_2805)
);

BUFx12f_ASAP7_75t_L g2806 ( 
.A(n_2625),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2717),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2743),
.B(n_2446),
.Y(n_2808)
);

AOI221xp5_ASAP7_75t_L g2809 ( 
.A1(n_2598),
.A2(n_2367),
.B1(n_2497),
.B2(n_2472),
.C(n_2562),
.Y(n_2809)
);

AOI22xp33_ASAP7_75t_L g2810 ( 
.A1(n_2693),
.A2(n_2497),
.B1(n_2367),
.B2(n_2571),
.Y(n_2810)
);

AOI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2735),
.A2(n_2618),
.B1(n_2583),
.B2(n_2642),
.Y(n_2811)
);

AOI221xp5_ASAP7_75t_L g2812 ( 
.A1(n_2621),
.A2(n_2364),
.B1(n_2349),
.B2(n_2521),
.C(n_2530),
.Y(n_2812)
);

OR2x2_ASAP7_75t_L g2813 ( 
.A(n_2713),
.B(n_2440),
.Y(n_2813)
);

AOI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2735),
.A2(n_2432),
.B1(n_2430),
.B2(n_2431),
.Y(n_2814)
);

OAI22x1_ASAP7_75t_L g2815 ( 
.A1(n_2676),
.A2(n_2363),
.B1(n_2532),
.B2(n_2577),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2683),
.Y(n_2816)
);

CKINVDCx5p33_ASAP7_75t_R g2817 ( 
.A(n_2769),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2707),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2761),
.B(n_2446),
.Y(n_2819)
);

AOI22xp33_ASAP7_75t_L g2820 ( 
.A1(n_2642),
.A2(n_2571),
.B1(n_2374),
.B2(n_2501),
.Y(n_2820)
);

BUFx3_ASAP7_75t_L g2821 ( 
.A(n_2647),
.Y(n_2821)
);

OA21x2_ASAP7_75t_L g2822 ( 
.A1(n_2747),
.A2(n_2519),
.B(n_2516),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2634),
.B(n_2374),
.Y(n_2823)
);

OAI22xp33_ASAP7_75t_L g2824 ( 
.A1(n_2641),
.A2(n_2340),
.B1(n_2326),
.B2(n_2344),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_SL g2825 ( 
.A(n_2615),
.B(n_2524),
.Y(n_2825)
);

NAND2x1p5_ASAP7_75t_L g2826 ( 
.A(n_2672),
.B(n_2438),
.Y(n_2826)
);

AOI22xp33_ASAP7_75t_L g2827 ( 
.A1(n_2628),
.A2(n_2459),
.B1(n_2521),
.B2(n_2530),
.Y(n_2827)
);

AOI22xp33_ASAP7_75t_L g2828 ( 
.A1(n_2586),
.A2(n_2551),
.B1(n_2536),
.B2(n_2557),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2617),
.B(n_2447),
.Y(n_2829)
);

HB1xp67_ASAP7_75t_L g2830 ( 
.A(n_2658),
.Y(n_2830)
);

HB1xp67_ASAP7_75t_L g2831 ( 
.A(n_2716),
.Y(n_2831)
);

OAI22xp5_ASAP7_75t_L g2832 ( 
.A1(n_2730),
.A2(n_2315),
.B1(n_2434),
.B2(n_2361),
.Y(n_2832)
);

INVx2_ASAP7_75t_SL g2833 ( 
.A(n_2680),
.Y(n_2833)
);

AOI221xp5_ASAP7_75t_L g2834 ( 
.A1(n_2609),
.A2(n_2484),
.B1(n_2511),
.B2(n_2508),
.C(n_2509),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2741),
.Y(n_2835)
);

AOI21xp5_ASAP7_75t_L g2836 ( 
.A1(n_2700),
.A2(n_2365),
.B(n_2325),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2617),
.B(n_2447),
.Y(n_2837)
);

AOI22xp5_ASAP7_75t_L g2838 ( 
.A1(n_2596),
.A2(n_2431),
.B1(n_2430),
.B2(n_2303),
.Y(n_2838)
);

OAI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2588),
.A2(n_2573),
.B(n_2502),
.Y(n_2839)
);

NOR3xp33_ASAP7_75t_SL g2840 ( 
.A(n_2584),
.B(n_2484),
.C(n_2511),
.Y(n_2840)
);

OAI22xp5_ASAP7_75t_L g2841 ( 
.A1(n_2730),
.A2(n_2324),
.B1(n_2325),
.B2(n_2344),
.Y(n_2841)
);

AOI22xp33_ASAP7_75t_L g2842 ( 
.A1(n_2638),
.A2(n_2561),
.B1(n_2506),
.B2(n_2503),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2756),
.Y(n_2843)
);

AOI22xp33_ASAP7_75t_L g2844 ( 
.A1(n_2641),
.A2(n_2596),
.B1(n_2681),
.B2(n_2678),
.Y(n_2844)
);

BUFx3_ASAP7_75t_L g2845 ( 
.A(n_2691),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2754),
.B(n_2535),
.Y(n_2846)
);

OAI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2585),
.A2(n_2641),
.B1(n_2657),
.B2(n_2592),
.Y(n_2847)
);

OAI21x1_ASAP7_75t_L g2848 ( 
.A1(n_2705),
.A2(n_2581),
.B(n_2579),
.Y(n_2848)
);

INVx6_ASAP7_75t_L g2849 ( 
.A(n_2615),
.Y(n_2849)
);

AND2x4_ASAP7_75t_L g2850 ( 
.A(n_2646),
.B(n_2383),
.Y(n_2850)
);

OAI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_2592),
.A2(n_2324),
.B1(n_2326),
.B2(n_2340),
.Y(n_2851)
);

INVxp33_ASAP7_75t_L g2852 ( 
.A(n_2655),
.Y(n_2852)
);

AOI22xp33_ASAP7_75t_L g2853 ( 
.A1(n_2637),
.A2(n_2570),
.B1(n_2575),
.B2(n_2467),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2607),
.Y(n_2854)
);

OAI22xp5_ASAP7_75t_L g2855 ( 
.A1(n_2592),
.A2(n_2423),
.B1(n_2377),
.B2(n_2371),
.Y(n_2855)
);

AND2x2_ASAP7_75t_SL g2856 ( 
.A(n_2677),
.B(n_2577),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2631),
.B(n_2458),
.Y(n_2857)
);

OAI22xp33_ASAP7_75t_L g2858 ( 
.A1(n_2657),
.A2(n_2423),
.B1(n_2377),
.B2(n_2371),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2752),
.B(n_2538),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2637),
.A2(n_2470),
.B1(n_2303),
.B2(n_2305),
.Y(n_2860)
);

OAI22xp33_ASAP7_75t_L g2861 ( 
.A1(n_2657),
.A2(n_2458),
.B1(n_2305),
.B2(n_2560),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2607),
.Y(n_2862)
);

INVx4_ASAP7_75t_SL g2863 ( 
.A(n_2686),
.Y(n_2863)
);

INVx2_ASAP7_75t_SL g2864 ( 
.A(n_2712),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2694),
.B(n_2538),
.Y(n_2865)
);

AOI22xp33_ASAP7_75t_L g2866 ( 
.A1(n_2689),
.A2(n_2307),
.B1(n_2567),
.B2(n_2560),
.Y(n_2866)
);

AOI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2663),
.A2(n_2567),
.B1(n_2555),
.B2(n_2486),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2631),
.B(n_2493),
.Y(n_2868)
);

OAI211xp5_ASAP7_75t_SL g2869 ( 
.A1(n_2651),
.A2(n_2383),
.B(n_2404),
.C(n_2555),
.Y(n_2869)
);

NOR2x1_ASAP7_75t_R g2870 ( 
.A(n_2722),
.B(n_2733),
.Y(n_2870)
);

AND2x4_ASAP7_75t_L g2871 ( 
.A(n_2690),
.B(n_2404),
.Y(n_2871)
);

OAI221xp5_ASAP7_75t_L g2872 ( 
.A1(n_2685),
.A2(n_2486),
.B1(n_2454),
.B2(n_2538),
.C(n_2554),
.Y(n_2872)
);

OAI22xp33_ASAP7_75t_L g2873 ( 
.A1(n_2702),
.A2(n_2554),
.B1(n_2480),
.B2(n_2464),
.Y(n_2873)
);

BUFx2_ASAP7_75t_L g2874 ( 
.A(n_2606),
.Y(n_2874)
);

OAI22xp33_ASAP7_75t_L g2875 ( 
.A1(n_2702),
.A2(n_2554),
.B1(n_2480),
.B2(n_2464),
.Y(n_2875)
);

NAND2xp33_ASAP7_75t_R g2876 ( 
.A(n_2709),
.B(n_405),
.Y(n_2876)
);

INVx3_ASAP7_75t_L g2877 ( 
.A(n_2662),
.Y(n_2877)
);

BUFx12f_ASAP7_75t_L g2878 ( 
.A(n_2718),
.Y(n_2878)
);

CKINVDCx20_ASAP7_75t_R g2879 ( 
.A(n_2684),
.Y(n_2879)
);

AOI21x1_ASAP7_75t_L g2880 ( 
.A1(n_2692),
.A2(n_2574),
.B(n_2552),
.Y(n_2880)
);

AND2x4_ASAP7_75t_L g2881 ( 
.A(n_2690),
.B(n_2549),
.Y(n_2881)
);

AOI22xp33_ASAP7_75t_SL g2882 ( 
.A1(n_2688),
.A2(n_2534),
.B1(n_2546),
.B2(n_2545),
.Y(n_2882)
);

INVx4_ASAP7_75t_L g2883 ( 
.A(n_2746),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2654),
.Y(n_2884)
);

OAI221xp5_ASAP7_75t_L g2885 ( 
.A1(n_2609),
.A2(n_2418),
.B1(n_2425),
.B2(n_2480),
.C(n_2549),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2661),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2661),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2736),
.Y(n_2888)
);

AOI22xp5_ASAP7_75t_L g2889 ( 
.A1(n_2770),
.A2(n_2548),
.B1(n_2418),
.B2(n_2425),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2726),
.B(n_2493),
.Y(n_2890)
);

NAND2x1p5_ASAP7_75t_L g2891 ( 
.A(n_2672),
.B(n_2418),
.Y(n_2891)
);

AOI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_2742),
.A2(n_2322),
.B(n_2381),
.Y(n_2892)
);

OAI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2710),
.A2(n_2492),
.B1(n_2495),
.B2(n_2515),
.Y(n_2893)
);

O2A1O1Ixp33_ASAP7_75t_SL g2894 ( 
.A1(n_2740),
.A2(n_2515),
.B(n_2495),
.C(n_2481),
.Y(n_2894)
);

AND2x2_ASAP7_75t_L g2895 ( 
.A(n_2698),
.B(n_406),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2688),
.B(n_2626),
.Y(n_2896)
);

AOI22xp5_ASAP7_75t_L g2897 ( 
.A1(n_2770),
.A2(n_2481),
.B1(n_2381),
.B2(n_409),
.Y(n_2897)
);

OAI22xp33_ASAP7_75t_L g2898 ( 
.A1(n_2710),
.A2(n_2381),
.B1(n_408),
.B2(n_409),
.Y(n_2898)
);

BUFx12f_ASAP7_75t_L g2899 ( 
.A(n_2721),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2639),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2653),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2764),
.Y(n_2902)
);

OAI22xp5_ASAP7_75t_L g2903 ( 
.A1(n_2758),
.A2(n_406),
.B1(n_408),
.B2(n_412),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2614),
.B(n_412),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2649),
.A2(n_2623),
.B1(n_2614),
.B2(n_2745),
.Y(n_2905)
);

HB1xp67_ASAP7_75t_L g2906 ( 
.A(n_2701),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2886),
.B(n_2887),
.Y(n_2907)
);

AOI22xp33_ASAP7_75t_L g2908 ( 
.A1(n_2811),
.A2(n_2649),
.B1(n_2737),
.B2(n_2706),
.Y(n_2908)
);

OAI22xp5_ASAP7_75t_L g2909 ( 
.A1(n_2811),
.A2(n_2758),
.B1(n_2762),
.B2(n_2737),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2846),
.B(n_2682),
.Y(n_2910)
);

AO21x2_ASAP7_75t_L g2911 ( 
.A1(n_2880),
.A2(n_2648),
.B(n_2768),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2776),
.Y(n_2912)
);

OAI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2810),
.A2(n_2814),
.B1(n_2804),
.B2(n_2798),
.Y(n_2913)
);

OAI22xp33_ASAP7_75t_L g2914 ( 
.A1(n_2814),
.A2(n_2674),
.B1(n_2746),
.B2(n_2751),
.Y(n_2914)
);

OAI22xp33_ASAP7_75t_L g2915 ( 
.A1(n_2876),
.A2(n_2674),
.B1(n_2746),
.B2(n_2751),
.Y(n_2915)
);

OAI22xp33_ASAP7_75t_L g2916 ( 
.A1(n_2787),
.A2(n_2751),
.B1(n_2742),
.B2(n_2759),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2788),
.B(n_2682),
.Y(n_2917)
);

AOI22xp33_ASAP7_75t_L g2918 ( 
.A1(n_2790),
.A2(n_2597),
.B1(n_2739),
.B2(n_2656),
.Y(n_2918)
);

AOI22xp5_ASAP7_75t_L g2919 ( 
.A1(n_2799),
.A2(n_2844),
.B1(n_2847),
.B2(n_2800),
.Y(n_2919)
);

AOI21xp33_ASAP7_75t_L g2920 ( 
.A1(n_2815),
.A2(n_2650),
.B(n_2620),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2774),
.A2(n_2602),
.B(n_2766),
.Y(n_2921)
);

BUFx2_ASAP7_75t_L g2922 ( 
.A(n_2789),
.Y(n_2922)
);

OAI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_2809),
.A2(n_2699),
.B1(n_2687),
.B2(n_2719),
.Y(n_2923)
);

AOI21xp5_ASAP7_75t_L g2924 ( 
.A1(n_2823),
.A2(n_2719),
.B(n_2711),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2831),
.Y(n_2925)
);

CKINVDCx5p33_ASAP7_75t_R g2926 ( 
.A(n_2791),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2781),
.Y(n_2927)
);

OR2x2_ASAP7_75t_L g2928 ( 
.A(n_2780),
.B(n_2744),
.Y(n_2928)
);

OAI22xp5_ASAP7_75t_L g2929 ( 
.A1(n_2820),
.A2(n_2838),
.B1(n_2860),
.B2(n_2827),
.Y(n_2929)
);

AOI221xp5_ASAP7_75t_L g2930 ( 
.A1(n_2805),
.A2(n_2666),
.B1(n_2665),
.B2(n_2759),
.C(n_2725),
.Y(n_2930)
);

OAI221xp5_ASAP7_75t_L g2931 ( 
.A1(n_2840),
.A2(n_2728),
.B1(n_2665),
.B2(n_2755),
.C(n_2679),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2784),
.Y(n_2932)
);

AOI22xp33_ASAP7_75t_L g2933 ( 
.A1(n_2786),
.A2(n_2679),
.B1(n_2636),
.B2(n_2738),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2830),
.B(n_2682),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2888),
.B(n_2660),
.Y(n_2935)
);

AOI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_2812),
.A2(n_2660),
.B1(n_2753),
.B2(n_2636),
.Y(n_2936)
);

AOI322xp5_ASAP7_75t_L g2937 ( 
.A1(n_2865),
.A2(n_2753),
.A3(n_2671),
.B1(n_2659),
.B2(n_2664),
.C1(n_2733),
.C2(n_419),
.Y(n_2937)
);

AOI221xp5_ASAP7_75t_L g2938 ( 
.A1(n_2778),
.A2(n_2714),
.B1(n_2594),
.B2(n_2723),
.C(n_2659),
.Y(n_2938)
);

OAI22xp33_ASAP7_75t_SL g2939 ( 
.A1(n_2849),
.A2(n_2864),
.B1(n_2874),
.B2(n_2789),
.Y(n_2939)
);

AOI21xp33_ASAP7_75t_L g2940 ( 
.A1(n_2896),
.A2(n_2763),
.B(n_2604),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2792),
.Y(n_2941)
);

INVx2_ASAP7_75t_SL g2942 ( 
.A(n_2821),
.Y(n_2942)
);

AOI22xp33_ASAP7_75t_SL g2943 ( 
.A1(n_2903),
.A2(n_2856),
.B1(n_2849),
.B2(n_2885),
.Y(n_2943)
);

OR2x2_ASAP7_75t_L g2944 ( 
.A(n_2782),
.B(n_2664),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2906),
.B(n_2608),
.Y(n_2945)
);

AOI221xp5_ASAP7_75t_L g2946 ( 
.A1(n_2884),
.A2(n_2731),
.B1(n_2750),
.B2(n_2708),
.C(n_2667),
.Y(n_2946)
);

OAI211xp5_ASAP7_75t_L g2947 ( 
.A1(n_2866),
.A2(n_2593),
.B(n_2734),
.C(n_2727),
.Y(n_2947)
);

NOR2xp33_ASAP7_75t_L g2948 ( 
.A(n_2801),
.B(n_2671),
.Y(n_2948)
);

OAI22xp33_ASAP7_75t_L g2949 ( 
.A1(n_2903),
.A2(n_2593),
.B1(n_2727),
.B2(n_2765),
.Y(n_2949)
);

AOI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2836),
.A2(n_2861),
.B(n_2858),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_2832),
.A2(n_2633),
.B1(n_2771),
.B2(n_2767),
.Y(n_2951)
);

A2O1A1Ixp33_ASAP7_75t_L g2952 ( 
.A1(n_2795),
.A2(n_2852),
.B(n_2889),
.C(n_2877),
.Y(n_2952)
);

AOI22xp33_ASAP7_75t_L g2953 ( 
.A1(n_2841),
.A2(n_2851),
.B1(n_2855),
.B2(n_2890),
.Y(n_2953)
);

AOI211xp5_ASAP7_75t_L g2954 ( 
.A1(n_2870),
.A2(n_2704),
.B(n_2582),
.C(n_2587),
.Y(n_2954)
);

AOI22xp33_ASAP7_75t_L g2955 ( 
.A1(n_2841),
.A2(n_2640),
.B1(n_2632),
.B2(n_2748),
.Y(n_2955)
);

AO22x1_ASAP7_75t_L g2956 ( 
.A1(n_2783),
.A2(n_2765),
.B1(n_2760),
.B2(n_2667),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2796),
.Y(n_2957)
);

AOI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_2824),
.A2(n_2748),
.B1(n_2732),
.B2(n_2765),
.Y(n_2958)
);

AOI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2838),
.A2(n_2748),
.B1(n_2605),
.B2(n_2599),
.Y(n_2959)
);

OAI222xp33_ASAP7_75t_L g2960 ( 
.A1(n_2783),
.A2(n_2905),
.B1(n_2889),
.B2(n_2897),
.C1(n_2893),
.C2(n_2807),
.Y(n_2960)
);

OAI21x1_ASAP7_75t_L g2961 ( 
.A1(n_2848),
.A2(n_2715),
.B(n_2697),
.Y(n_2961)
);

AND2x2_ASAP7_75t_L g2962 ( 
.A(n_2895),
.B(n_2624),
.Y(n_2962)
);

AND2x2_ASAP7_75t_L g2963 ( 
.A(n_2777),
.B(n_2624),
.Y(n_2963)
);

AOI222xp33_ASAP7_75t_L g2964 ( 
.A1(n_2863),
.A2(n_413),
.B1(n_414),
.B2(n_415),
.C1(n_416),
.C2(n_417),
.Y(n_2964)
);

NAND3xp33_ASAP7_75t_L g2965 ( 
.A(n_2902),
.B(n_2760),
.C(n_416),
.Y(n_2965)
);

INVx3_ASAP7_75t_L g2966 ( 
.A(n_2883),
.Y(n_2966)
);

OAI221xp5_ASAP7_75t_L g2967 ( 
.A1(n_2842),
.A2(n_2760),
.B1(n_417),
.B2(n_419),
.C(n_420),
.Y(n_2967)
);

AOI22xp33_ASAP7_75t_L g2968 ( 
.A1(n_2834),
.A2(n_2748),
.B1(n_2600),
.B2(n_2622),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2816),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_SL g2970 ( 
.A(n_2873),
.B(n_2703),
.Y(n_2970)
);

AOI222xp33_ASAP7_75t_L g2971 ( 
.A1(n_2863),
.A2(n_413),
.B1(n_420),
.B2(n_421),
.C1(n_422),
.C2(n_423),
.Y(n_2971)
);

OAI22xp5_ASAP7_75t_L g2972 ( 
.A1(n_2897),
.A2(n_2645),
.B1(n_2591),
.B2(n_423),
.Y(n_2972)
);

INVx4_ASAP7_75t_L g2973 ( 
.A(n_2826),
.Y(n_2973)
);

INVx5_ASAP7_75t_SL g2974 ( 
.A(n_2881),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2867),
.A2(n_421),
.B1(n_422),
.B2(n_424),
.Y(n_2975)
);

HB1xp67_ASAP7_75t_L g2976 ( 
.A(n_2818),
.Y(n_2976)
);

AOI22xp33_ASAP7_75t_L g2977 ( 
.A1(n_2828),
.A2(n_2696),
.B1(n_2695),
.B2(n_426),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2859),
.A2(n_424),
.B1(n_425),
.B2(n_426),
.Y(n_2978)
);

INVx6_ASAP7_75t_L g2979 ( 
.A(n_2775),
.Y(n_2979)
);

INVx5_ASAP7_75t_L g2980 ( 
.A(n_2878),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2835),
.Y(n_2981)
);

AOI22xp33_ASAP7_75t_L g2982 ( 
.A1(n_2854),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_2982)
);

AND2x4_ASAP7_75t_L g2983 ( 
.A(n_2794),
.B(n_429),
.Y(n_2983)
);

INVxp67_ASAP7_75t_L g2984 ( 
.A(n_2845),
.Y(n_2984)
);

AOI22xp33_ASAP7_75t_L g2985 ( 
.A1(n_2862),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_2985)
);

OAI22xp33_ASAP7_75t_SL g2986 ( 
.A1(n_2779),
.A2(n_431),
.B1(n_433),
.B2(n_434),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_2817),
.Y(n_2987)
);

OAI211xp5_ASAP7_75t_L g2988 ( 
.A1(n_2825),
.A2(n_433),
.B(n_434),
.C(n_436),
.Y(n_2988)
);

AND2x2_ASAP7_75t_L g2989 ( 
.A(n_2963),
.B(n_2868),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2910),
.B(n_2891),
.Y(n_2990)
);

OR2x2_ASAP7_75t_L g2991 ( 
.A(n_2925),
.B(n_2813),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2941),
.B(n_2843),
.Y(n_2992)
);

AND2x2_ASAP7_75t_L g2993 ( 
.A(n_2917),
.B(n_2934),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2981),
.Y(n_2994)
);

AOI22xp33_ASAP7_75t_L g2995 ( 
.A1(n_2913),
.A2(n_2919),
.B1(n_2929),
.B2(n_2916),
.Y(n_2995)
);

HB1xp67_ASAP7_75t_L g2996 ( 
.A(n_2976),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2912),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2907),
.B(n_2857),
.Y(n_2998)
);

AOI21xp5_ASAP7_75t_L g2999 ( 
.A1(n_2950),
.A2(n_2875),
.B(n_2894),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2962),
.B(n_2891),
.Y(n_3000)
);

INVx2_ASAP7_75t_SL g3001 ( 
.A(n_2922),
.Y(n_3001)
);

BUFx6f_ASAP7_75t_L g3002 ( 
.A(n_2961),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2957),
.Y(n_3003)
);

NOR2x1_ASAP7_75t_L g3004 ( 
.A(n_2973),
.B(n_2883),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2927),
.Y(n_3005)
);

INVx2_ASAP7_75t_SL g3006 ( 
.A(n_2979),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2932),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2969),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2953),
.B(n_2900),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2959),
.Y(n_3010)
);

INVx2_ASAP7_75t_SL g3011 ( 
.A(n_2979),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2947),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2911),
.Y(n_3013)
);

OR2x2_ASAP7_75t_L g3014 ( 
.A(n_2928),
.B(n_2785),
.Y(n_3014)
);

HB1xp67_ASAP7_75t_L g3015 ( 
.A(n_2944),
.Y(n_3015)
);

BUFx2_ASAP7_75t_L g3016 ( 
.A(n_2956),
.Y(n_3016)
);

AND2x4_ASAP7_75t_L g3017 ( 
.A(n_2924),
.B(n_2901),
.Y(n_3017)
);

NAND2xp33_ASAP7_75t_R g3018 ( 
.A(n_2987),
.B(n_2877),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2911),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2972),
.Y(n_3020)
);

OAI321xp33_ASAP7_75t_L g3021 ( 
.A1(n_2913),
.A2(n_2872),
.A3(n_2898),
.B1(n_2839),
.B2(n_2904),
.C(n_2853),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2972),
.Y(n_3022)
);

NOR2xp33_ASAP7_75t_L g3023 ( 
.A(n_2942),
.B(n_2779),
.Y(n_3023)
);

CKINVDCx5p33_ASAP7_75t_R g3024 ( 
.A(n_2926),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2966),
.Y(n_3025)
);

AND2x2_ASAP7_75t_L g3026 ( 
.A(n_2940),
.B(n_2892),
.Y(n_3026)
);

BUFx3_ASAP7_75t_L g3027 ( 
.A(n_2973),
.Y(n_3027)
);

INVxp67_ASAP7_75t_SL g3028 ( 
.A(n_2949),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2935),
.B(n_2822),
.Y(n_3029)
);

AND2x2_ASAP7_75t_L g3030 ( 
.A(n_2933),
.B(n_2822),
.Y(n_3030)
);

BUFx2_ASAP7_75t_SL g3031 ( 
.A(n_3027),
.Y(n_3031)
);

HB1xp67_ASAP7_75t_L g3032 ( 
.A(n_2996),
.Y(n_3032)
);

OAI221xp5_ASAP7_75t_L g3033 ( 
.A1(n_2995),
.A2(n_2943),
.B1(n_2952),
.B2(n_2929),
.C(n_2908),
.Y(n_3033)
);

INVx3_ASAP7_75t_L g3034 ( 
.A(n_3002),
.Y(n_3034)
);

OAI22xp5_ASAP7_75t_L g3035 ( 
.A1(n_3027),
.A2(n_2918),
.B1(n_2915),
.B2(n_2936),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_3008),
.Y(n_3036)
);

BUFx2_ASAP7_75t_L g3037 ( 
.A(n_3016),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_3008),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2997),
.Y(n_3039)
);

OAI22xp33_ASAP7_75t_L g3040 ( 
.A1(n_3027),
.A2(n_2914),
.B1(n_2980),
.B2(n_2909),
.Y(n_3040)
);

AND2x2_ASAP7_75t_L g3041 ( 
.A(n_3029),
.B(n_2989),
.Y(n_3041)
);

HB1xp67_ASAP7_75t_L g3042 ( 
.A(n_3001),
.Y(n_3042)
);

OAI22xp5_ASAP7_75t_L g3043 ( 
.A1(n_3004),
.A2(n_2909),
.B1(n_2923),
.B2(n_2983),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_3029),
.B(n_2970),
.Y(n_3044)
);

OAI211xp5_ASAP7_75t_L g3045 ( 
.A1(n_3028),
.A2(n_2964),
.B(n_2971),
.C(n_2937),
.Y(n_3045)
);

NOR2x2_ASAP7_75t_L g3046 ( 
.A(n_3018),
.B(n_2980),
.Y(n_3046)
);

OAI21x1_ASAP7_75t_L g3047 ( 
.A1(n_3013),
.A2(n_3019),
.B(n_3012),
.Y(n_3047)
);

AOI22xp33_ASAP7_75t_L g3048 ( 
.A1(n_3020),
.A2(n_2923),
.B1(n_2930),
.B2(n_2964),
.Y(n_3048)
);

AOI22xp5_ASAP7_75t_L g3049 ( 
.A1(n_3020),
.A2(n_2971),
.B1(n_2975),
.B2(n_2983),
.Y(n_3049)
);

OAI221xp5_ASAP7_75t_L g3050 ( 
.A1(n_3012),
.A2(n_3022),
.B1(n_2999),
.B2(n_3001),
.C(n_2920),
.Y(n_3050)
);

HB1xp67_ASAP7_75t_L g3051 ( 
.A(n_3015),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_3003),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_R g3053 ( 
.A(n_3024),
.B(n_2803),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_3003),
.Y(n_3054)
);

NAND2xp33_ASAP7_75t_SL g3055 ( 
.A(n_3016),
.B(n_2879),
.Y(n_3055)
);

OAI22xp33_ASAP7_75t_L g3056 ( 
.A1(n_3006),
.A2(n_2980),
.B1(n_2931),
.B2(n_2966),
.Y(n_3056)
);

NOR2xp33_ASAP7_75t_R g3057 ( 
.A(n_3006),
.B(n_2980),
.Y(n_3057)
);

BUFx3_ASAP7_75t_L g3058 ( 
.A(n_3011),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2989),
.B(n_2920),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_3009),
.B(n_2938),
.Y(n_3060)
);

AND2x4_ASAP7_75t_L g3061 ( 
.A(n_3017),
.B(n_2955),
.Y(n_3061)
);

OR2x2_ASAP7_75t_L g3062 ( 
.A(n_2991),
.B(n_2984),
.Y(n_3062)
);

AND2x2_ASAP7_75t_L g3063 ( 
.A(n_2993),
.B(n_2990),
.Y(n_3063)
);

AND2x2_ASAP7_75t_L g3064 ( 
.A(n_2993),
.B(n_2946),
.Y(n_3064)
);

OAI211xp5_ASAP7_75t_L g3065 ( 
.A1(n_3004),
.A2(n_2948),
.B(n_2954),
.C(n_2988),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2997),
.Y(n_3066)
);

OAI221xp5_ASAP7_75t_L g3067 ( 
.A1(n_3022),
.A2(n_2939),
.B1(n_2967),
.B2(n_2978),
.C(n_2975),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_R g3068 ( 
.A(n_3011),
.B(n_2773),
.Y(n_3068)
);

AOI22xp33_ASAP7_75t_L g3069 ( 
.A1(n_3009),
.A2(n_2965),
.B1(n_2945),
.B2(n_2794),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_3038),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_3038),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_3041),
.B(n_3044),
.Y(n_3072)
);

INVx3_ASAP7_75t_L g3073 ( 
.A(n_3034),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_3064),
.B(n_2994),
.Y(n_3074)
);

HB1xp67_ASAP7_75t_L g3075 ( 
.A(n_3051),
.Y(n_3075)
);

INVx2_ASAP7_75t_L g3076 ( 
.A(n_3036),
.Y(n_3076)
);

AND2x2_ASAP7_75t_L g3077 ( 
.A(n_3041),
.B(n_2990),
.Y(n_3077)
);

AND2x4_ASAP7_75t_L g3078 ( 
.A(n_3061),
.B(n_3017),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_3052),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_3044),
.B(n_3030),
.Y(n_3080)
);

HB1xp67_ASAP7_75t_L g3081 ( 
.A(n_3032),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_3064),
.B(n_2994),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_3059),
.B(n_3005),
.Y(n_3083)
);

INVxp67_ASAP7_75t_L g3084 ( 
.A(n_3047),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_3052),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_3063),
.B(n_3030),
.Y(n_3086)
);

AND2x2_ASAP7_75t_L g3087 ( 
.A(n_3063),
.B(n_3061),
.Y(n_3087)
);

CKINVDCx5p33_ASAP7_75t_R g3088 ( 
.A(n_3068),
.Y(n_3088)
);

AND2x4_ASAP7_75t_L g3089 ( 
.A(n_3061),
.B(n_3017),
.Y(n_3089)
);

INVx1_ASAP7_75t_SL g3090 ( 
.A(n_3046),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_3061),
.B(n_3026),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_3054),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_3054),
.Y(n_3093)
);

BUFx6f_ASAP7_75t_L g3094 ( 
.A(n_3034),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_3042),
.B(n_3037),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_3039),
.Y(n_3096)
);

AND2x2_ASAP7_75t_L g3097 ( 
.A(n_3037),
.B(n_3026),
.Y(n_3097)
);

INVxp67_ASAP7_75t_SL g3098 ( 
.A(n_3047),
.Y(n_3098)
);

OR2x2_ASAP7_75t_L g3099 ( 
.A(n_3062),
.B(n_2991),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3066),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_3083),
.B(n_3066),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_3091),
.B(n_3058),
.Y(n_3102)
);

INVxp67_ASAP7_75t_SL g3103 ( 
.A(n_3081),
.Y(n_3103)
);

OAI21x1_ASAP7_75t_L g3104 ( 
.A1(n_3073),
.A2(n_3034),
.B(n_3060),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_3083),
.B(n_3005),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_3096),
.Y(n_3106)
);

INVxp67_ASAP7_75t_SL g3107 ( 
.A(n_3081),
.Y(n_3107)
);

INVxp67_ASAP7_75t_SL g3108 ( 
.A(n_3075),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_3074),
.B(n_3007),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_3091),
.B(n_3058),
.Y(n_3110)
);

OR2x2_ASAP7_75t_L g3111 ( 
.A(n_3074),
.B(n_3062),
.Y(n_3111)
);

AND2x2_ASAP7_75t_L g3112 ( 
.A(n_3091),
.B(n_3058),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_3076),
.Y(n_3113)
);

INVx1_ASAP7_75t_SL g3114 ( 
.A(n_3075),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_3097),
.B(n_3087),
.Y(n_3115)
);

AND2x2_ASAP7_75t_L g3116 ( 
.A(n_3097),
.B(n_3010),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_3082),
.B(n_3007),
.Y(n_3117)
);

OR2x2_ASAP7_75t_L g3118 ( 
.A(n_3082),
.B(n_3014),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_3076),
.Y(n_3119)
);

OAI21xp5_ASAP7_75t_SL g3120 ( 
.A1(n_3090),
.A2(n_3043),
.B(n_3045),
.Y(n_3120)
);

INVx2_ASAP7_75t_SL g3121 ( 
.A(n_3090),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_3108),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_3108),
.Y(n_3123)
);

INVx3_ASAP7_75t_SL g3124 ( 
.A(n_3121),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_3120),
.B(n_3097),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_3120),
.B(n_3080),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_3116),
.B(n_3080),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_3103),
.Y(n_3128)
);

AND2x2_ASAP7_75t_L g3129 ( 
.A(n_3121),
.B(n_3115),
.Y(n_3129)
);

OAI221xp5_ASAP7_75t_L g3130 ( 
.A1(n_3107),
.A2(n_3055),
.B1(n_3033),
.B2(n_3050),
.C(n_3043),
.Y(n_3130)
);

NAND5xp2_ASAP7_75t_SL g3131 ( 
.A(n_3102),
.B(n_3088),
.C(n_3065),
.D(n_3048),
.E(n_3049),
.Y(n_3131)
);

AND2x2_ASAP7_75t_L g3132 ( 
.A(n_3115),
.B(n_3087),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_3111),
.Y(n_3133)
);

OR2x2_ASAP7_75t_L g3134 ( 
.A(n_3118),
.B(n_3099),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_3111),
.Y(n_3135)
);

AND2x2_ASAP7_75t_L g3136 ( 
.A(n_3116),
.B(n_3087),
.Y(n_3136)
);

HB1xp67_ASAP7_75t_L g3137 ( 
.A(n_3114),
.Y(n_3137)
);

AND2x4_ASAP7_75t_L g3138 ( 
.A(n_3114),
.B(n_3078),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_3109),
.B(n_3080),
.Y(n_3139)
);

NOR2x1_ASAP7_75t_L g3140 ( 
.A(n_3102),
.B(n_3031),
.Y(n_3140)
);

NOR2x1_ASAP7_75t_L g3141 ( 
.A(n_3110),
.B(n_3031),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3118),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_3113),
.Y(n_3143)
);

OR2x2_ASAP7_75t_L g3144 ( 
.A(n_3109),
.B(n_3099),
.Y(n_3144)
);

INVxp33_ASAP7_75t_L g3145 ( 
.A(n_3110),
.Y(n_3145)
);

OR2x2_ASAP7_75t_L g3146 ( 
.A(n_3117),
.B(n_3095),
.Y(n_3146)
);

A2O1A1Ixp33_ASAP7_75t_L g3147 ( 
.A1(n_3130),
.A2(n_3140),
.B(n_3141),
.C(n_3125),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_3137),
.Y(n_3148)
);

AOI21xp33_ASAP7_75t_L g3149 ( 
.A1(n_3137),
.A2(n_3084),
.B(n_3098),
.Y(n_3149)
);

OAI22xp5_ASAP7_75t_L g3150 ( 
.A1(n_3126),
.A2(n_3112),
.B1(n_3089),
.B2(n_3078),
.Y(n_3150)
);

INVx1_ASAP7_75t_SL g3151 ( 
.A(n_3124),
.Y(n_3151)
);

OA21x2_ASAP7_75t_L g3152 ( 
.A1(n_3122),
.A2(n_3084),
.B(n_3104),
.Y(n_3152)
);

OAI22xp5_ASAP7_75t_L g3153 ( 
.A1(n_3145),
.A2(n_3112),
.B1(n_3078),
.B2(n_3089),
.Y(n_3153)
);

INVxp67_ASAP7_75t_L g3154 ( 
.A(n_3123),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_3124),
.B(n_3117),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3128),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_3133),
.B(n_3105),
.Y(n_3157)
);

AOI31xp33_ASAP7_75t_SL g3158 ( 
.A1(n_3131),
.A2(n_3023),
.A3(n_3069),
.B(n_3053),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_3129),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3134),
.Y(n_3160)
);

INVxp67_ASAP7_75t_L g3161 ( 
.A(n_3135),
.Y(n_3161)
);

AOI22xp33_ASAP7_75t_L g3162 ( 
.A1(n_3138),
.A2(n_3035),
.B1(n_3078),
.B2(n_3089),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_3145),
.B(n_2806),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_3132),
.B(n_3095),
.Y(n_3164)
);

OAI221xp5_ASAP7_75t_L g3165 ( 
.A1(n_3142),
.A2(n_3035),
.B1(n_3098),
.B2(n_3049),
.C(n_3067),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_L g3166 ( 
.A(n_3144),
.B(n_3105),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_3148),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_3151),
.Y(n_3168)
);

AOI22xp5_ASAP7_75t_L g3169 ( 
.A1(n_3165),
.A2(n_3138),
.B1(n_3132),
.B2(n_3089),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_3159),
.B(n_3136),
.Y(n_3170)
);

AOI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_3162),
.A2(n_3138),
.B1(n_3040),
.B2(n_3146),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_3160),
.B(n_3136),
.Y(n_3172)
);

OAI21xp5_ASAP7_75t_L g3173 ( 
.A1(n_3147),
.A2(n_3104),
.B(n_3127),
.Y(n_3173)
);

OAI21xp33_ASAP7_75t_L g3174 ( 
.A1(n_3155),
.A2(n_3139),
.B(n_3143),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3156),
.Y(n_3175)
);

OAI21xp5_ASAP7_75t_L g3176 ( 
.A1(n_3154),
.A2(n_2986),
.B(n_3104),
.Y(n_3176)
);

OAI22xp33_ASAP7_75t_L g3177 ( 
.A1(n_3153),
.A2(n_3056),
.B1(n_3073),
.B2(n_3143),
.Y(n_3177)
);

AOI21xp33_ASAP7_75t_SL g3178 ( 
.A1(n_3154),
.A2(n_2833),
.B(n_3101),
.Y(n_3178)
);

OR2x2_ASAP7_75t_L g3179 ( 
.A(n_3161),
.B(n_3101),
.Y(n_3179)
);

NAND3xp33_ASAP7_75t_L g3180 ( 
.A(n_3149),
.B(n_3094),
.C(n_2985),
.Y(n_3180)
);

AOI32xp33_ASAP7_75t_L g3181 ( 
.A1(n_3163),
.A2(n_3086),
.A3(n_3073),
.B1(n_3072),
.B2(n_3021),
.Y(n_3181)
);

AOI221xp5_ASAP7_75t_L g3182 ( 
.A1(n_3161),
.A2(n_2960),
.B1(n_3119),
.B2(n_3113),
.C(n_3086),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_3166),
.B(n_3086),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_3168),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3172),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_3167),
.B(n_3157),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_3175),
.B(n_3164),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_3170),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_3171),
.B(n_3150),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_3179),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_SL g3191 ( 
.A(n_3181),
.B(n_3158),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_3180),
.Y(n_3192)
);

INVxp67_ASAP7_75t_L g3193 ( 
.A(n_3169),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3174),
.Y(n_3194)
);

OR2x2_ASAP7_75t_L g3195 ( 
.A(n_3183),
.B(n_3152),
.Y(n_3195)
);

INVxp67_ASAP7_75t_L g3196 ( 
.A(n_3176),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_3177),
.B(n_3057),
.Y(n_3197)
);

AOI22xp33_ASAP7_75t_SL g3198 ( 
.A1(n_3176),
.A2(n_3152),
.B1(n_3094),
.B2(n_3073),
.Y(n_3198)
);

BUFx6f_ASAP7_75t_L g3199 ( 
.A(n_3184),
.Y(n_3199)
);

AND2x2_ASAP7_75t_L g3200 ( 
.A(n_3188),
.B(n_3178),
.Y(n_3200)
);

AO22x2_ASAP7_75t_L g3201 ( 
.A1(n_3185),
.A2(n_3173),
.B1(n_3182),
.B2(n_3119),
.Y(n_3201)
);

OAI21xp5_ASAP7_75t_L g3202 ( 
.A1(n_3196),
.A2(n_3191),
.B(n_3193),
.Y(n_3202)
);

NOR3xp33_ASAP7_75t_L g3203 ( 
.A(n_3194),
.B(n_2869),
.C(n_3034),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_3189),
.B(n_3113),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3192),
.B(n_3119),
.Y(n_3205)
);

OAI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3197),
.A2(n_3072),
.B1(n_3106),
.B2(n_3094),
.Y(n_3206)
);

OR2x2_ASAP7_75t_L g3207 ( 
.A(n_3187),
.B(n_3077),
.Y(n_3207)
);

XNOR2x2_ASAP7_75t_L g3208 ( 
.A(n_3186),
.B(n_3014),
.Y(n_3208)
);

NAND3xp33_ASAP7_75t_SL g3209 ( 
.A(n_3198),
.B(n_2982),
.C(n_2826),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_3190),
.B(n_3106),
.Y(n_3210)
);

AO221x1_ASAP7_75t_L g3211 ( 
.A1(n_3199),
.A2(n_3187),
.B1(n_3186),
.B2(n_3195),
.C(n_3094),
.Y(n_3211)
);

NOR2x1_ASAP7_75t_L g3212 ( 
.A(n_3202),
.B(n_3094),
.Y(n_3212)
);

NAND5xp2_ASAP7_75t_L g3213 ( 
.A(n_3200),
.B(n_2839),
.C(n_2958),
.D(n_2882),
.E(n_3010),
.Y(n_3213)
);

AOI221xp5_ASAP7_75t_L g3214 ( 
.A1(n_3204),
.A2(n_3094),
.B1(n_3019),
.B2(n_3013),
.C(n_3100),
.Y(n_3214)
);

OAI222xp33_ASAP7_75t_L g3215 ( 
.A1(n_3206),
.A2(n_3077),
.B1(n_3025),
.B2(n_3100),
.C1(n_2992),
.C2(n_2797),
.Y(n_3215)
);

OAI221xp5_ASAP7_75t_L g3216 ( 
.A1(n_3209),
.A2(n_3094),
.B1(n_2977),
.B2(n_2951),
.C(n_2793),
.Y(n_3216)
);

A2O1A1Ixp33_ASAP7_75t_L g3217 ( 
.A1(n_3205),
.A2(n_2921),
.B(n_2808),
.C(n_2802),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_SL g3218 ( 
.A(n_3203),
.B(n_3002),
.Y(n_3218)
);

INVx2_ASAP7_75t_SL g3219 ( 
.A(n_3210),
.Y(n_3219)
);

XNOR2xp5_ASAP7_75t_L g3220 ( 
.A(n_3208),
.B(n_436),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3220),
.Y(n_3221)
);

CKINVDCx16_ASAP7_75t_R g3222 ( 
.A(n_3219),
.Y(n_3222)
);

AOI22xp5_ASAP7_75t_L g3223 ( 
.A1(n_3211),
.A2(n_3201),
.B1(n_3207),
.B2(n_2899),
.Y(n_3223)
);

A2O1A1Ixp33_ASAP7_75t_L g3224 ( 
.A1(n_3212),
.A2(n_2819),
.B(n_3025),
.C(n_3071),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3222),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_3223),
.B(n_3217),
.Y(n_3226)
);

AND2x4_ASAP7_75t_L g3227 ( 
.A(n_3221),
.B(n_3218),
.Y(n_3227)
);

AOI21xp33_ASAP7_75t_SL g3228 ( 
.A1(n_3224),
.A2(n_3216),
.B(n_3213),
.Y(n_3228)
);

BUFx24_ASAP7_75t_SL g3229 ( 
.A(n_3223),
.Y(n_3229)
);

XNOR2xp5_ASAP7_75t_L g3230 ( 
.A(n_3229),
.B(n_3214),
.Y(n_3230)
);

OAI221xp5_ASAP7_75t_L g3231 ( 
.A1(n_3225),
.A2(n_3215),
.B1(n_2998),
.B2(n_2829),
.C(n_2837),
.Y(n_3231)
);

NAND2xp33_ASAP7_75t_L g3232 ( 
.A(n_3226),
.B(n_3002),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3230),
.B(n_3227),
.Y(n_3233)
);

INVxp33_ASAP7_75t_SL g3234 ( 
.A(n_3232),
.Y(n_3234)
);

AND2x4_ASAP7_75t_L g3235 ( 
.A(n_3231),
.B(n_3228),
.Y(n_3235)
);

OA22x2_ASAP7_75t_L g3236 ( 
.A1(n_3233),
.A2(n_3085),
.B1(n_3093),
.B2(n_3079),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_SL g3237 ( 
.A(n_3236),
.B(n_3235),
.Y(n_3237)
);

HB1xp67_ASAP7_75t_L g3238 ( 
.A(n_3237),
.Y(n_3238)
);

OAI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_3238),
.A2(n_3234),
.B(n_3092),
.Y(n_3239)
);

INVxp67_ASAP7_75t_L g3240 ( 
.A(n_3239),
.Y(n_3240)
);

AOI322xp5_ASAP7_75t_L g3241 ( 
.A1(n_3240),
.A2(n_3079),
.A3(n_3092),
.B1(n_3093),
.B2(n_3085),
.C1(n_3071),
.C2(n_3070),
.Y(n_3241)
);

OAI221xp5_ASAP7_75t_R g3242 ( 
.A1(n_3241),
.A2(n_2968),
.B1(n_438),
.B2(n_437),
.C(n_2974),
.Y(n_3242)
);

AOI211xp5_ASAP7_75t_L g3243 ( 
.A1(n_3242),
.A2(n_2850),
.B(n_2871),
.C(n_3000),
.Y(n_3243)
);


endmodule