module fake_netlist_6_3400_n_186 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_186);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_186;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_145;
wire n_92;
wire n_42;
wire n_133;
wire n_96;
wire n_160;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_1),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

OR2x6_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2x1p5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_34),
.B(n_2),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_3),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

AND3x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_5),
.C(n_6),
.Y(n_68)
);

CKINVDCx6p67_ASAP7_75t_R g69 ( 
.A(n_33),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_5),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g76 ( 
.A(n_51),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_53),
.C(n_52),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

O2A1O1Ixp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_42),
.B(n_41),
.C(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_46),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_44),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_35),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_72),
.B(n_65),
.C(n_76),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_78),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_69),
.Y(n_97)
);

AO31x2_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_72),
.A3(n_65),
.B(n_73),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_76),
.B(n_74),
.C(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_60),
.B1(n_64),
.B2(n_63),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_60),
.B(n_62),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_60),
.B(n_62),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_93),
.B(n_81),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_90),
.B(n_82),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_93),
.Y(n_107)
);

O2A1O1Ixp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_75),
.B(n_70),
.C(n_73),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_85),
.B(n_81),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_77),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_89),
.Y(n_111)
);

AOI21x1_ASAP7_75t_SL g112 ( 
.A1(n_103),
.A2(n_60),
.B(n_68),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_98),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_96),
.B(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_119),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_110),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_110),
.Y(n_133)
);

NOR2xp67_ASAP7_75t_SL g134 ( 
.A(n_123),
.B(n_117),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_97),
.B1(n_100),
.B2(n_60),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_128),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_68),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_37),
.A3(n_71),
.B1(n_56),
.B2(n_89),
.Y(n_142)
);

NOR4xp25_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_94),
.C(n_71),
.D(n_70),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

AOI211xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_69),
.B(n_79),
.C(n_70),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_133),
.B(n_116),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_139),
.Y(n_147)
);

OAI211xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_67),
.B(n_132),
.C(n_69),
.Y(n_148)
);

AOI211x1_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_140),
.B(n_142),
.C(n_67),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_101),
.B(n_102),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_129),
.B1(n_136),
.B2(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_136),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_129),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_133),
.B(n_109),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_134),
.C(n_103),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_98),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_147),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_61),
.C(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_61),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_151),
.A2(n_112),
.B(n_75),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_98),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_75),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

AND3x4_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_149),
.C(n_9),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_150),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_154),
.C(n_108),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_109),
.Y(n_169)
);

NAND4xp75_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_108),
.C(n_10),
.D(n_11),
.Y(n_170)
);

AND3x2_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_8),
.C(n_12),
.Y(n_171)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_26),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_161),
.B1(n_156),
.B2(n_92),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_112),
.C(n_81),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_8),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_19),
.C2(n_20),
.Y(n_175)
);

OAI211xp5_ASAP7_75t_SL g176 ( 
.A1(n_165),
.A2(n_13),
.B(n_14),
.C(n_85),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_85),
.B1(n_22),
.B2(n_82),
.C(n_90),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_82),
.A3(n_90),
.B1(n_92),
.B2(n_96),
.C1(n_169),
.C2(n_174),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_166),
.B1(n_173),
.B2(n_170),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_181),
.A2(n_176),
.B1(n_178),
.B2(n_90),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_96),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_181),
.Y(n_185)
);

AOI22x1_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_180),
.B1(n_183),
.B2(n_92),
.Y(n_186)
);


endmodule