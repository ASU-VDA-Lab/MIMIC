module fake_aes_5603_n_469 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_469);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_469;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_141;
wire n_119;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g62 ( .A(n_59), .Y(n_62) );
INVxp67_ASAP7_75t_SL g63 ( .A(n_6), .Y(n_63) );
BUFx3_ASAP7_75t_L g64 ( .A(n_48), .Y(n_64) );
INVxp67_ASAP7_75t_L g65 ( .A(n_49), .Y(n_65) );
HB1xp67_ASAP7_75t_L g66 ( .A(n_21), .Y(n_66) );
CKINVDCx5p33_ASAP7_75t_R g67 ( .A(n_50), .Y(n_67) );
CKINVDCx20_ASAP7_75t_R g68 ( .A(n_41), .Y(n_68) );
INVxp67_ASAP7_75t_SL g69 ( .A(n_4), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_37), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_20), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_36), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_8), .Y(n_73) );
HB1xp67_ASAP7_75t_L g74 ( .A(n_32), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_2), .Y(n_75) );
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_40), .Y(n_76) );
INVxp67_ASAP7_75t_SL g77 ( .A(n_53), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_26), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_28), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_51), .Y(n_80) );
CKINVDCx14_ASAP7_75t_R g81 ( .A(n_14), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_46), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_61), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_0), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_38), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_45), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_54), .Y(n_87) );
CKINVDCx14_ASAP7_75t_R g88 ( .A(n_9), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_35), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_5), .Y(n_91) );
INVxp33_ASAP7_75t_L g92 ( .A(n_8), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_56), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_58), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_42), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_39), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_55), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_0), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_68), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_76), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_81), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_88), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_62), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_64), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_64), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_62), .Y(n_106) );
NOR2xp33_ASAP7_75t_R g107 ( .A(n_67), .B(n_27), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_91), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_91), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_66), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_92), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_64), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_80), .Y(n_113) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_70), .A2(n_25), .B(n_60), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_71), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_85), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_74), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_71), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_72), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_115), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_111), .B(n_65), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_104), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_114), .Y(n_125) );
OR2x2_ASAP7_75t_L g126 ( .A(n_108), .B(n_63), .Y(n_126) );
NOR2x1p5_ASAP7_75t_L g127 ( .A(n_109), .B(n_63), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_104), .Y(n_128) );
NAND3xp33_ASAP7_75t_L g129 ( .A(n_103), .B(n_98), .C(n_73), .Y(n_129) );
NOR2x1p5_ASAP7_75t_L g130 ( .A(n_99), .B(n_69), .Y(n_130) );
BUFx3_ASAP7_75t_L g131 ( .A(n_105), .Y(n_131) );
OAI221xp5_ASAP7_75t_L g132 ( .A1(n_103), .A2(n_69), .B1(n_84), .B2(n_98), .C(n_73), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_115), .Y(n_133) );
AO22x2_ASAP7_75t_L g134 ( .A1(n_106), .A2(n_83), .B1(n_72), .B2(n_89), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_110), .A2(n_75), .B1(n_84), .B2(n_65), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_115), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_106), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_100), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_105), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_104), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_117), .B(n_96), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_105), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_117), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_120), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_120), .B(n_75), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_131), .Y(n_148) );
INVx4_ASAP7_75t_L g149 ( .A(n_147), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_147), .B(n_113), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_147), .B(n_121), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_137), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_137), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_147), .B(n_121), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_134), .A2(n_104), .B1(n_112), .B2(n_83), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_140), .B(n_118), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_141), .B(n_101), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_141), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
INVx5_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_128), .Y(n_164) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_145), .A2(n_114), .B(n_90), .Y(n_165) );
INVx6_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_146), .B(n_102), .Y(n_168) );
AND2x6_ASAP7_75t_SL g169 ( .A(n_123), .B(n_78), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_138), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_122), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
INVx3_ASAP7_75t_SL g177 ( .A(n_134), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_122), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_134), .A2(n_119), .B1(n_96), .B2(n_79), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_126), .B(n_97), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_152), .A2(n_139), .B(n_131), .Y(n_181) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_173), .Y(n_182) );
OAI222xp33_ASAP7_75t_L g183 ( .A1(n_179), .A2(n_135), .B1(n_132), .B2(n_126), .C1(n_143), .C2(n_136), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_149), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_177), .A2(n_127), .B1(n_130), .B2(n_133), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_152), .A2(n_131), .B(n_139), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_149), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
BUFx5_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_171), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_151), .B(n_127), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_149), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_177), .A2(n_130), .B1(n_129), .B2(n_136), .Y(n_193) );
BUFx4f_ASAP7_75t_L g194 ( .A(n_177), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_174), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_153), .Y(n_196) );
OAI21xp33_ASAP7_75t_L g197 ( .A1(n_179), .A2(n_133), .B(n_139), .Y(n_197) );
INVx2_ASAP7_75t_SL g198 ( .A(n_149), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_148), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_173), .A2(n_144), .B1(n_77), .B2(n_125), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_151), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_151), .A2(n_154), .B1(n_161), .B2(n_160), .Y(n_202) );
O2A1O1Ixp5_ASAP7_75t_L g203 ( .A1(n_158), .A2(n_144), .B(n_142), .C(n_90), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_154), .A2(n_125), .B1(n_94), .B2(n_89), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_169), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_174), .Y(n_206) );
OR2x2_ASAP7_75t_L g207 ( .A(n_158), .B(n_1), .Y(n_207) );
INVxp67_ASAP7_75t_L g208 ( .A(n_180), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_154), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_154), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_157), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_159), .B(n_168), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_150), .A2(n_78), .B(n_79), .C(n_82), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_203), .A2(n_170), .B(n_161), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_196), .A2(n_165), .B(n_160), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_212), .B(n_157), .Y(n_216) );
NAND3xp33_ASAP7_75t_SL g217 ( .A(n_205), .B(n_155), .C(n_107), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_202), .B(n_170), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_189), .Y(n_219) );
HB1xp67_ASAP7_75t_SL g220 ( .A(n_190), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_210), .A2(n_159), .B1(n_168), .B2(n_178), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_210), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_194), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_202), .A2(n_178), .B1(n_175), .B2(n_166), .Y(n_224) );
AOI221xp5_ASAP7_75t_L g225 ( .A1(n_183), .A2(n_155), .B1(n_175), .B2(n_82), .C(n_94), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_211), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_196), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_208), .B(n_169), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_189), .B(n_178), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_189), .B(n_188), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_189), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_189), .B(n_178), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_201), .A2(n_166), .B1(n_148), .B2(n_162), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_189), .B(n_162), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_209), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_182), .B(n_162), .Y(n_236) );
OAI221xp5_ASAP7_75t_L g237 ( .A1(n_207), .A2(n_86), .B1(n_87), .B2(n_93), .C(n_95), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_191), .B(n_162), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_185), .B(n_162), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_205), .A2(n_166), .B1(n_148), .B2(n_162), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_220), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_228), .A2(n_197), .B1(n_193), .B2(n_194), .Y(n_242) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_215), .A2(n_165), .B(n_186), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_216), .B(n_184), .Y(n_244) );
AOI221xp5_ASAP7_75t_L g245 ( .A1(n_216), .A2(n_213), .B1(n_190), .B2(n_184), .C(n_204), .Y(n_245) );
OAI22xp33_ASAP7_75t_L g246 ( .A1(n_237), .A2(n_200), .B1(n_198), .B2(n_187), .Y(n_246) );
OAI22xp33_ASAP7_75t_L g247 ( .A1(n_237), .A2(n_198), .B1(n_187), .B2(n_184), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_218), .A2(n_192), .B1(n_199), .B2(n_166), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_218), .A2(n_192), .B1(n_199), .B2(n_166), .Y(n_249) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_215), .A2(n_165), .B(n_181), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_227), .B(n_195), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_227), .Y(n_252) );
AOI21xp33_ASAP7_75t_L g253 ( .A1(n_239), .A2(n_104), .B(n_112), .Y(n_253) );
AOI21xp33_ASAP7_75t_L g254 ( .A1(n_219), .A2(n_104), .B(n_112), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_226), .B(n_162), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_219), .B(n_195), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_226), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_219), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_223), .B(n_174), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_214), .A2(n_114), .B(n_142), .Y(n_260) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_214), .A2(n_86), .B(n_87), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_235), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_220), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_247), .A2(n_221), .B1(n_225), .B2(n_217), .Y(n_264) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_253), .A2(n_225), .B(n_230), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_252), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_257), .B(n_235), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_257), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_252), .B(n_229), .Y(n_269) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_251), .Y(n_270) );
OAI21xp33_ASAP7_75t_L g271 ( .A1(n_242), .A2(n_217), .B(n_224), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_258), .B(n_231), .Y(n_272) );
INVx4_ASAP7_75t_L g273 ( .A(n_251), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_245), .A2(n_223), .B1(n_238), .B2(n_222), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_262), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_262), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_243), .Y(n_277) );
OAI221xp5_ASAP7_75t_L g278 ( .A1(n_245), .A2(n_240), .B1(n_230), .B2(n_223), .C(n_234), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_246), .A2(n_223), .B1(n_222), .B2(n_236), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_261), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_244), .B(n_231), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_258), .B(n_261), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_244), .A2(n_229), .B1(n_236), .B2(n_232), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_258), .B(n_231), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_263), .A2(n_229), .B1(n_232), .B2(n_234), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_266), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_266), .Y(n_287) );
OAI33xp33_ASAP7_75t_L g288 ( .A1(n_268), .A2(n_263), .A3(n_241), .B1(n_95), .B2(n_93), .B3(n_255), .Y(n_288) );
AOI21xp5_ASAP7_75t_SL g289 ( .A1(n_265), .A2(n_261), .B(n_259), .Y(n_289) );
AND2x2_ASAP7_75t_SL g290 ( .A(n_273), .B(n_261), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_266), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_275), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_275), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_276), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_270), .B(n_261), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_273), .B(n_255), .Y(n_297) );
INVxp67_ASAP7_75t_SL g298 ( .A(n_282), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_276), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_269), .B(n_248), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_273), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_269), .B(n_249), .Y(n_302) );
INVxp67_ASAP7_75t_SL g303 ( .A(n_282), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_282), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_273), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_277), .Y(n_306) );
NAND4xp25_ASAP7_75t_L g307 ( .A(n_271), .B(n_93), .C(n_95), .D(n_253), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_281), .B(n_250), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_272), .B(n_250), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_267), .B(n_250), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_277), .B(n_250), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_280), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_305), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_305), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_304), .B(n_277), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_292), .B(n_280), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_304), .B(n_272), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_306), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_298), .B(n_272), .Y(n_319) );
NOR3xp33_ASAP7_75t_SL g320 ( .A(n_288), .B(n_307), .C(n_271), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_303), .B(n_283), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_301), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_306), .Y(n_323) );
NAND2x1_ASAP7_75t_L g324 ( .A(n_287), .B(n_267), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_292), .B(n_265), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_286), .Y(n_326) );
NOR2x1p5_ASAP7_75t_L g327 ( .A(n_296), .B(n_281), .Y(n_327) );
NAND3xp33_ASAP7_75t_L g328 ( .A(n_289), .B(n_274), .C(n_264), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_309), .B(n_283), .Y(n_329) );
NOR3xp33_ASAP7_75t_L g330 ( .A(n_293), .B(n_278), .C(n_284), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_309), .B(n_265), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_294), .B(n_265), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_286), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_287), .Y(n_335) );
NOR2x1_ASAP7_75t_SL g336 ( .A(n_297), .B(n_284), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_312), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_300), .A2(n_278), .B1(n_285), .B2(n_279), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_312), .B(n_265), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_311), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_294), .Y(n_341) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_297), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_308), .B(n_243), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g344 ( .A1(n_289), .A2(n_254), .B(n_112), .C(n_256), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_295), .B(n_243), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_299), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_299), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_310), .B(n_112), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_291), .B(n_112), .Y(n_349) );
NAND3xp33_ASAP7_75t_L g350 ( .A(n_290), .B(n_254), .C(n_114), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_291), .B(n_260), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_308), .B(n_260), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_344), .B(n_290), .C(n_302), .Y(n_354) );
OAI221xp5_ASAP7_75t_SL g355 ( .A1(n_338), .A2(n_290), .B1(n_233), .B2(n_4), .C(n_5), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_342), .B(n_311), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_344), .B(n_311), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_319), .B(n_2), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_328), .A2(n_125), .B1(n_260), .B2(n_174), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_332), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_327), .A2(n_125), .B1(n_6), .B2(n_7), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_353), .B(n_3), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_327), .B(n_10), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_330), .A2(n_174), .B1(n_206), .B2(n_195), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_322), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g366 ( .A1(n_336), .A2(n_206), .B1(n_195), .B2(n_13), .Y(n_366) );
INVxp67_ASAP7_75t_L g367 ( .A(n_336), .Y(n_367) );
OAI21xp33_ASAP7_75t_L g368 ( .A1(n_320), .A2(n_11), .B(n_12), .Y(n_368) );
OAI322xp33_ASAP7_75t_SL g369 ( .A1(n_341), .A2(n_347), .A3(n_346), .B1(n_333), .B2(n_325), .C1(n_316), .C2(n_337), .Y(n_369) );
OAI21xp33_ASAP7_75t_L g370 ( .A1(n_320), .A2(n_11), .B(n_12), .Y(n_370) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_324), .B(n_13), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_313), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_321), .B(n_15), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_313), .B(n_15), .Y(n_375) );
AOI21xp33_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_16), .B(n_17), .Y(n_376) );
NAND2x1_ASAP7_75t_L g377 ( .A(n_335), .B(n_206), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_321), .B(n_17), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_314), .A2(n_18), .B1(n_19), .B2(n_174), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_314), .A2(n_18), .B1(n_19), .B2(n_176), .Y(n_380) );
AOI33xp33_ASAP7_75t_L g381 ( .A1(n_329), .A2(n_176), .A3(n_172), .B1(n_167), .B2(n_164), .B3(n_163), .Y(n_381) );
OAI21xp33_ASAP7_75t_L g382 ( .A1(n_331), .A2(n_176), .B(n_172), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_317), .B(n_22), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_348), .A2(n_167), .B(n_164), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_318), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_337), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_337), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_339), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_340), .B(n_23), .Y(n_389) );
A2O1A1Ixp33_ASAP7_75t_L g390 ( .A1(n_368), .A2(n_350), .B(n_343), .C(n_316), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_357), .A2(n_350), .B(n_352), .Y(n_391) );
OAI21xp33_ASAP7_75t_SL g392 ( .A1(n_367), .A2(n_325), .B(n_333), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_375), .B(n_343), .Y(n_393) );
NOR3xp33_ASAP7_75t_SL g394 ( .A(n_370), .B(n_352), .C(n_345), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_373), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_388), .B(n_315), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_365), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_360), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_375), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_356), .B(n_351), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_386), .Y(n_401) );
NOR3xp33_ASAP7_75t_L g402 ( .A(n_361), .B(n_349), .C(n_318), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_372), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_374), .B(n_323), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_387), .Y(n_405) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_371), .B(n_349), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_369), .A2(n_323), .B1(n_326), .B2(n_334), .C(n_164), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_372), .B(n_334), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_358), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_385), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_362), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_363), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_383), .B(n_24), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_377), .Y(n_414) );
INVxp67_ASAP7_75t_L g415 ( .A(n_378), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_354), .B(n_29), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_366), .A2(n_163), .B(n_156), .Y(n_417) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_355), .B(n_163), .C(n_156), .D(n_33), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_381), .Y(n_419) );
NAND4xp25_ASAP7_75t_L g420 ( .A(n_407), .B(n_376), .C(n_380), .D(n_379), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_412), .Y(n_421) );
OAI21xp5_ASAP7_75t_L g422 ( .A1(n_392), .A2(n_379), .B(n_380), .Y(n_422) );
INVxp67_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_407), .B(n_382), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_398), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_390), .A2(n_389), .B(n_384), .Y(n_426) );
INVx6_ASAP7_75t_L g427 ( .A(n_408), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_408), .Y(n_428) );
NAND2x1_ASAP7_75t_SL g429 ( .A(n_414), .B(n_389), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_394), .A2(n_364), .B(n_359), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_391), .B(n_156), .Y(n_431) );
AOI211xp5_ASAP7_75t_L g432 ( .A1(n_418), .A2(n_393), .B(n_399), .C(n_402), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_411), .B(n_30), .C(n_31), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_415), .B(n_34), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_403), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_396), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_419), .A2(n_43), .B1(n_44), .B2(n_47), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_409), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_415), .B(n_52), .Y(n_439) );
NOR2xp33_ASAP7_75t_R g440 ( .A(n_435), .B(n_413), .Y(n_440) );
AOI211x1_ASAP7_75t_SL g441 ( .A1(n_422), .A2(n_416), .B(n_404), .C(n_406), .Y(n_441) );
AOI321xp33_ASAP7_75t_L g442 ( .A1(n_432), .A2(n_416), .A3(n_400), .B1(n_404), .B2(n_417), .C(n_401), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_438), .Y(n_443) );
OAI21xp33_ASAP7_75t_SL g444 ( .A1(n_429), .A2(n_405), .B(n_410), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_425), .Y(n_445) );
XNOR2xp5_ASAP7_75t_L g446 ( .A(n_436), .B(n_420), .Y(n_446) );
OAI21xp33_ASAP7_75t_SL g447 ( .A1(n_430), .A2(n_431), .B(n_428), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_427), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_426), .B(n_424), .Y(n_449) );
OA211x2_ASAP7_75t_L g450 ( .A1(n_437), .A2(n_433), .B(n_434), .C(n_439), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_427), .B(n_437), .Y(n_451) );
NOR2xp33_ASAP7_75t_SL g452 ( .A(n_427), .B(n_435), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_435), .A2(n_395), .B1(n_422), .B2(n_438), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_421), .B(n_392), .Y(n_454) );
OAI211xp5_ASAP7_75t_L g455 ( .A1(n_422), .A2(n_432), .B(n_392), .C(n_423), .Y(n_455) );
OAI21x1_ASAP7_75t_L g456 ( .A1(n_454), .A2(n_446), .B(n_451), .Y(n_456) );
BUFx4f_ASAP7_75t_SL g457 ( .A(n_443), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_445), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_444), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_440), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_460), .A2(n_453), .B1(n_455), .B2(n_449), .Y(n_461) );
NAND4xp25_ASAP7_75t_L g462 ( .A(n_459), .B(n_450), .C(n_441), .D(n_442), .Y(n_462) );
INVx3_ASAP7_75t_SL g463 ( .A(n_457), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_461), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_463), .Y(n_465) );
OR2x6_ASAP7_75t_L g466 ( .A(n_465), .B(n_456), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_464), .Y(n_467) );
AOI322xp5_ASAP7_75t_L g468 ( .A1(n_467), .A2(n_459), .A3(n_447), .B1(n_456), .B2(n_462), .C1(n_448), .C2(n_452), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_468), .A2(n_466), .B(n_458), .Y(n_469) );
endmodule