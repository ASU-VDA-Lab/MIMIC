module real_jpeg_33033_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_261;
wire n_86;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_0),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_0),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_0),
.Y(n_313)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_0),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_1),
.B(n_60),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_1),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_1),
.B(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_1),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_1),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_1),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_1),
.B(n_432),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_1),
.Y(n_455)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_2),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_2),
.B(n_262),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_2),
.B(n_448),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_SL g478 ( 
.A(n_2),
.B(n_479),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx11_ASAP7_75t_R g552 ( 
.A(n_3),
.Y(n_552)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_4),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_4),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_4),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_4),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_4),
.B(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_6),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_6),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_6),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_8),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_9),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_9),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_9),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_9),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_9),
.B(n_128),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_9),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_9),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_10),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_10),
.B(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_10),
.B(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_10),
.Y(n_295)
);

AND2x2_ASAP7_75t_SL g446 ( 
.A(n_10),
.B(n_198),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_10),
.B(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_10),
.B(n_490),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_11),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_11),
.Y(n_143)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_11),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_12),
.Y(n_302)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_13),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_14),
.B(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_14),
.A2(n_124),
.B1(n_297),
.B2(n_299),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_14),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_14),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_14),
.B(n_358),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_14),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_14),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_14),
.B(n_495),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_19),
.B(n_20),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_16),
.Y(n_165)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_16),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

NAND2x1_ASAP7_75t_L g71 ( 
.A(n_17),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_17),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_17),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_17),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_17),
.B(n_167),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_249),
.B(n_532),
.C(n_553),
.Y(n_20)
);

NOR2xp67_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_168),
.Y(n_21)
);

OAI211xp5_ASAP7_75t_L g532 ( 
.A1(n_22),
.A2(n_533),
.B(n_536),
.C(n_551),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_105),
.Y(n_22)
);

NAND2xp33_ASAP7_75t_SL g538 ( 
.A(n_23),
.B(n_105),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_88),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_55),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_25),
.B(n_55),
.C(n_88),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.C(n_49),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_26),
.B(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.C(n_36),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_27),
.A2(n_28),
.B1(n_32),
.B2(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_27),
.B(n_115),
.C(n_119),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_27),
.A2(n_28),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_27),
.A2(n_28),
.B1(n_272),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_28),
.B(n_272),
.C(n_275),
.Y(n_271)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_31),
.Y(n_159)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_31),
.Y(n_198)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_32),
.A2(n_113),
.B1(n_543),
.B2(n_544),
.Y(n_542)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_36),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_36),
.A2(n_63),
.B1(n_70),
.B2(n_71),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_36),
.A2(n_63),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_36),
.A2(n_63),
.B1(n_261),
.B2(n_263),
.Y(n_260)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_38),
.Y(n_238)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_40),
.B(n_49),
.Y(n_91)
);

NOR2xp67_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_47),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_48),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_50),
.B(n_94),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_50),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_53),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_54),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_54),
.Y(n_240)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_54),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_75),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_57),
.B(n_62),
.C(n_75),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_61),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.C(n_70),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_63),
.B(n_258),
.C(n_261),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_64),
.B(n_119),
.C(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_66),
.B(n_140),
.Y(n_192)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_68),
.Y(n_326)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_71),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_70),
.A2(n_71),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_71),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_71),
.Y(n_548)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_74),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_76),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_123),
.C(n_127),
.Y(n_122)
);

XOR2x2_ASAP7_75t_L g144 ( 
.A(n_77),
.B(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_80),
.Y(n_294)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_83),
.B(n_196),
.C(n_199),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_83),
.A2(n_84),
.B1(n_166),
.B2(n_189),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_83),
.B(n_546),
.C(n_547),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_84),
.B(n_226),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_SL g555 ( 
.A(n_84),
.B(n_113),
.C(n_166),
.Y(n_555)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.C(n_103),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_103),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_100),
.Y(n_92)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_97),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_97),
.B(n_154),
.C(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_97),
.B(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_99),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_99),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_130),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_106),
.B(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_122),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_110),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_114),
.B(n_122),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_115),
.B(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_119),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_119),
.B(n_230),
.Y(n_316)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_121),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_121),
.Y(n_430)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_121),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_127),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_127),
.A2(n_146),
.B1(n_215),
.B2(n_342),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_130),
.A2(n_131),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_148),
.C(n_152),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.C(n_144),
.Y(n_132)
);

XOR2x2_ASAP7_75t_L g246 ( 
.A(n_133),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_136),
.A2(n_230),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_136),
.B(n_230),
.Y(n_435)
);

OAI21xp33_ASAP7_75t_L g466 ( 
.A1(n_136),
.A2(n_230),
.B(n_435),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_137),
.A2(n_138),
.B1(n_144),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_143),
.Y(n_365)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_144),
.Y(n_248)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_146),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_152),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_161),
.C(n_166),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_153)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_156),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_179),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_154),
.B(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_154),
.B(n_428),
.Y(n_462)
);

INVx8_ASAP7_75t_L g504 ( 
.A(n_155),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_157),
.B(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_157),
.B(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_157),
.B(n_329),
.C(n_334),
.Y(n_343)
);

OR2x2_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_162),
.B1(n_166),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_165),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_178),
.C(n_181),
.Y(n_177)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_166),
.A2(n_181),
.B1(n_182),
.B2(n_189),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_205),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_169),
.A2(n_534),
.B(n_535),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_202),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_170),
.B(n_202),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_R g170 ( 
.A(n_171),
.B(n_173),
.C(n_175),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_185),
.C(n_190),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_177),
.A2(n_186),
.B1(n_187),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_178),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_179),
.B(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_179),
.B(n_265),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_180),
.Y(n_497)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g243 ( 
.A(n_190),
.B(n_244),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_195),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_191),
.B(n_195),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_193),
.B(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_200),
.Y(n_226)
);

INVxp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_206),
.B(n_208),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_243),
.C(n_246),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_209),
.B(n_400),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_227),
.C(n_241),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_210),
.B(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_224),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g383 ( 
.A(n_211),
.B(n_384),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_213),
.A2(n_214),
.B1(n_224),
.B2(n_225),
.Y(n_384)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.C(n_220),
.Y(n_214)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_215),
.Y(n_342)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_220),
.Y(n_340)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_227),
.B(n_241),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_236),
.C(n_239),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_228),
.B(n_380),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.C(n_233),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_284)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_232),
.Y(n_492)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_235),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_239),
.Y(n_381)
);

XNOR2x1_ASAP7_75t_L g400 ( 
.A(n_243),
.B(n_246),
.Y(n_400)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_412),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_386),
.B(n_408),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_368),
.B(n_385),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_344),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_254),
.B(n_344),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_304),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_255),
.B(n_305),
.C(n_336),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_281),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g372 ( 
.A(n_256),
.B(n_282),
.C(n_285),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_264),
.C(n_270),
.Y(n_256)
);

XOR2x2_ASAP7_75t_L g366 ( 
.A(n_257),
.B(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_261),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_264),
.B(n_271),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g334 ( 
.A(n_269),
.B(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_269),
.B(n_430),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_269),
.B(n_507),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_272),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_274),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_275),
.B(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_278),
.Y(n_444)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_280),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_296),
.B2(n_303),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_288),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_290),
.Y(n_483)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_291),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_292),
.Y(n_510)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_293),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_295),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_296),
.B(n_377),
.C(n_378),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_298),
.Y(n_456)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OA21x2_ASAP7_75t_SL g306 ( 
.A1(n_303),
.A2(n_307),
.B(n_311),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_336),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_314),
.C(n_327),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_327),
.Y(n_346)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx4f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_314),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_317),
.C(n_322),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_315),
.A2(n_316),
.B1(n_423),
.B2(n_424),
.Y(n_422)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_317),
.A2(n_318),
.B1(n_322),
.B2(n_323),
.Y(n_424)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2x2_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_334),
.Y(n_327)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

XOR2x2_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_343),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_339),
.C(n_343),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.C(n_366),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_345),
.B(n_416),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_366),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_353),
.C(n_354),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_350),
.B(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_353),
.A2(n_354),
.B1(n_355),
.B2(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_361),
.C(n_363),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_356),
.A2(n_357),
.B1(n_361),
.B2(n_362),
.Y(n_470)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_363),
.B(n_470),
.Y(n_469)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_369),
.B(n_531),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_371),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_372),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_383),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_382),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_394),
.C(n_395),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_379),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_382),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_406),
.C(n_407),
.Y(n_405)
);

NAND3xp33_ASAP7_75t_SL g412 ( 
.A(n_386),
.B(n_413),
.C(n_530),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_398),
.B1(n_401),
.B2(n_404),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_388),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_399),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_399),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.C(n_396),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_390),
.B(n_396),
.Y(n_403)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_405),
.Y(n_410)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_410),
.B(n_411),
.Y(n_408)
);

AO21x2_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_436),
.B(n_529),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_417),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_415),
.B(n_417),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_422),
.C(n_425),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_418),
.A2(n_419),
.B1(n_527),
.B2(n_528),
.Y(n_526)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_419),
.B(n_523),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_422),
.B(n_425),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_422),
.B(n_425),
.Y(n_528)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_431),
.C(n_434),
.Y(n_425)
);

XNOR2x1_ASAP7_75t_L g464 ( 
.A(n_426),
.B(n_465),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_431),
.A2(n_434),
.B1(n_466),
.B2(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_431),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_437),
.A2(n_521),
.B(n_525),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_472),
.B(n_520),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_463),
.Y(n_438)
);

NOR2x1_ASAP7_75t_L g520 ( 
.A(n_439),
.B(n_463),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_452),
.C(n_462),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_441),
.B(n_517),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_445),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_446),
.C(n_451),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_443),
.B(n_502),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_447),
.B1(n_450),
.B2(n_451),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_446),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_447),
.Y(n_451)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

AO22x1_ASAP7_75t_L g517 ( 
.A1(n_452),
.A2(n_453),
.B1(n_462),
.B2(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_457),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_454),
.A2(n_457),
.B1(n_458),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_462),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_468),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_464),
.B(n_469),
.C(n_471),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_514),
.B(n_519),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_498),
.B(n_513),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_487),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_475),
.B(n_487),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_477),
.B1(n_484),
.B2(n_485),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_478),
.B(n_481),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_478),
.B(n_481),
.C(n_484),
.Y(n_515)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_493),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_488),
.A2(n_489),
.B1(n_493),
.B2(n_494),
.Y(n_511)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx3_ASAP7_75t_SL g490 ( 
.A(n_491),
.Y(n_490)
);

INVx8_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_505),
.B(n_512),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_511),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_511),
.Y(n_512)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_516),
.Y(n_519)
);

NOR2x1p5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_524),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

NOR3xp33_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_539),
.C(n_545),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_550),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_549),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_545),
.Y(n_541)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_548),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_551),
.B(n_554),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_555),
.Y(n_554)
);


endmodule