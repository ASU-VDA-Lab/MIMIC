module fake_jpeg_20761_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_21),
.B1(n_22),
.B2(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx6p67_ASAP7_75t_R g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_7),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_10),
.B1(n_11),
.B2(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_34),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_21),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_27),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_27),
.B(n_12),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_8),
.B(n_15),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_47),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_31),
.C(n_35),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_38),
.Y(n_50)
);

XNOR2x1_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_29),
.B1(n_17),
.B2(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_42),
.Y(n_55)
);

AO21x1_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_54),
.B(n_49),
.Y(n_56)
);

AOI322xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_9),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.C1(n_6),
.C2(n_7),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_5),
.Y(n_58)
);


endmodule