module real_aes_9724_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_2014;
wire n_1314;
wire n_2003;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_2006;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_2021;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1994;
wire n_1225;
wire n_1441;
wire n_1382;
wire n_951;
wire n_875;
wire n_1199;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_2016;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_2022;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_2018;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_1600;
wire n_805;
wire n_619;
wire n_1250;
wire n_1284;
wire n_1095;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_2004;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_2024;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1940;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_2007;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_2012;
wire n_1018;
wire n_1563;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_1712;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_2020;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_2017;
wire n_1946;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_2009;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_2005;
wire n_508;
wire n_1141;
wire n_1985;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_2023;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_2015;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_2019;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_2013;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_2008;
wire n_1722;
wire n_528;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1078;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_2025;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_2011;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1931;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_1596;
wire n_987;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_2010;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_2026;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_729;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
XNOR2xp5_ASAP7_75t_L g870 ( .A(n_0), .B(n_871), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_1), .A2(n_342), .B1(n_1278), .B2(n_1279), .Y(n_1277) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1), .Y(n_1305) );
INVx1_ASAP7_75t_L g1033 ( .A(n_2), .Y(n_1033) );
CKINVDCx5p33_ASAP7_75t_R g1946 ( .A(n_3), .Y(n_1946) );
CKINVDCx5p33_ASAP7_75t_R g1963 ( .A(n_4), .Y(n_1963) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_5), .A2(n_266), .B1(n_527), .B2(n_604), .C(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g635 ( .A(n_5), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g1497 ( .A1(n_6), .A2(n_115), .B1(n_1444), .B2(n_1446), .Y(n_1497) );
INVx1_ASAP7_75t_L g1529 ( .A(n_6), .Y(n_1529) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_7), .A2(n_334), .B1(n_456), .B2(n_460), .Y(n_455) );
INVx1_ASAP7_75t_L g540 ( .A(n_7), .Y(n_540) );
INVxp33_ASAP7_75t_SL g1995 ( .A(n_8), .Y(n_1995) );
AOI22xp5_ASAP7_75t_SL g2019 ( .A1(n_8), .A2(n_318), .B1(n_1186), .B2(n_2020), .Y(n_2019) );
INVx1_ASAP7_75t_L g695 ( .A(n_9), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_9), .A2(n_163), .B1(n_666), .B2(n_752), .Y(n_751) );
CKINVDCx5p33_ASAP7_75t_R g1273 ( .A(n_10), .Y(n_1273) );
INVx1_ASAP7_75t_L g1137 ( .A(n_11), .Y(n_1137) );
INVx1_ASAP7_75t_L g1722 ( .A(n_12), .Y(n_1722) );
AOI22xp33_ASAP7_75t_L g1971 ( .A1(n_12), .A2(n_1972), .B1(n_1977), .B2(n_2023), .Y(n_1971) );
AO22x1_ASAP7_75t_L g1980 ( .A1(n_12), .A2(n_1722), .B1(n_1981), .B2(n_2022), .Y(n_1980) );
INVx1_ASAP7_75t_L g1587 ( .A(n_13), .Y(n_1587) );
AOI22xp33_ASAP7_75t_L g1606 ( .A1(n_13), .A2(n_126), .B1(n_1281), .B2(n_1607), .Y(n_1606) );
INVx1_ASAP7_75t_L g894 ( .A(n_14), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_14), .A2(n_212), .B1(n_905), .B2(n_906), .Y(n_904) );
AOI221xp5_ASAP7_75t_L g1222 ( .A1(n_15), .A2(n_33), .B1(n_656), .B2(n_1223), .C(n_1225), .Y(n_1222) );
INVx1_ASAP7_75t_L g1253 ( .A(n_15), .Y(n_1253) );
AOI22xp33_ASAP7_75t_SL g2004 ( .A1(n_16), .A2(n_256), .B1(n_622), .B2(n_2005), .Y(n_2004) );
AOI22xp33_ASAP7_75t_L g2014 ( .A1(n_16), .A2(n_256), .B1(n_2015), .B2(n_2017), .Y(n_2014) );
OAI22xp33_ASAP7_75t_L g1559 ( .A1(n_17), .A2(n_112), .B1(n_485), .B2(n_516), .Y(n_1559) );
AOI221xp5_ASAP7_75t_L g1565 ( .A1(n_17), .A2(n_112), .B1(n_1193), .B2(n_1395), .C(n_1566), .Y(n_1565) );
AOI221xp5_ASAP7_75t_L g1014 ( .A1(n_18), .A2(n_290), .B1(n_691), .B2(n_709), .C(n_775), .Y(n_1014) );
OAI22xp33_ASAP7_75t_L g1020 ( .A1(n_18), .A2(n_123), .B1(n_927), .B2(n_929), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1595 ( .A1(n_19), .A2(n_133), .B1(n_1403), .B2(n_1596), .Y(n_1595) );
AOI22xp33_ASAP7_75t_SL g1603 ( .A1(n_19), .A2(n_133), .B1(n_1197), .B2(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1173 ( .A(n_20), .Y(n_1173) );
AOI22xp33_ASAP7_75t_SL g1188 ( .A1(n_20), .A2(n_305), .B1(n_1189), .B2(n_1191), .Y(n_1188) );
INVx1_ASAP7_75t_L g425 ( .A(n_21), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g1443 ( .A1(n_22), .A2(n_79), .B1(n_1444), .B2(n_1446), .Y(n_1443) );
OAI22xp33_ASAP7_75t_L g1453 ( .A1(n_22), .A2(n_207), .B1(n_390), .B2(n_1352), .Y(n_1453) );
CKINVDCx16_ASAP7_75t_R g595 ( .A(n_23), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_24), .A2(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g715 ( .A(n_24), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g1698 ( .A1(n_25), .A2(n_144), .B1(n_1680), .B2(n_1688), .Y(n_1698) );
INVx1_ASAP7_75t_L g800 ( .A(n_26), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_26), .A2(n_139), .B1(n_581), .B2(n_658), .Y(n_854) );
AOI22xp33_ASAP7_75t_SL g1597 ( .A1(n_27), .A2(n_104), .B1(n_1403), .B2(n_1598), .Y(n_1597) );
INVxp67_ASAP7_75t_SL g1622 ( .A(n_27), .Y(n_1622) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_28), .A2(n_152), .B1(n_1217), .B2(n_1218), .Y(n_1216) );
INVx1_ASAP7_75t_L g1238 ( .A(n_28), .Y(n_1238) );
INVx1_ASAP7_75t_L g1438 ( .A(n_29), .Y(n_1438) );
OAI222xp33_ASAP7_75t_L g1450 ( .A1(n_29), .A2(n_253), .B1(n_352), .B2(n_706), .C1(n_1451), .C2(n_1452), .Y(n_1450) );
CKINVDCx5p33_ASAP7_75t_R g1219 ( .A(n_30), .Y(n_1219) );
AOI22xp33_ASAP7_75t_SL g1397 ( .A1(n_31), .A2(n_150), .B1(n_1185), .B2(n_1279), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_31), .A2(n_150), .B1(n_600), .B2(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g618 ( .A(n_32), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g667 ( .A1(n_32), .A2(n_325), .B1(n_668), .B2(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g1249 ( .A(n_33), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_34), .A2(n_80), .B1(n_600), .B2(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g638 ( .A(n_34), .Y(n_638) );
INVx1_ASAP7_75t_L g610 ( .A(n_35), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_35), .A2(n_188), .B1(n_660), .B2(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g1381 ( .A(n_36), .Y(n_1381) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_36), .A2(n_355), .B1(n_609), .B2(n_1407), .Y(n_1406) );
NOR2xp33_ASAP7_75t_L g1496 ( .A(n_37), .B(n_1442), .Y(n_1496) );
INVx1_ASAP7_75t_L g1527 ( .A(n_37), .Y(n_1527) );
INVx1_ASAP7_75t_L g1928 ( .A(n_38), .Y(n_1928) );
AOI221xp5_ASAP7_75t_L g1953 ( .A1(n_38), .A2(n_175), .B1(n_1213), .B2(n_1214), .C(n_1954), .Y(n_1953) );
CKINVDCx5p33_ASAP7_75t_R g1151 ( .A(n_39), .Y(n_1151) );
INVx1_ASAP7_75t_L g381 ( .A(n_40), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g1679 ( .A1(n_41), .A2(n_138), .B1(n_1680), .B2(n_1688), .Y(n_1679) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_42), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_43), .A2(n_131), .B1(n_546), .B2(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g652 ( .A(n_43), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g1440 ( .A1(n_44), .A2(n_132), .B1(n_1441), .B2(n_1442), .Y(n_1440) );
AOI22xp33_ASAP7_75t_SL g1461 ( .A1(n_44), .A2(n_132), .B1(n_600), .B2(n_1405), .Y(n_1461) );
AOI21xp33_ASAP7_75t_L g690 ( .A1(n_45), .A2(n_623), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g748 ( .A(n_45), .Y(n_748) );
INVx1_ASAP7_75t_L g1036 ( .A(n_46), .Y(n_1036) );
OAI211xp5_ASAP7_75t_SL g1062 ( .A1(n_46), .A2(n_516), .B(n_1063), .C(n_1068), .Y(n_1062) );
INVx1_ASAP7_75t_L g1794 ( .A(n_47), .Y(n_1794) );
AOI22xp5_ASAP7_75t_L g1921 ( .A1(n_48), .A2(n_1922), .B1(n_1964), .B2(n_1965), .Y(n_1921) );
CKINVDCx5p33_ASAP7_75t_R g1964 ( .A(n_48), .Y(n_1964) );
INVx1_ASAP7_75t_L g1991 ( .A(n_49), .Y(n_1991) );
XOR2xp5_ASAP7_75t_L g405 ( .A(n_50), .B(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_SL g1588 ( .A(n_51), .Y(n_1588) );
OAI22xp33_ASAP7_75t_L g1613 ( .A1(n_51), .A2(n_197), .B1(n_1385), .B2(n_1614), .Y(n_1613) );
INVx1_ASAP7_75t_L g1629 ( .A(n_52), .Y(n_1629) );
AOI22xp33_ASAP7_75t_L g1658 ( .A1(n_52), .A2(n_232), .B1(n_1329), .B2(n_1407), .Y(n_1658) );
INVxp33_ASAP7_75t_SL g2001 ( .A(n_53), .Y(n_2001) );
AOI22xp33_ASAP7_75t_L g2021 ( .A1(n_53), .A2(n_316), .B1(n_731), .B2(n_2015), .Y(n_2021) );
INVx1_ASAP7_75t_L g1320 ( .A(n_54), .Y(n_1320) );
AOI22xp33_ASAP7_75t_L g1361 ( .A1(n_54), .A2(n_308), .B1(n_815), .B2(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1455 ( .A(n_55), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1469 ( .A1(n_55), .A2(n_249), .B1(n_750), .B2(n_1375), .Y(n_1469) );
AOI22xp33_ASAP7_75t_L g1655 ( .A1(n_56), .A2(n_167), .B1(n_1298), .B2(n_1329), .Y(n_1655) );
AOI22xp33_ASAP7_75t_L g1661 ( .A1(n_56), .A2(n_167), .B1(n_1189), .B2(n_1395), .Y(n_1661) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_57), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_58), .A2(n_269), .B1(n_1281), .B2(n_1282), .Y(n_1280) );
INVx1_ASAP7_75t_L g1302 ( .A(n_58), .Y(n_1302) );
INVx1_ASAP7_75t_L g1935 ( .A(n_59), .Y(n_1935) );
AOI22xp33_ASAP7_75t_L g1961 ( .A1(n_59), .A2(n_149), .B1(n_581), .B2(n_993), .Y(n_1961) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_60), .Y(n_816) );
AOI22x1_ASAP7_75t_SL g1430 ( .A1(n_61), .A2(n_1431), .B1(n_1470), .B2(n_1471), .Y(n_1430) );
INVx1_ASAP7_75t_L g1470 ( .A(n_61), .Y(n_1470) );
INVx1_ASAP7_75t_L g1106 ( .A(n_62), .Y(n_1106) );
INVx1_ASAP7_75t_L g1205 ( .A(n_63), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1699 ( .A1(n_63), .A2(n_82), .B1(n_1692), .B2(n_1696), .Y(n_1699) );
INVx1_ASAP7_75t_L g989 ( .A(n_64), .Y(n_989) );
OAI221xp5_ASAP7_75t_L g1000 ( .A1(n_64), .A2(n_485), .B1(n_512), .B2(n_1001), .C(n_1007), .Y(n_1000) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_65), .A2(n_267), .B1(n_456), .B2(n_460), .Y(n_1043) );
INVx1_ASAP7_75t_L g1066 ( .A(n_65), .Y(n_1066) );
INVx1_ASAP7_75t_L g509 ( .A(n_66), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_66), .A2(n_251), .B1(n_568), .B2(n_571), .Y(n_567) );
INVx1_ASAP7_75t_L g951 ( .A(n_67), .Y(n_951) );
INVx1_ASAP7_75t_L g1390 ( .A(n_68), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_68), .A2(n_204), .B1(n_1403), .B2(n_1405), .Y(n_1402) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_69), .A2(n_257), .B1(n_626), .B2(n_627), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_69), .A2(n_257), .B1(n_656), .B2(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g1347 ( .A(n_70), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g1374 ( .A1(n_70), .A2(n_299), .B1(n_750), .B2(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1350 ( .A(n_71), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1373 ( .A1(n_71), .A2(n_332), .B1(n_581), .B2(n_663), .Y(n_1373) );
INVx1_ASAP7_75t_L g496 ( .A(n_72), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_72), .A2(n_213), .B1(n_574), .B2(n_577), .Y(n_573) );
INVx1_ASAP7_75t_L g1543 ( .A(n_73), .Y(n_1543) );
AOI221xp5_ASAP7_75t_L g1561 ( .A1(n_73), .A2(n_278), .B1(n_1395), .B2(n_1562), .C(n_1564), .Y(n_1561) );
AOI22xp33_ASAP7_75t_L g1732 ( .A1(n_74), .A2(n_222), .B1(n_1680), .B2(n_1688), .Y(n_1732) );
OAI22xp33_ASAP7_75t_L g1147 ( .A1(n_75), .A2(n_339), .B1(n_549), .B2(n_554), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_75), .A2(n_339), .B1(n_1196), .B2(n_1197), .Y(n_1195) );
AO22x1_ASAP7_75t_SL g1701 ( .A1(n_76), .A2(n_147), .B1(n_1680), .B2(n_1688), .Y(n_1701) );
INVx1_ASAP7_75t_L g1326 ( .A(n_77), .Y(n_1326) );
OAI22xp5_ASAP7_75t_L g1336 ( .A1(n_77), .A2(n_353), .B1(n_1337), .B2(n_1339), .Y(n_1336) );
AOI22xp33_ASAP7_75t_L g1653 ( .A1(n_78), .A2(n_214), .B1(n_1403), .B2(n_1654), .Y(n_1653) );
AOI22xp33_ASAP7_75t_L g1660 ( .A1(n_78), .A2(n_214), .B1(n_658), .B2(n_1604), .Y(n_1660) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_79), .A2(n_162), .B1(n_1329), .B2(n_1359), .Y(n_1462) );
INVx1_ASAP7_75t_L g636 ( .A(n_80), .Y(n_636) );
INVxp33_ASAP7_75t_SL g1083 ( .A(n_81), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_81), .A2(n_368), .B1(n_1122), .B2(n_1124), .Y(n_1121) );
INVx1_ASAP7_75t_L g466 ( .A(n_83), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g1230 ( .A(n_84), .Y(n_1230) );
CKINVDCx5p33_ASAP7_75t_R g1266 ( .A(n_85), .Y(n_1266) );
AOI22xp33_ASAP7_75t_SL g1459 ( .A1(n_86), .A2(n_170), .B1(n_691), .B2(n_1329), .Y(n_1459) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_86), .A2(n_170), .B1(n_581), .B2(n_582), .Y(n_1466) );
AOI22xp5_ASAP7_75t_L g1733 ( .A1(n_87), .A2(n_246), .B1(n_1696), .B2(n_1712), .Y(n_1733) );
CKINVDCx5p33_ASAP7_75t_R g941 ( .A(n_88), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_89), .A2(n_272), .B1(n_838), .B2(n_1127), .Y(n_1220) );
OAI221xp5_ASAP7_75t_L g1244 ( .A1(n_89), .A2(n_272), .B1(n_783), .B2(n_788), .C(n_1087), .Y(n_1244) );
INVx1_ASAP7_75t_L g1039 ( .A(n_90), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_90), .A2(n_248), .B1(n_905), .B2(n_906), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1283 ( .A1(n_91), .A2(n_370), .B1(n_1193), .B2(n_1282), .Y(n_1283) );
OAI221xp5_ASAP7_75t_L g1300 ( .A1(n_91), .A2(n_485), .B1(n_1061), .B2(n_1301), .C(n_1304), .Y(n_1300) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_92), .Y(n_829) );
INVx1_ASAP7_75t_L g1630 ( .A(n_93), .Y(n_1630) );
AOI22xp33_ASAP7_75t_L g1657 ( .A1(n_93), .A2(n_191), .B1(n_1005), .B2(n_1403), .Y(n_1657) );
INVx1_ASAP7_75t_L g1927 ( .A(n_94), .Y(n_1927) );
AOI22xp33_ASAP7_75t_L g1955 ( .A1(n_94), .A2(n_241), .B1(n_668), .B2(n_1956), .Y(n_1955) );
INVx1_ASAP7_75t_L g1990 ( .A(n_95), .Y(n_1990) );
AOI22xp33_ASAP7_75t_SL g2008 ( .A1(n_95), .A2(n_142), .B1(n_607), .B2(n_2005), .Y(n_2008) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_96), .Y(n_887) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_97), .Y(n_1097) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_97), .A2(n_371), .B1(n_574), .B2(n_1132), .C(n_1133), .Y(n_1131) );
INVx1_ASAP7_75t_L g1987 ( .A(n_98), .Y(n_1987) );
INVx1_ASAP7_75t_L g944 ( .A(n_99), .Y(n_944) );
OAI221xp5_ASAP7_75t_L g954 ( .A1(n_99), .A2(n_485), .B1(n_512), .B2(n_955), .C(n_958), .Y(n_954) );
XNOR2x2_ASAP7_75t_L g1534 ( .A(n_100), .B(n_1535), .Y(n_1534) );
AOI22xp5_ASAP7_75t_L g1711 ( .A1(n_100), .A2(n_130), .B1(n_1696), .B2(n_1712), .Y(n_1711) );
INVxp67_ASAP7_75t_SL g1582 ( .A(n_101), .Y(n_1582) );
AOI22xp33_ASAP7_75t_L g1609 ( .A1(n_101), .A2(n_282), .B1(n_993), .B2(n_1604), .Y(n_1609) );
OAI221xp5_ASAP7_75t_L g1932 ( .A1(n_102), .A2(n_137), .B1(n_783), .B2(n_788), .C(n_1087), .Y(n_1932) );
OAI22xp5_ASAP7_75t_L g1958 ( .A1(n_102), .A2(n_137), .B1(n_838), .B2(n_1127), .Y(n_1958) );
CKINVDCx5p33_ASAP7_75t_R g1552 ( .A(n_103), .Y(n_1552) );
INVxp33_ASAP7_75t_L g1621 ( .A(n_104), .Y(n_1621) );
INVx1_ASAP7_75t_L g424 ( .A(n_105), .Y(n_424) );
BUFx2_ASAP7_75t_L g469 ( .A(n_105), .Y(n_469) );
BUFx2_ASAP7_75t_L g474 ( .A(n_105), .Y(n_474) );
OR2x2_ASAP7_75t_L g787 ( .A(n_105), .B(n_479), .Y(n_787) );
AOI22xp33_ASAP7_75t_SL g1460 ( .A1(n_106), .A2(n_263), .B1(n_626), .B2(n_1405), .Y(n_1460) );
AOI22xp33_ASAP7_75t_L g1464 ( .A1(n_106), .A2(n_263), .B1(n_669), .B2(n_1465), .Y(n_1464) );
INVx1_ASAP7_75t_L g683 ( .A(n_107), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_107), .A2(n_153), .B1(n_669), .B2(n_758), .Y(n_757) );
OAI22xp33_ASAP7_75t_L g949 ( .A1(n_108), .A2(n_120), .B1(n_410), .B2(n_427), .Y(n_949) );
INVx1_ASAP7_75t_L g971 ( .A(n_108), .Y(n_971) );
INVx1_ASAP7_75t_L g1796 ( .A(n_109), .Y(n_1796) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_110), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g1394 ( .A1(n_111), .A2(n_365), .B1(n_1189), .B2(n_1395), .Y(n_1394) );
AOI22xp33_ASAP7_75t_SL g1411 ( .A1(n_111), .A2(n_365), .B1(n_1407), .B2(n_1412), .Y(n_1411) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_113), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_114), .A2(n_375), .B1(n_626), .B2(n_627), .Y(n_1360) );
AOI22xp33_ASAP7_75t_SL g1369 ( .A1(n_114), .A2(n_375), .B1(n_1370), .B2(n_1371), .Y(n_1369) );
INVx1_ASAP7_75t_L g1489 ( .A(n_115), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_116), .A2(n_177), .B1(n_1325), .B2(n_1385), .Y(n_1384) );
OAI22xp33_ASAP7_75t_L g1421 ( .A1(n_116), .A2(n_177), .B1(n_1339), .B2(n_1422), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1728 ( .A1(n_117), .A2(n_327), .B1(n_1680), .B2(n_1688), .Y(n_1728) );
CKINVDCx5p33_ASAP7_75t_R g1541 ( .A(n_118), .Y(n_1541) );
INVx1_ASAP7_75t_L g1269 ( .A(n_119), .Y(n_1269) );
AOI221xp5_ASAP7_75t_L g1295 ( .A1(n_119), .A2(n_315), .B1(n_527), .B2(n_1296), .C(n_1298), .Y(n_1295) );
INVx1_ASAP7_75t_L g970 ( .A(n_120), .Y(n_970) );
OAI221xp5_ASAP7_75t_L g1085 ( .A1(n_121), .A2(n_206), .B1(n_783), .B2(n_1086), .C(n_1087), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_121), .A2(n_206), .B1(n_1127), .B2(n_1129), .Y(n_1126) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_122), .A2(n_208), .B1(n_621), .B2(n_622), .C(n_623), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_122), .A2(n_208), .B1(n_660), .B2(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g1012 ( .A(n_123), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1599 ( .A1(n_124), .A2(n_220), .B1(n_1407), .B2(n_1600), .Y(n_1599) );
INVxp67_ASAP7_75t_SL g1612 ( .A(n_124), .Y(n_1612) );
INVx1_ASAP7_75t_L g1322 ( .A(n_125), .Y(n_1322) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_125), .A2(n_145), .B1(n_622), .B2(n_1365), .Y(n_1364) );
INVxp33_ASAP7_75t_L g1584 ( .A(n_126), .Y(n_1584) );
AOI22xp33_ASAP7_75t_L g1691 ( .A1(n_127), .A2(n_293), .B1(n_1692), .B2(n_1696), .Y(n_1691) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_128), .A2(n_485), .B1(n_490), .B2(n_502), .C(n_512), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_128), .A2(n_287), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_129), .A2(n_294), .B1(n_581), .B2(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1254 ( .A(n_129), .Y(n_1254) );
INVx1_ASAP7_75t_L g651 ( .A(n_131), .Y(n_651) );
XNOR2x2_ASAP7_75t_L g1312 ( .A(n_134), .B(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1992 ( .A(n_135), .Y(n_1992) );
INVx1_ASAP7_75t_L g948 ( .A(n_136), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_136), .A2(n_244), .B1(n_905), .B2(n_906), .Y(n_953) );
INVx1_ASAP7_75t_L g809 ( .A(n_139), .Y(n_809) );
INVx1_ASAP7_75t_L g1035 ( .A(n_140), .Y(n_1035) );
OAI221xp5_ASAP7_75t_L g1049 ( .A1(n_140), .A2(n_485), .B1(n_1050), .B2(n_1055), .C(n_1061), .Y(n_1049) );
XNOR2xp5_ASAP7_75t_L g931 ( .A(n_141), .B(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g1704 ( .A(n_141), .Y(n_1704) );
INVxp33_ASAP7_75t_SL g1984 ( .A(n_142), .Y(n_1984) );
CKINVDCx5p33_ASAP7_75t_R g986 ( .A(n_143), .Y(n_986) );
INVx1_ASAP7_75t_L g1316 ( .A(n_145), .Y(n_1316) );
OA22x2_ASAP7_75t_L g1476 ( .A1(n_146), .A2(n_1477), .B1(n_1532), .B2(n_1533), .Y(n_1476) );
INVxp67_ASAP7_75t_SL g1533 ( .A(n_146), .Y(n_1533) );
XNOR2xp5_ASAP7_75t_L g1260 ( .A(n_148), .B(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1941 ( .A(n_149), .Y(n_1941) );
CKINVDCx5p33_ASAP7_75t_R g1159 ( .A(n_151), .Y(n_1159) );
INVx1_ASAP7_75t_L g1243 ( .A(n_152), .Y(n_1243) );
INVx1_ASAP7_75t_L g684 ( .A(n_153), .Y(n_684) );
INVx1_ASAP7_75t_L g454 ( .A(n_154), .Y(n_454) );
INVx1_ASAP7_75t_L g1645 ( .A(n_155), .Y(n_1645) );
AOI22xp33_ASAP7_75t_SL g1663 ( .A1(n_155), .A2(n_335), .B1(n_1395), .B2(n_1664), .Y(n_1663) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_156), .A2(n_180), .B1(n_1285), .B2(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1424 ( .A(n_156), .Y(n_1424) );
CKINVDCx5p33_ASAP7_75t_R g1547 ( .A(n_157), .Y(n_1547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_158), .A2(n_309), .B1(n_549), .B2(n_554), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_158), .A2(n_309), .B1(n_584), .B2(n_587), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_159), .A2(n_216), .B1(n_1185), .B2(n_1285), .Y(n_1284) );
OAI22xp5_ASAP7_75t_L g1309 ( .A1(n_159), .A2(n_216), .B1(n_549), .B2(n_554), .Y(n_1309) );
INVx1_ASAP7_75t_L g1169 ( .A(n_160), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_160), .A2(n_310), .B1(n_1185), .B2(n_1186), .Y(n_1184) );
CKINVDCx5p33_ASAP7_75t_R g1270 ( .A(n_161), .Y(n_1270) );
INVx1_ASAP7_75t_L g1435 ( .A(n_162), .Y(n_1435) );
INVx1_ASAP7_75t_L g688 ( .A(n_163), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g1490 ( .A(n_164), .Y(n_1490) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_165), .Y(n_705) );
XOR2xp5_ASAP7_75t_L g1073 ( .A(n_166), .B(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1684 ( .A(n_168), .Y(n_1684) );
OAI22xp33_ASAP7_75t_L g994 ( .A1(n_169), .A2(n_356), .B1(n_995), .B2(n_997), .Y(n_994) );
INVx1_ASAP7_75t_L g1016 ( .A(n_169), .Y(n_1016) );
INVx1_ASAP7_75t_L g1640 ( .A(n_171), .Y(n_1640) );
AOI22xp33_ASAP7_75t_L g1665 ( .A1(n_171), .A2(n_211), .B1(n_442), .B2(n_658), .Y(n_1665) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_172), .A2(n_374), .B1(n_657), .B2(n_896), .Y(n_987) );
INVx1_ASAP7_75t_L g1003 ( .A(n_172), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g1790 ( .A1(n_173), .A2(n_268), .B1(n_1791), .B2(n_1792), .C(n_1793), .Y(n_1790) );
INVx1_ASAP7_75t_L g1178 ( .A(n_174), .Y(n_1178) );
INVx1_ASAP7_75t_L g1930 ( .A(n_175), .Y(n_1930) );
INVx1_ASAP7_75t_L g1585 ( .A(n_176), .Y(n_1585) );
INVx1_ASAP7_75t_L g803 ( .A(n_178), .Y(n_803) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_178), .A2(n_224), .B1(n_576), .B2(n_849), .C(n_852), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g2006 ( .A1(n_179), .A2(n_321), .B1(n_537), .B2(n_1362), .Y(n_2006) );
AOI22xp33_ASAP7_75t_L g2010 ( .A1(n_179), .A2(n_321), .B1(n_2011), .B2(n_2012), .Y(n_2010) );
INVx1_ASAP7_75t_L g1426 ( .A(n_180), .Y(n_1426) );
INVx1_ASAP7_75t_L g1030 ( .A(n_181), .Y(n_1030) );
INVx1_ASAP7_75t_L g1685 ( .A(n_182), .Y(n_1685) );
NAND2xp5_ASAP7_75t_L g1690 ( .A(n_182), .B(n_1683), .Y(n_1690) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_183), .A2(n_326), .B1(n_600), .B2(n_703), .C(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g728 ( .A(n_183), .Y(n_728) );
INVx1_ASAP7_75t_L g991 ( .A(n_184), .Y(n_991) );
OAI211xp5_ASAP7_75t_SL g1009 ( .A1(n_184), .A2(n_516), .B(n_1010), .C(n_1015), .Y(n_1009) );
INVxp33_ASAP7_75t_SL g1985 ( .A(n_185), .Y(n_1985) );
AOI22xp33_ASAP7_75t_L g2007 ( .A1(n_185), .A2(n_275), .B1(n_1362), .B2(n_1943), .Y(n_2007) );
INVx1_ASAP7_75t_L g777 ( .A(n_186), .Y(n_777) );
AOI21xp33_ASAP7_75t_L g844 ( .A1(n_186), .A2(n_845), .B(n_846), .Y(n_844) );
INVx2_ASAP7_75t_L g393 ( .A(n_187), .Y(n_393) );
INVx1_ASAP7_75t_L g629 ( .A(n_188), .Y(n_629) );
INVx1_ASAP7_75t_L g779 ( .A(n_189), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_189), .A2(n_243), .B1(n_579), .B2(n_657), .Y(n_843) );
AO221x2_ASAP7_75t_L g1716 ( .A1(n_190), .A2(n_231), .B1(n_1692), .B2(n_1717), .C(n_1718), .Y(n_1716) );
INVx1_ASAP7_75t_L g1633 ( .A(n_191), .Y(n_1633) );
CKINVDCx5p33_ASAP7_75t_R g1510 ( .A(n_192), .Y(n_1510) );
BUFx3_ASAP7_75t_L g432 ( .A(n_193), .Y(n_432) );
INVx1_ASAP7_75t_L g459 ( .A(n_193), .Y(n_459) );
INVx1_ASAP7_75t_L g1013 ( .A(n_194), .Y(n_1013) );
OAI22xp33_ASAP7_75t_L g1019 ( .A1(n_194), .A2(n_290), .B1(n_460), .B2(n_925), .Y(n_1019) );
CKINVDCx5p33_ASAP7_75t_R g1503 ( .A(n_195), .Y(n_1503) );
OAI22xp33_ASAP7_75t_L g900 ( .A1(n_196), .A2(n_351), .B1(n_410), .B2(n_427), .Y(n_900) );
INVx1_ASAP7_75t_L g920 ( .A(n_196), .Y(n_920) );
INVx1_ASAP7_75t_L g1590 ( .A(n_197), .Y(n_1590) );
CKINVDCx5p33_ASAP7_75t_R g1494 ( .A(n_198), .Y(n_1494) );
INVxp33_ASAP7_75t_SL g1080 ( .A(n_199), .Y(n_1080) );
AOI221xp5_ASAP7_75t_L g1117 ( .A1(n_199), .A2(n_320), .B1(n_581), .B2(n_849), .C(n_1118), .Y(n_1117) );
AOI221xp5_ASAP7_75t_L g918 ( .A1(n_200), .A2(n_364), .B1(n_708), .B2(n_709), .C(n_775), .Y(n_918) );
OAI22xp33_ASAP7_75t_L g926 ( .A1(n_200), .A2(n_217), .B1(n_927), .B2(n_929), .Y(n_926) );
INVx1_ASAP7_75t_L g965 ( .A(n_201), .Y(n_965) );
OAI22xp33_ASAP7_75t_L g974 ( .A1(n_201), .A2(n_203), .B1(n_927), .B2(n_929), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g1558 ( .A1(n_202), .A2(n_345), .B1(n_905), .B2(n_906), .Y(n_1558) );
INVx1_ASAP7_75t_L g1568 ( .A(n_202), .Y(n_1568) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_203), .A2(n_234), .B1(n_609), .B2(n_708), .C(n_709), .Y(n_968) );
INVx1_ASAP7_75t_L g1391 ( .A(n_204), .Y(n_1391) );
OAI221xp5_ASAP7_75t_L g1634 ( .A1(n_205), .A2(n_277), .B1(n_1385), .B2(n_1635), .C(n_1636), .Y(n_1634) );
INVx1_ASAP7_75t_L g1643 ( .A(n_205), .Y(n_1643) );
AOI22xp33_ASAP7_75t_L g1467 ( .A1(n_207), .A2(n_253), .B1(n_1135), .B2(n_1468), .Y(n_1467) );
CKINVDCx5p33_ASAP7_75t_R g1948 ( .A(n_209), .Y(n_1948) );
AOI221xp5_ASAP7_75t_L g1211 ( .A1(n_210), .A2(n_218), .B1(n_1212), .B2(n_1213), .C(n_1214), .Y(n_1211) );
INVx1_ASAP7_75t_L g1242 ( .A(n_210), .Y(n_1242) );
INVx1_ASAP7_75t_L g1641 ( .A(n_211), .Y(n_1641) );
INVx1_ASAP7_75t_L g897 ( .A(n_212), .Y(n_897) );
INVx1_ASAP7_75t_L g501 ( .A(n_213), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g1154 ( .A(n_215), .Y(n_1154) );
INVx1_ASAP7_75t_L g915 ( .A(n_217), .Y(n_915) );
INVx1_ASAP7_75t_L g1240 ( .A(n_218), .Y(n_1240) );
INVx1_ASAP7_75t_L g420 ( .A(n_219), .Y(n_420) );
INVx1_ASAP7_75t_L g566 ( .A(n_219), .Y(n_566) );
INVxp33_ASAP7_75t_L g1618 ( .A(n_220), .Y(n_1618) );
OAI22xp33_ASAP7_75t_L g1044 ( .A1(n_221), .A2(n_297), .B1(n_927), .B2(n_929), .Y(n_1044) );
AOI221xp5_ASAP7_75t_L g1067 ( .A1(n_221), .A2(n_267), .B1(n_606), .B2(n_709), .C(n_775), .Y(n_1067) );
CKINVDCx5p33_ASAP7_75t_R g1514 ( .A(n_223), .Y(n_1514) );
INVx1_ASAP7_75t_L g805 ( .A(n_224), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g1945 ( .A(n_225), .Y(n_1945) );
INVx1_ASAP7_75t_L g1108 ( .A(n_226), .Y(n_1108) );
CKINVDCx5p33_ASAP7_75t_R g1161 ( .A(n_227), .Y(n_1161) );
XOR2x2_ASAP7_75t_L g1144 ( .A(n_228), .B(n_1145), .Y(n_1144) );
CKINVDCx5p33_ASAP7_75t_R g1949 ( .A(n_229), .Y(n_1949) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_230), .Y(n_1388) );
INVx1_ASAP7_75t_L g1637 ( .A(n_232), .Y(n_1637) );
INVxp67_ASAP7_75t_SL g1098 ( .A(n_233), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_233), .A2(n_322), .B1(n_750), .B2(n_1135), .Y(n_1134) );
OAI22xp33_ASAP7_75t_L g973 ( .A1(n_234), .A2(n_341), .B1(n_460), .B2(n_925), .Y(n_973) );
INVx1_ASAP7_75t_L g1937 ( .A(n_235), .Y(n_1937) );
AOI221xp5_ASAP7_75t_L g1960 ( .A1(n_235), .A2(n_254), .B1(n_1212), .B2(n_1225), .C(n_1370), .Y(n_1960) );
AOI22xp5_ASAP7_75t_L g1710 ( .A1(n_236), .A2(n_302), .B1(n_1680), .B2(n_1688), .Y(n_1710) );
CKINVDCx5p33_ASAP7_75t_R g680 ( .A(n_237), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g1556 ( .A(n_238), .Y(n_1556) );
OAI221xp5_ASAP7_75t_L g1569 ( .A1(n_238), .A2(n_410), .B1(n_427), .B2(n_647), .C(n_1570), .Y(n_1569) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_239), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g1729 ( .A1(n_240), .A2(n_328), .B1(n_1696), .B2(n_1712), .Y(n_1729) );
INVx1_ASAP7_75t_L g1931 ( .A(n_241), .Y(n_1931) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_242), .Y(n_678) );
INVx1_ASAP7_75t_L g769 ( .A(n_243), .Y(n_769) );
INVx1_ASAP7_75t_L g947 ( .A(n_244), .Y(n_947) );
INVx1_ASAP7_75t_L g449 ( .A(n_245), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g1032 ( .A(n_247), .Y(n_1032) );
INVx1_ASAP7_75t_L g1038 ( .A(n_248), .Y(n_1038) );
INVx1_ASAP7_75t_L g1456 ( .A(n_249), .Y(n_1456) );
CKINVDCx5p33_ASAP7_75t_R g1158 ( .A(n_250), .Y(n_1158) );
INVx1_ASAP7_75t_L g507 ( .A(n_251), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g878 ( .A(n_252), .Y(n_878) );
INVx1_ASAP7_75t_L g1940 ( .A(n_254), .Y(n_1940) );
CKINVDCx5p33_ASAP7_75t_R g1632 ( .A(n_255), .Y(n_1632) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_258), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_259), .A2(n_340), .B1(n_607), .B2(n_1359), .Y(n_1358) );
AOI22xp33_ASAP7_75t_SL g1372 ( .A1(n_259), .A2(n_340), .B1(n_568), .B2(n_663), .Y(n_1372) );
INVx1_ASAP7_75t_L g1706 ( .A(n_260), .Y(n_1706) );
CKINVDCx16_ASAP7_75t_R g1576 ( .A(n_261), .Y(n_1576) );
INVx1_ASAP7_75t_L g889 ( .A(n_262), .Y(n_889) );
OAI221xp5_ASAP7_75t_L g907 ( .A1(n_262), .A2(n_485), .B1(n_512), .B2(n_908), .C(n_909), .Y(n_907) );
INVx1_ASAP7_75t_L g979 ( .A(n_264), .Y(n_979) );
CKINVDCx20_ASAP7_75t_R g1719 ( .A(n_265), .Y(n_1719) );
INVx1_ASAP7_75t_L g640 ( .A(n_266), .Y(n_640) );
INVx1_ASAP7_75t_L g1303 ( .A(n_269), .Y(n_1303) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_270), .Y(n_884) );
INVx1_ASAP7_75t_L g1028 ( .A(n_271), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g1549 ( .A(n_273), .Y(n_1549) );
OAI22xp5_ASAP7_75t_L g1481 ( .A1(n_274), .A2(n_295), .B1(n_1482), .B2(n_1484), .Y(n_1481) );
INVx1_ASAP7_75t_L g1521 ( .A(n_274), .Y(n_1521) );
INVxp33_ASAP7_75t_SL g1988 ( .A(n_275), .Y(n_1988) );
INVx1_ASAP7_75t_L g984 ( .A(n_276), .Y(n_984) );
AOI21xp33_ASAP7_75t_L g1008 ( .A1(n_276), .A2(n_606), .B(n_623), .Y(n_1008) );
INVx1_ASAP7_75t_L g1644 ( .A(n_277), .Y(n_1644) );
AOI21xp33_ASAP7_75t_L g1544 ( .A1(n_278), .A2(n_480), .B(n_623), .Y(n_1544) );
OAI221xp5_ASAP7_75t_L g1148 ( .A1(n_279), .A2(n_516), .B1(n_1149), .B2(n_1155), .C(n_1160), .Y(n_1148) );
AOI22xp33_ASAP7_75t_SL g1192 ( .A1(n_279), .A2(n_350), .B1(n_1191), .B2(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1234 ( .A(n_280), .Y(n_1234) );
OAI211xp5_ASAP7_75t_L g1485 ( .A1(n_281), .A2(n_801), .B(n_1486), .C(n_1487), .Y(n_1485) );
INVx1_ASAP7_75t_L g1518 ( .A(n_281), .Y(n_1518) );
INVx1_ASAP7_75t_L g1581 ( .A(n_282), .Y(n_1581) );
CKINVDCx5p33_ASAP7_75t_R g1232 ( .A(n_283), .Y(n_1232) );
XNOR2xp5_ASAP7_75t_L g976 ( .A(n_284), .B(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_SL g992 ( .A1(n_285), .A2(n_314), .B1(n_877), .B2(n_993), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_285), .A2(n_314), .B1(n_549), .B2(n_554), .Y(n_999) );
BUFx3_ASAP7_75t_L g415 ( .A(n_286), .Y(n_415) );
INVx1_ASAP7_75t_L g445 ( .A(n_286), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_287), .A2(n_516), .B1(n_523), .B2(n_532), .C(n_541), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_288), .Y(n_681) );
INVx1_ASAP7_75t_L g1046 ( .A(n_289), .Y(n_1046) );
INVx1_ASAP7_75t_L g891 ( .A(n_291), .Y(n_891) );
OAI211xp5_ASAP7_75t_L g912 ( .A1(n_291), .A2(n_516), .B(n_913), .C(n_919), .Y(n_912) );
AO22x2_ASAP7_75t_L g1625 ( .A1(n_292), .A2(n_1626), .B1(n_1666), .B2(n_1667), .Y(n_1625) );
INVxp67_ASAP7_75t_L g1666 ( .A(n_292), .Y(n_1666) );
XNOR2xp5_ASAP7_75t_L g1022 ( .A(n_293), .B(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1247 ( .A(n_294), .Y(n_1247) );
INVx1_ASAP7_75t_L g1520 ( .A(n_295), .Y(n_1520) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_296), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_296), .B(n_358), .Y(n_479) );
AND2x2_ASAP7_75t_L g487 ( .A(n_296), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g531 ( .A(n_296), .Y(n_531) );
INVx1_ASAP7_75t_L g1065 ( .A(n_297), .Y(n_1065) );
AOI21xp33_ASAP7_75t_L g1550 ( .A1(n_298), .A2(n_708), .B(n_709), .Y(n_1550) );
INVx1_ASAP7_75t_L g1572 ( .A(n_298), .Y(n_1572) );
INVx1_ASAP7_75t_L g1344 ( .A(n_299), .Y(n_1344) );
XNOR2xp5_ASAP7_75t_L g1377 ( .A(n_300), .B(n_1378), .Y(n_1377) );
INVx2_ASAP7_75t_L g422 ( .A(n_301), .Y(n_422) );
OR2x2_ASAP7_75t_L g448 ( .A(n_301), .B(n_420), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g1233 ( .A(n_303), .Y(n_1233) );
INVx1_ASAP7_75t_L g917 ( .A(n_304), .Y(n_917) );
OAI22xp33_ASAP7_75t_L g924 ( .A1(n_304), .A2(n_364), .B1(n_460), .B2(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g1176 ( .A(n_305), .Y(n_1176) );
CKINVDCx5p33_ASAP7_75t_R g1539 ( .A(n_306), .Y(n_1539) );
CKINVDCx5p33_ASAP7_75t_R g1508 ( .A(n_307), .Y(n_1508) );
INVx1_ASAP7_75t_L g1317 ( .A(n_308), .Y(n_1317) );
INVx1_ASAP7_75t_L g1166 ( .A(n_310), .Y(n_1166) );
INVx1_ASAP7_75t_L g902 ( .A(n_311), .Y(n_902) );
INVx1_ASAP7_75t_L g945 ( .A(n_312), .Y(n_945) );
OAI211xp5_ASAP7_75t_L g963 ( .A1(n_312), .A2(n_516), .B(n_964), .C(n_969), .Y(n_963) );
INVx1_ASAP7_75t_L g1103 ( .A(n_313), .Y(n_1103) );
INVx1_ASAP7_75t_L g1267 ( .A(n_315), .Y(n_1267) );
INVx1_ASAP7_75t_L g1998 ( .A(n_316), .Y(n_1998) );
CKINVDCx5p33_ASAP7_75t_R g1546 ( .A(n_317), .Y(n_1546) );
INVxp33_ASAP7_75t_SL g1996 ( .A(n_318), .Y(n_1996) );
INVx1_ASAP7_75t_L g764 ( .A(n_319), .Y(n_764) );
INVxp33_ASAP7_75t_L g1082 ( .A(n_320), .Y(n_1082) );
INVxp33_ASAP7_75t_L g1090 ( .A(n_322), .Y(n_1090) );
CKINVDCx5p33_ASAP7_75t_R g1515 ( .A(n_323), .Y(n_1515) );
AOI22xp33_ASAP7_75t_L g1414 ( .A1(n_324), .A2(n_344), .B1(n_1395), .B2(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1428 ( .A(n_324), .Y(n_1428) );
INVx1_ASAP7_75t_L g617 ( .A(n_325), .Y(n_617) );
INVx1_ASAP7_75t_L g720 ( .A(n_326), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g1593 ( .A1(n_329), .A2(n_372), .B1(n_1407), .B2(n_1594), .Y(n_1593) );
AOI22xp33_ASAP7_75t_L g1605 ( .A1(n_329), .A2(n_372), .B1(n_1189), .B2(n_1383), .Y(n_1605) );
CKINVDCx5p33_ASAP7_75t_R g1274 ( .A(n_330), .Y(n_1274) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_331), .Y(n_819) );
INVx1_ASAP7_75t_L g1332 ( .A(n_332), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_333), .Y(n_937) );
INVx1_ASAP7_75t_L g525 ( .A(n_334), .Y(n_525) );
INVx1_ASAP7_75t_L g1650 ( .A(n_335), .Y(n_1650) );
INVx1_ASAP7_75t_L g433 ( .A(n_336), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g1319 ( .A(n_337), .Y(n_1319) );
OAI22xp33_ASAP7_75t_L g1041 ( .A1(n_338), .A2(n_363), .B1(n_995), .B2(n_997), .Y(n_1041) );
INVx1_ASAP7_75t_L g1070 ( .A(n_338), .Y(n_1070) );
INVx1_ASAP7_75t_L g967 ( .A(n_341), .Y(n_967) );
INVx1_ASAP7_75t_L g1306 ( .A(n_342), .Y(n_1306) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_343), .Y(n_938) );
INVx1_ASAP7_75t_L g1420 ( .A(n_344), .Y(n_1420) );
INVx1_ASAP7_75t_L g1567 ( .A(n_345), .Y(n_1567) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_346), .B(n_381), .Y(n_1687) );
AND3x2_ASAP7_75t_L g1695 ( .A(n_346), .B(n_381), .C(n_1684), .Y(n_1695) );
INVx2_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_348), .Y(n_880) );
INVx1_ASAP7_75t_L g940 ( .A(n_349), .Y(n_940) );
AOI21xp33_ASAP7_75t_L g960 ( .A1(n_349), .A2(n_623), .B(n_961), .Y(n_960) );
OAI221xp5_ASAP7_75t_L g1163 ( .A1(n_350), .A2(n_485), .B1(n_512), .B2(n_1164), .C(n_1170), .Y(n_1163) );
INVx1_ASAP7_75t_L g922 ( .A(n_351), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g1437 ( .A(n_352), .Y(n_1437) );
INVx1_ASAP7_75t_L g1323 ( .A(n_353), .Y(n_1323) );
INVx1_ASAP7_75t_L g1287 ( .A(n_354), .Y(n_1287) );
INVx1_ASAP7_75t_L g1387 ( .A(n_355), .Y(n_1387) );
INVx1_ASAP7_75t_L g1017 ( .A(n_356), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g782 ( .A1(n_357), .A2(n_359), .B1(n_783), .B2(n_788), .C(n_791), .Y(n_782) );
OAI221xp5_ASAP7_75t_L g834 ( .A1(n_357), .A2(n_359), .B1(n_835), .B2(n_838), .C(n_840), .Y(n_834) );
INVx1_ASAP7_75t_L g396 ( .A(n_358), .Y(n_396) );
INVx2_ASAP7_75t_L g488 ( .A(n_358), .Y(n_488) );
AO22x2_ASAP7_75t_L g674 ( .A1(n_360), .A2(n_675), .B1(n_760), .B2(n_761), .Y(n_674) );
INVxp67_ASAP7_75t_SL g760 ( .A(n_360), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g1480 ( .A(n_361), .Y(n_1480) );
INVx1_ASAP7_75t_L g1111 ( .A(n_362), .Y(n_1111) );
INVx1_ASAP7_75t_L g1069 ( .A(n_363), .Y(n_1069) );
INVx1_ASAP7_75t_L g1555 ( .A(n_366), .Y(n_1555) );
HB1xp67_ASAP7_75t_L g1570 ( .A(n_366), .Y(n_1570) );
OAI211xp5_ASAP7_75t_L g1498 ( .A1(n_367), .A2(n_1439), .B(n_1499), .C(n_1501), .Y(n_1498) );
INVx1_ASAP7_75t_L g1530 ( .A(n_367), .Y(n_1530) );
INVxp33_ASAP7_75t_SL g1078 ( .A(n_368), .Y(n_1078) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_369), .B(n_643), .Y(n_642) );
OAI211xp5_ASAP7_75t_SL g1289 ( .A1(n_370), .A2(n_516), .B(n_1290), .C(n_1299), .Y(n_1289) );
INVxp33_ASAP7_75t_SL g1094 ( .A(n_371), .Y(n_1094) );
CKINVDCx5p33_ASAP7_75t_R g1162 ( .A(n_373), .Y(n_1162) );
INVx1_ASAP7_75t_L g1006 ( .A(n_374), .Y(n_1006) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_397), .B(n_1670), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
AND2x4_ASAP7_75t_L g1976 ( .A(n_379), .B(n_385), .Y(n_1976) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_SL g1970 ( .A(n_380), .Y(n_1970) );
NAND2xp5_ASAP7_75t_L g2026 ( .A(n_380), .B(n_382), .Y(n_2026) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g1969 ( .A(n_382), .B(n_1970), .Y(n_1969) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x6_ASAP7_75t_L g1353 ( .A(n_387), .B(n_469), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1478 ( .A(n_387), .B(n_469), .Y(n_1478) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g511 ( .A(n_388), .B(n_396), .Y(n_511) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g623 ( .A(n_389), .B(n_624), .Y(n_623) );
INVx8_ASAP7_75t_L g1349 ( .A(n_390), .Y(n_1349) );
OR2x6_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .Y(n_390) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_391), .Y(n_508) );
INVx2_ASAP7_75t_SL g799 ( .A(n_391), .Y(n_799) );
OR2x2_ASAP7_75t_L g827 ( .A(n_391), .B(n_787), .Y(n_827) );
INVx1_ASAP7_75t_L g911 ( .A(n_391), .Y(n_911) );
BUFx2_ASAP7_75t_L g1058 ( .A(n_391), .Y(n_1058) );
INVx2_ASAP7_75t_SL g1093 ( .A(n_391), .Y(n_1093) );
OR2x6_ASAP7_75t_L g1352 ( .A(n_391), .B(n_1343), .Y(n_1352) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g482 ( .A(n_393), .B(n_394), .Y(n_482) );
INVx2_ASAP7_75t_L g495 ( .A(n_393), .Y(n_495) );
AND2x4_ASAP7_75t_L g499 ( .A(n_393), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g506 ( .A(n_393), .Y(n_506) );
INVx1_ASAP7_75t_L g522 ( .A(n_393), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_394), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g500 ( .A(n_394), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_394), .Y(n_505) );
INVx1_ASAP7_75t_L g544 ( .A(n_394), .Y(n_544) );
INVx1_ASAP7_75t_L g553 ( .A(n_394), .Y(n_553) );
AND2x4_ASAP7_75t_L g1338 ( .A(n_395), .B(n_544), .Y(n_1338) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_396), .B(n_1340), .Y(n_1339) );
OR2x2_ASAP7_75t_L g1452 ( .A(n_396), .B(n_1340), .Y(n_1452) );
XNOR2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_1139), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_1072), .B2(n_1138), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
XNOR2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_868), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_672), .B2(n_867), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_593), .B2(n_594), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND4xp75_ASAP7_75t_SL g406 ( .A(n_407), .B(n_465), .C(n_483), .D(n_561), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_440), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_425), .B1(n_426), .B2(n_433), .C(n_434), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g1272 ( .A1(n_409), .A2(n_426), .B1(n_1273), .B2(n_1274), .Y(n_1272) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g650 ( .A(n_410), .Y(n_650) );
INVx2_ASAP7_75t_L g996 ( .A(n_410), .Y(n_996) );
INVx1_ASAP7_75t_L g1182 ( .A(n_410), .Y(n_1182) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_411), .B(n_416), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g837 ( .A(n_412), .Y(n_837) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g736 ( .A(n_413), .Y(n_736) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g453 ( .A(n_414), .B(n_431), .Y(n_453) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g438 ( .A(n_415), .B(n_432), .Y(n_438) );
AND2x4_ASAP7_75t_L g458 ( .A(n_415), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
OR2x6_ASAP7_75t_L g427 ( .A(n_417), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g439 ( .A(n_417), .Y(n_439) );
OR2x2_ASAP7_75t_L g997 ( .A(n_417), .B(n_428), .Y(n_997) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_418), .B(n_423), .Y(n_417) );
AND2x2_ASAP7_75t_L g470 ( .A(n_418), .B(n_453), .Y(n_470) );
AND2x4_ASAP7_75t_L g836 ( .A(n_418), .B(n_837), .Y(n_836) );
AND2x2_ASAP7_75t_L g839 ( .A(n_418), .B(n_429), .Y(n_839) );
INVx1_ASAP7_75t_L g859 ( .A(n_418), .Y(n_859) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_418), .B(n_837), .Y(n_1128) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g592 ( .A(n_421), .B(n_566), .Y(n_592) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g565 ( .A(n_422), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g718 ( .A(n_422), .Y(n_718) );
INVx1_ASAP7_75t_L g723 ( .A(n_422), .Y(n_723) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_422), .Y(n_727) );
OR2x6_ASAP7_75t_L g823 ( .A(n_423), .B(n_529), .Y(n_823) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g447 ( .A(n_424), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g772 ( .A(n_424), .B(n_487), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_425), .A2(n_433), .B1(n_542), .B2(n_545), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_426), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g1181 ( .A1(n_426), .A2(n_1161), .B1(n_1162), .B2(n_1182), .Y(n_1181) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g1129 ( .A(n_428), .B(n_859), .Y(n_1129) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x6_ASAP7_75t_L g737 ( .A(n_430), .B(n_723), .Y(n_737) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g444 ( .A(n_432), .B(n_445), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g872 ( .A(n_434), .B(n_873), .C(n_900), .Y(n_872) );
NOR3xp33_ASAP7_75t_L g933 ( .A(n_434), .B(n_934), .C(n_949), .Y(n_933) );
NOR3xp33_ASAP7_75t_SL g980 ( .A(n_434), .B(n_981), .C(n_994), .Y(n_980) );
NOR3xp33_ASAP7_75t_SL g1024 ( .A(n_434), .B(n_1025), .C(n_1041), .Y(n_1024) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_439), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g1212 ( .A(n_436), .Y(n_1212) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g740 ( .A(n_437), .B(n_741), .Y(n_740) );
BUFx6f_ASAP7_75t_L g851 ( .A(n_437), .Y(n_851) );
BUFx6f_ASAP7_75t_L g1383 ( .A(n_437), .Y(n_1383) );
INVx2_ASAP7_75t_L g1396 ( .A(n_437), .Y(n_1396) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_438), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_439), .B(n_648), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_449), .B1(n_450), .B2(n_454), .C(n_455), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_441), .A2(n_450), .B1(n_635), .B2(n_636), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g1202 ( .A1(n_441), .A2(n_450), .B1(n_1154), .B2(n_1158), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_441), .A2(n_450), .B1(n_1269), .B2(n_1270), .Y(n_1268) );
AOI222xp33_ASAP7_75t_L g1571 ( .A1(n_441), .A2(n_450), .B1(n_468), .B2(n_1546), .C1(n_1552), .C2(n_1572), .Y(n_1571) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_446), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g1417 ( .A(n_443), .Y(n_1417) );
OAI22xp5_ASAP7_75t_L g1519 ( .A1(n_443), .A2(n_1520), .B1(n_1521), .B2(n_1522), .Y(n_1519) );
INVx2_ASAP7_75t_SL g2020 ( .A(n_443), .Y(n_2020) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_444), .Y(n_576) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_444), .Y(n_586) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_444), .Y(n_657) );
AND2x6_ASAP7_75t_L g721 ( .A(n_444), .B(n_722), .Y(n_721) );
BUFx6f_ASAP7_75t_L g758 ( .A(n_444), .Y(n_758) );
BUFx3_ASAP7_75t_L g877 ( .A(n_444), .Y(n_877) );
BUFx2_ASAP7_75t_L g1278 ( .A(n_444), .Y(n_1278) );
BUFx2_ASAP7_75t_L g1604 ( .A(n_444), .Y(n_1604) );
INVx1_ASAP7_75t_L g464 ( .A(n_445), .Y(n_464) );
AND2x2_ASAP7_75t_L g450 ( .A(n_446), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g456 ( .A(n_447), .B(n_457), .Y(n_456) );
OR2x6_ASAP7_75t_L g460 ( .A(n_447), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g925 ( .A(n_447), .B(n_457), .Y(n_925) );
OR2x2_ASAP7_75t_L g927 ( .A(n_447), .B(n_928), .Y(n_927) );
OR2x2_ASAP7_75t_L g929 ( .A(n_447), .B(n_930), .Y(n_929) );
INVx2_ASAP7_75t_L g833 ( .A(n_448), .Y(n_833) );
OR2x2_ASAP7_75t_L g862 ( .A(n_448), .B(n_747), .Y(n_862) );
OR2x2_ASAP7_75t_L g864 ( .A(n_448), .B(n_865), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_449), .A2(n_533), .B1(n_536), .B2(n_540), .Y(n_532) );
INVx2_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g581 ( .A(n_452), .Y(n_581) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx6_ASAP7_75t_L g570 ( .A(n_453), .Y(n_570) );
AND2x4_ASAP7_75t_L g725 ( .A(n_453), .B(n_726), .Y(n_725) );
BUFx2_ASAP7_75t_L g1281 ( .A(n_453), .Y(n_1281) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_454), .A2(n_508), .B1(n_524), .B2(n_525), .C(n_526), .Y(n_523) );
CKINVDCx6p67_ASAP7_75t_R g639 ( .A(n_456), .Y(n_639) );
INVx2_ASAP7_75t_L g1957 ( .A(n_457), .Y(n_1957) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_458), .Y(n_579) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_458), .Y(n_589) );
INVx1_ASAP7_75t_L g670 ( .A(n_458), .Y(n_670) );
INVx2_ASAP7_75t_L g865 ( .A(n_458), .Y(n_865) );
INVx1_ASAP7_75t_L g463 ( .A(n_459), .Y(n_463) );
CKINVDCx6p67_ASAP7_75t_R g641 ( .A(n_460), .Y(n_641) );
BUFx3_ASAP7_75t_L g1517 ( .A(n_461), .Y(n_1517) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g756 ( .A(n_462), .Y(n_756) );
BUFx4f_ASAP7_75t_L g842 ( .A(n_462), .Y(n_842) );
BUFx2_ASAP7_75t_L g886 ( .A(n_462), .Y(n_886) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
OR2x2_ASAP7_75t_L g747 ( .A(n_463), .B(n_464), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g643 ( .A(n_467), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_467), .B(n_902), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_467), .B(n_951), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_467), .B(n_979), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_467), .B(n_1046), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_467), .B(n_1178), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_467), .B(n_1287), .Y(n_1286) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_471), .Y(n_467) );
INVx2_ASAP7_75t_L g828 ( .A(n_468), .Y(n_828) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
AND2x4_ASAP7_75t_L g591 ( .A(n_469), .B(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g899 ( .A(n_469), .B(n_592), .Y(n_899) );
NOR2xp67_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
INVx2_ASAP7_75t_L g1114 ( .A(n_472), .Y(n_1114) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OR2x6_ASAP7_75t_L g563 ( .A(n_473), .B(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g632 ( .A(n_473), .Y(n_632) );
OR2x2_ASAP7_75t_L g874 ( .A(n_473), .B(n_564), .Y(n_874) );
OAI31xp33_ASAP7_75t_L g1146 ( .A1(n_473), .A2(n_1147), .A3(n_1148), .B(n_1163), .Y(n_1146) );
AND2x4_ASAP7_75t_L g1357 ( .A(n_473), .B(n_511), .Y(n_1357) );
OR2x2_ASAP7_75t_L g1399 ( .A(n_473), .B(n_1400), .Y(n_1399) );
AND2x4_ASAP7_75t_L g1458 ( .A(n_473), .B(n_511), .Y(n_1458) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g560 ( .A(n_474), .Y(n_560) );
OR2x6_ASAP7_75t_L g796 ( .A(n_474), .B(n_623), .Y(n_796) );
INVx1_ASAP7_75t_L g679 ( .A(n_475), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .Y(n_475) );
AND2x2_ASAP7_75t_L g542 ( .A(n_476), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g921 ( .A(n_476), .B(n_543), .Y(n_921) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR2x6_ASAP7_75t_L g512 ( .A(n_477), .B(n_513), .Y(n_512) );
OR2x6_ASAP7_75t_L g546 ( .A(n_477), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g615 ( .A(n_477), .Y(n_615) );
OR2x2_ASAP7_75t_L g1061 ( .A(n_477), .B(n_513), .Y(n_1061) );
INVx1_ASAP7_75t_L g1557 ( .A(n_477), .Y(n_1557) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g1407 ( .A(n_480), .Y(n_1407) );
INVx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g606 ( .A(n_481), .Y(n_606) );
INVx2_ASAP7_75t_L g708 ( .A(n_481), .Y(n_708) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_482), .Y(n_489) );
OAI31xp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_515), .A3(n_548), .B(n_558), .Y(n_483) );
CKINVDCx6p67_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_486), .A2(n_620), .B1(n_625), .B2(n_629), .C(n_630), .Y(n_619) );
AOI222xp33_ASAP7_75t_L g677 ( .A1(n_486), .A2(n_517), .B1(n_678), .B2(n_679), .C1(n_680), .C2(n_681), .Y(n_677) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
INVx2_ASAP7_75t_L g519 ( .A(n_487), .Y(n_519) );
AND2x2_ASAP7_75t_L g550 ( .A(n_487), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g530 ( .A(n_488), .Y(n_530) );
INVx1_ASAP7_75t_L g624 ( .A(n_488), .Y(n_624) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_489), .Y(n_691) );
INVx3_ASAP7_75t_L g962 ( .A(n_489), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_496), .B1(n_497), .B2(n_501), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_491), .A2(n_628), .B1(n_878), .B2(n_880), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g1526 ( .A1(n_491), .A2(n_810), .B1(n_1503), .B2(n_1527), .Y(n_1526) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g1002 ( .A(n_492), .Y(n_1002) );
INVx2_ASAP7_75t_L g1011 ( .A(n_492), .Y(n_1011) );
INVx2_ASAP7_75t_L g1064 ( .A(n_492), .Y(n_1064) );
BUFx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g808 ( .A(n_493), .Y(n_808) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g535 ( .A(n_494), .Y(n_535) );
BUFx2_ASAP7_75t_L g694 ( .A(n_494), .Y(n_694) );
INVx1_ASAP7_75t_L g547 ( .A(n_495), .Y(n_547) );
AND2x4_ASAP7_75t_L g551 ( .A(n_495), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_SL g602 ( .A(n_498), .Y(n_602) );
INVx4_ASAP7_75t_L g628 ( .A(n_498), .Y(n_628) );
BUFx3_ASAP7_75t_L g815 ( .A(n_498), .Y(n_815) );
INVx2_ASAP7_75t_SL g916 ( .A(n_498), .Y(n_916) );
INVx2_ASAP7_75t_SL g966 ( .A(n_498), .Y(n_966) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx3_ASAP7_75t_L g539 ( .A(n_499), .Y(n_539) );
INVx1_ASAP7_75t_L g557 ( .A(n_499), .Y(n_557) );
INVx1_ASAP7_75t_L g1308 ( .A(n_499), .Y(n_1308) );
AND2x4_ASAP7_75t_L g521 ( .A(n_500), .B(n_522), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_507), .B1(n_508), .B2(n_509), .C(n_510), .Y(n_502) );
BUFx3_ASAP7_75t_L g689 ( .A(n_503), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g909 ( .A1(n_503), .A2(n_510), .B1(n_884), .B2(n_887), .C(n_910), .Y(n_909) );
BUFx3_ASAP7_75t_L g959 ( .A(n_503), .Y(n_959) );
INVx2_ASAP7_75t_L g1110 ( .A(n_503), .Y(n_1110) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_L g514 ( .A(n_505), .B(n_506), .Y(n_514) );
INVx1_ASAP7_75t_L g1340 ( .A(n_506), .Y(n_1340) );
BUFx2_ASAP7_75t_L g818 ( .A(n_508), .Y(n_818) );
INVx1_ASAP7_75t_L g1153 ( .A(n_508), .Y(n_1153) );
INVx1_ASAP7_75t_L g1175 ( .A(n_508), .Y(n_1175) );
OAI22xp33_ASAP7_75t_L g1524 ( .A1(n_508), .A2(n_1171), .B1(n_1514), .B2(n_1515), .Y(n_1524) );
OAI22xp33_ASAP7_75t_L g1528 ( .A1(n_508), .A2(n_1109), .B1(n_1529), .B2(n_1530), .Y(n_1528) );
BUFx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g1060 ( .A(n_511), .Y(n_1060) );
INVx2_ASAP7_75t_L g630 ( .A(n_512), .Y(n_630) );
HB1xp67_ASAP7_75t_L g1095 ( .A(n_513), .Y(n_1095) );
INVx1_ASAP7_75t_L g1172 ( .A(n_513), .Y(n_1172) );
NAND2xp5_ASAP7_75t_L g1553 ( .A(n_513), .B(n_1554), .Y(n_1553) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g524 ( .A(n_514), .Y(n_524) );
INVx2_ASAP7_75t_L g706 ( .A(n_514), .Y(n_706) );
BUFx2_ASAP7_75t_L g802 ( .A(n_514), .Y(n_802) );
INVx8_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_517), .A2(n_599), .B1(n_603), .B2(n_610), .C(n_611), .Y(n_598) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
AND2x4_ASAP7_75t_L g555 ( .A(n_518), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g1297 ( .A(n_520), .Y(n_1297) );
BUFx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_521), .Y(n_609) );
BUFx3_ASAP7_75t_L g775 ( .A(n_521), .Y(n_775) );
BUFx6f_ASAP7_75t_L g1331 ( .A(n_521), .Y(n_1331) );
AND2x4_ASAP7_75t_L g1333 ( .A(n_521), .B(n_1334), .Y(n_1333) );
BUFx2_ASAP7_75t_L g1648 ( .A(n_521), .Y(n_1648) );
OAI221xp5_ASAP7_75t_L g1055 ( .A1(n_524), .A2(n_1032), .B1(n_1033), .B2(n_1056), .C(n_1059), .Y(n_1055) );
OAI21xp5_ASAP7_75t_L g1542 ( .A1(n_524), .A2(n_1543), .B(n_1544), .Y(n_1542) );
OAI221xp5_ASAP7_75t_L g1149 ( .A1(n_526), .A2(n_1150), .B1(n_1151), .B2(n_1152), .C(n_1154), .Y(n_1149) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g709 ( .A(n_529), .Y(n_709) );
NAND2x1p5_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g1335 ( .A(n_530), .Y(n_1335) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_L g1291 ( .A(n_534), .Y(n_1291) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g914 ( .A(n_535), .Y(n_914) );
INVx2_ASAP7_75t_L g1157 ( .A(n_535), .Y(n_1157) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_SL g811 ( .A(n_538), .Y(n_811) );
INVx2_ASAP7_75t_L g1005 ( .A(n_538), .Y(n_1005) );
INVx2_ASAP7_75t_L g1105 ( .A(n_538), .Y(n_1105) );
INVx2_ASAP7_75t_L g1168 ( .A(n_538), .Y(n_1168) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx3_ASAP7_75t_L g697 ( .A(n_539), .Y(n_697) );
INVx3_ASAP7_75t_L g1054 ( .A(n_539), .Y(n_1054) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_542), .A2(n_545), .B1(n_700), .B2(n_701), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_542), .A2(n_545), .B1(n_1016), .B2(n_1017), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_542), .A2(n_545), .B1(n_1161), .B2(n_1162), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1299 ( .A1(n_542), .A2(n_545), .B1(n_1273), .B2(n_1274), .Y(n_1299) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g614 ( .A(n_544), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g1554 ( .A1(n_544), .A2(n_790), .B1(n_1555), .B2(n_1556), .Y(n_1554) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_545), .A2(n_920), .B1(n_921), .B2(n_922), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_545), .A2(n_921), .B1(n_970), .B2(n_971), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_545), .A2(n_921), .B1(n_1069), .B2(n_1070), .Y(n_1068) );
CKINVDCx11_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g790 ( .A(n_547), .Y(n_790) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_550), .A2(n_555), .B1(n_617), .B2(n_618), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_550), .A2(n_555), .B1(n_683), .B2(n_684), .Y(n_682) );
INVx3_ASAP7_75t_L g905 ( .A(n_550), .Y(n_905) );
BUFx2_ASAP7_75t_L g600 ( .A(n_551), .Y(n_600) );
BUFx2_ASAP7_75t_L g626 ( .A(n_551), .Y(n_626) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_551), .Y(n_781) );
AND2x4_ASAP7_75t_L g1342 ( .A(n_551), .B(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1404 ( .A(n_551), .Y(n_1404) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx3_ASAP7_75t_L g906 ( .A(n_555), .Y(n_906) );
INVx1_ASAP7_75t_L g1294 ( .A(n_556), .Y(n_1294) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI31xp33_ASAP7_75t_L g903 ( .A1(n_558), .A2(n_904), .A3(n_907), .B(n_912), .Y(n_903) );
OAI31xp33_ASAP7_75t_L g952 ( .A1(n_558), .A2(n_953), .A3(n_954), .B(n_963), .Y(n_952) );
OAI31xp33_ASAP7_75t_L g998 ( .A1(n_558), .A2(n_999), .A3(n_1000), .B(n_1009), .Y(n_998) );
BUFx8_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g1208 ( .A(n_559), .Y(n_1208) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g711 ( .A(n_560), .B(n_712), .Y(n_711) );
AND2x4_ASAP7_75t_L g1447 ( .A(n_560), .B(n_712), .Y(n_1447) );
AOI33xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_567), .A3(n_573), .B1(n_580), .B2(n_583), .B3(n_590), .Y(n_561) );
AOI33xp33_ASAP7_75t_L g1183 ( .A1(n_562), .A2(n_1184), .A3(n_1188), .B1(n_1192), .B2(n_1195), .B3(n_1198), .Y(n_1183) );
AOI33xp33_ASAP7_75t_L g2009 ( .A1(n_562), .A2(n_591), .A3(n_2010), .B1(n_2014), .B2(n_2019), .B3(n_2021), .Y(n_2009) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_563), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_563), .A2(n_743), .B1(n_753), .B2(n_759), .Y(n_742) );
INVx2_ASAP7_75t_L g1276 ( .A(n_563), .Y(n_1276) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx3_ASAP7_75t_L g853 ( .A(n_565), .Y(n_853) );
INVx1_ASAP7_75t_L g1133 ( .A(n_565), .Y(n_1133) );
INVx2_ASAP7_75t_SL g1227 ( .A(n_565), .Y(n_1227) );
INVx1_ASAP7_75t_L g1400 ( .A(n_565), .Y(n_1400) );
INVx1_ASAP7_75t_L g712 ( .A(n_566), .Y(n_712) );
BUFx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g1135 ( .A(n_569), .Y(n_1135) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g662 ( .A(n_570), .Y(n_662) );
INVx2_ASAP7_75t_L g719 ( .A(n_570), .Y(n_719) );
INVx2_ASAP7_75t_SL g845 ( .A(n_570), .Y(n_845) );
INVx2_ASAP7_75t_L g1190 ( .A(n_570), .Y(n_1190) );
BUFx6f_ASAP7_75t_L g1194 ( .A(n_570), .Y(n_1194) );
HB1xp67_ASAP7_75t_L g1563 ( .A(n_570), .Y(n_1563) );
INVx1_ASAP7_75t_L g1664 ( .A(n_570), .Y(n_1664) );
AOI222xp33_ASAP7_75t_L g1321 ( .A1(n_571), .A2(n_737), .B1(n_1322), .B2(n_1323), .C1(n_1324), .C2(n_1326), .Y(n_1321) );
BUFx4f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx3_ASAP7_75t_L g582 ( .A(n_572), .Y(n_582) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_572), .Y(n_648) );
INVx2_ASAP7_75t_SL g664 ( .A(n_572), .Y(n_664) );
INVx1_ASAP7_75t_L g732 ( .A(n_572), .Y(n_732) );
AND2x4_ASAP7_75t_L g856 ( .A(n_572), .B(n_833), .Y(n_856) );
INVx1_ASAP7_75t_L g1608 ( .A(n_572), .Y(n_1608) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_575), .A2(n_895), .B1(n_1038), .B2(n_1039), .Y(n_1037) );
INVx1_ASAP7_75t_L g1217 ( .A(n_575), .Y(n_1217) );
INVx1_ASAP7_75t_L g1465 ( .A(n_575), .Y(n_1465) );
OAI22xp5_ASAP7_75t_L g1564 ( .A1(n_575), .A2(n_670), .B1(n_1539), .B2(n_1541), .Y(n_1564) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
BUFx3_ASAP7_75t_L g668 ( .A(n_576), .Y(n_668) );
AND2x4_ASAP7_75t_L g832 ( .A(n_576), .B(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g1123 ( .A(n_576), .Y(n_1123) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_579), .Y(n_658) );
INVx1_ASAP7_75t_L g879 ( .A(n_579), .Y(n_879) );
INVx1_ASAP7_75t_L g1029 ( .A(n_579), .Y(n_1029) );
BUFx3_ASAP7_75t_L g1229 ( .A(n_579), .Y(n_1229) );
AOI222xp33_ASAP7_75t_L g1989 ( .A1(n_582), .A2(n_737), .B1(n_1324), .B2(n_1990), .C1(n_1991), .C2(n_1992), .Y(n_1989) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g752 ( .A(n_585), .Y(n_752) );
INVx1_ASAP7_75t_L g1196 ( .A(n_585), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1566 ( .A1(n_585), .A2(n_1187), .B1(n_1567), .B2(n_1568), .Y(n_1566) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g893 ( .A(n_586), .Y(n_893) );
INVx2_ASAP7_75t_SL g936 ( .A(n_586), .Y(n_936) );
AOI322xp5_ASAP7_75t_L g1501 ( .A1(n_586), .A2(n_737), .A3(n_1490), .B1(n_1494), .B2(n_1502), .C1(n_1503), .C2(n_1504), .Y(n_1501) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g1371 ( .A(n_588), .Y(n_1371) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x6_ASAP7_75t_L g729 ( .A(n_589), .B(n_717), .Y(n_729) );
BUFx6f_ASAP7_75t_L g896 ( .A(n_589), .Y(n_896) );
BUFx6f_ASAP7_75t_L g993 ( .A(n_589), .Y(n_993) );
HB1xp67_ASAP7_75t_L g1197 ( .A(n_589), .Y(n_1197) );
INVx1_ASAP7_75t_L g1522 ( .A(n_589), .Y(n_1522) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_590), .Y(n_759) );
BUFx4f_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx4f_ASAP7_75t_L g671 ( .A(n_591), .Y(n_671) );
INVx4_ASAP7_75t_L g1040 ( .A(n_591), .Y(n_1040) );
AOI33xp33_ASAP7_75t_L g1463 ( .A1(n_591), .A2(n_654), .A3(n_1464), .B1(n_1466), .B2(n_1467), .B3(n_1469), .Y(n_1463) );
AOI221xp5_ASAP7_75t_L g1560 ( .A1(n_591), .A2(n_1276), .B1(n_1561), .B2(n_1565), .C(n_1569), .Y(n_1560) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_592), .Y(n_846) );
INVx2_ASAP7_75t_SL g1120 ( .A(n_592), .Y(n_1120) );
INVx2_ASAP7_75t_L g1215 ( .A(n_592), .Y(n_1215) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
XNOR2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NOR4xp75_ASAP7_75t_L g596 ( .A(n_597), .B(n_633), .C(n_642), .D(n_644), .Y(n_596) );
AOI31xp33_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_616), .A3(n_619), .B(n_631), .Y(n_597) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g621 ( .A(n_606), .Y(n_621) );
AND2x4_ASAP7_75t_L g778 ( .A(n_606), .B(n_772), .Y(n_778) );
AOI211xp5_ASAP7_75t_L g1419 ( .A1(n_607), .A2(n_1333), .B(n_1420), .C(n_1421), .Y(n_1419) );
INVx2_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g622 ( .A(n_608), .Y(n_622) );
INVx2_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
BUFx6f_ASAP7_75t_L g1594 ( .A(n_609), .Y(n_1594) );
NAND2x1p5_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
NAND2x1_ASAP7_75t_SL g785 ( .A(n_613), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI222xp33_ASAP7_75t_L g1586 ( .A1(n_622), .A2(n_1491), .B1(n_1587), .B2(n_1588), .C1(n_1589), .C2(n_1590), .Y(n_1586) );
INVx1_ASAP7_75t_L g1343 ( .A(n_624), .Y(n_1343) );
INVx2_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g703 ( .A(n_628), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g1010 ( .A1(n_628), .A2(n_1011), .B1(n_1012), .B2(n_1013), .C(n_1014), .Y(n_1010) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_628), .A2(n_1064), .B1(n_1065), .B2(n_1066), .C(n_1067), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_628), .A2(n_1219), .B1(n_1233), .B2(n_1251), .Y(n_1255) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_630), .B(n_686), .C(n_702), .Y(n_685) );
INVx2_ASAP7_75t_L g866 ( .A(n_631), .Y(n_866) );
CKINVDCx8_ASAP7_75t_R g631 ( .A(n_632), .Y(n_631) );
AOI221x1_ASAP7_75t_SL g675 ( .A1(n_632), .A2(n_676), .B1(n_710), .B2(n_713), .C(n_742), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_637), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B1(n_640), .B2(n_641), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_639), .A2(n_641), .B1(n_1151), .B2(n_1159), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_639), .A2(n_641), .B1(n_1266), .B2(n_1267), .Y(n_1265) );
AOI22xp5_ASAP7_75t_L g1573 ( .A1(n_639), .A2(n_641), .B1(n_1547), .B2(n_1549), .Y(n_1573) );
NAND3xp33_ASAP7_75t_SL g644 ( .A(n_645), .B(n_649), .C(n_653), .Y(n_644) );
NAND3xp33_ASAP7_75t_SL g1180 ( .A(n_645), .B(n_1181), .C(n_1183), .Y(n_1180) );
NAND3xp33_ASAP7_75t_L g1271 ( .A(n_645), .B(n_1272), .C(n_1275), .Y(n_1271) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_648), .Y(n_666) );
BUFx2_ASAP7_75t_SL g1132 ( .A(n_648), .Y(n_1132) );
INVx1_ASAP7_75t_L g2018 ( .A(n_648), .Y(n_2018) );
AOI33xp33_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .A3(n_659), .B1(n_665), .B2(n_667), .B3(n_671), .Y(n_653) );
AOI33xp33_ASAP7_75t_L g1368 ( .A1(n_654), .A2(n_671), .A3(n_1369), .B1(n_1372), .B2(n_1373), .B3(n_1374), .Y(n_1368) );
BUFx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g1027 ( .A(n_657), .Y(n_1027) );
BUFx3_ASAP7_75t_L g1370 ( .A(n_657), .Y(n_1370) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_663), .B(n_1435), .Y(n_1434) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g1191 ( .A(n_664), .Y(n_1191) );
INVx1_ASAP7_75t_L g1282 ( .A(n_664), .Y(n_1282) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g750 ( .A(n_670), .Y(n_750) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_670), .A2(n_936), .B1(n_937), .B2(n_938), .Y(n_935) );
INVx1_ASAP7_75t_L g867 ( .A(n_672), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B1(n_762), .B2(n_763), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g761 ( .A(n_675), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_682), .C(n_685), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_678), .A2(n_725), .B1(n_728), .B2(n_729), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g753 ( .A1(n_680), .A2(n_681), .B1(n_745), .B2(n_754), .C(n_757), .Y(n_753) );
OAI21xp5_ASAP7_75t_SL g686 ( .A1(n_687), .A2(n_692), .B(n_699), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B(n_690), .Y(n_687) );
BUFx3_ASAP7_75t_L g1938 ( .A(n_689), .Y(n_1938) );
INVx1_ASAP7_75t_L g1366 ( .A(n_691), .Y(n_1366) );
A2O1A1Ixp33_ASAP7_75t_L g1551 ( .A1(n_691), .A2(n_1552), .B(n_1553), .C(n_1557), .Y(n_1551) );
HB1xp67_ASAP7_75t_L g2005 ( .A(n_691), .Y(n_2005) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .B1(n_696), .B2(n_698), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_693), .A2(n_1103), .B1(n_1104), .B2(n_1106), .Y(n_1102) );
BUFx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g957 ( .A(n_694), .Y(n_957) );
OR2x2_ASAP7_75t_L g1482 ( .A(n_694), .B(n_1483), .Y(n_1482) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_696), .A2(n_937), .B1(n_938), .B2(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_L g771 ( .A(n_697), .B(n_772), .Y(n_771) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_698), .A2(n_744), .B1(n_748), .B2(n_749), .C(n_751), .Y(n_743) );
AOI222xp33_ASAP7_75t_L g730 ( .A1(n_700), .A2(n_701), .B1(n_705), .B2(n_731), .C1(n_733), .C2(n_737), .Y(n_730) );
OAI21xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_706), .B(n_707), .Y(n_704) );
OAI21xp33_ASAP7_75t_L g1548 ( .A1(n_706), .A2(n_1549), .B(n_1550), .Y(n_1548) );
OAI22xp33_ASAP7_75t_L g1947 ( .A1(n_706), .A2(n_910), .B1(n_1948), .B2(n_1949), .Y(n_1947) );
BUFx3_ASAP7_75t_L g1359 ( .A(n_708), .Y(n_1359) );
AOI211x1_ASAP7_75t_L g1313 ( .A1(n_710), .A2(n_1314), .B(n_1327), .C(n_1354), .Y(n_1313) );
AOI221x1_ASAP7_75t_L g1626 ( .A1(n_710), .A2(n_1578), .B1(n_1627), .B2(n_1638), .C(n_1651), .Y(n_1626) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AO211x2_ASAP7_75t_L g1378 ( .A1(n_711), .A2(n_1379), .B(n_1392), .C(n_1418), .Y(n_1378) );
AOI221xp5_ASAP7_75t_L g1981 ( .A1(n_711), .A2(n_1578), .B1(n_1982), .B2(n_1993), .C(n_2002), .Y(n_1981) );
NAND4xp25_ASAP7_75t_SL g713 ( .A(n_714), .B(n_724), .C(n_730), .D(n_738), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_720), .B2(n_721), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_716), .A2(n_721), .B1(n_1316), .B2(n_1317), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_716), .A2(n_725), .B1(n_1387), .B2(n_1388), .Y(n_1386) );
AOI22xp33_ASAP7_75t_L g1628 ( .A1(n_716), .A2(n_729), .B1(n_1629), .B2(n_1630), .Y(n_1628) );
AND2x4_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
AND2x4_ASAP7_75t_L g1619 ( .A(n_717), .B(n_719), .Y(n_1619) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_718), .B(n_1616), .Y(n_1615) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_721), .A2(n_729), .B1(n_1390), .B2(n_1391), .Y(n_1389) );
CKINVDCx6p67_ASAP7_75t_R g1441 ( .A(n_721), .Y(n_1441) );
AOI22xp33_ASAP7_75t_L g1620 ( .A1(n_721), .A2(n_729), .B1(n_1621), .B2(n_1622), .Y(n_1620) );
AOI221xp5_ASAP7_75t_L g1631 ( .A1(n_721), .A2(n_725), .B1(n_1632), .B2(n_1633), .C(n_1634), .Y(n_1631) );
AOI22xp33_ASAP7_75t_L g1983 ( .A1(n_721), .A2(n_1619), .B1(n_1984), .B2(n_1985), .Y(n_1983) );
INVx1_ASAP7_75t_L g741 ( .A(n_722), .Y(n_741) );
INVx1_ASAP7_75t_L g1445 ( .A(n_722), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_722), .B(n_1383), .Y(n_1500) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_725), .A2(n_729), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
INVx4_ASAP7_75t_L g1446 ( .A(n_725), .Y(n_1446) );
AOI22xp33_ASAP7_75t_L g1617 ( .A1(n_725), .A2(n_1585), .B1(n_1618), .B2(n_1619), .Y(n_1617) );
AOI22xp33_ASAP7_75t_L g1986 ( .A1(n_725), .A2(n_729), .B1(n_1987), .B2(n_1988), .Y(n_1986) );
AND2x4_ASAP7_75t_L g734 ( .A(n_726), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_SL g1504 ( .A(n_726), .B(n_735), .Y(n_1504) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx4_ASAP7_75t_L g1442 ( .A(n_729), .Y(n_1442) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx4f_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g1325 ( .A(n_734), .Y(n_1325) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_734), .A2(n_737), .B1(n_1437), .B2(n_1438), .Y(n_1436) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g1616 ( .A(n_736), .Y(n_1616) );
INVx3_ASAP7_75t_L g1385 ( .A(n_737), .Y(n_1385) );
BUFx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND4xp25_ASAP7_75t_SL g1314 ( .A(n_739), .B(n_1315), .C(n_1318), .D(n_1321), .Y(n_1314) );
NAND4xp25_ASAP7_75t_L g1982 ( .A(n_739), .B(n_1983), .C(n_1986), .D(n_1989), .Y(n_1982) );
INVx5_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI211xp5_ASAP7_75t_L g1380 ( .A1(n_740), .A2(n_1381), .B(n_1382), .C(n_1384), .Y(n_1380) );
CKINVDCx8_ASAP7_75t_R g1439 ( .A(n_740), .Y(n_1439) );
AOI211xp5_ASAP7_75t_L g1611 ( .A1(n_740), .A2(n_1500), .B(n_1612), .C(n_1613), .Y(n_1611) );
OAI21xp33_ASAP7_75t_L g1636 ( .A1(n_741), .A2(n_851), .B(n_1637), .Y(n_1636) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g883 ( .A(n_747), .Y(n_883) );
BUFx2_ASAP7_75t_L g983 ( .A(n_747), .Y(n_983) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_747), .B(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_754), .A2(n_943), .B1(n_944), .B2(n_945), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g1031 ( .A1(n_754), .A2(n_882), .B1(n_1032), .B2(n_1033), .Y(n_1031) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
BUFx2_ASAP7_75t_L g990 ( .A(n_756), .Y(n_990) );
INVx1_ASAP7_75t_L g930 ( .A(n_758), .Y(n_930) );
BUFx4f_ASAP7_75t_L g1185 ( .A(n_758), .Y(n_1185) );
BUFx2_ASAP7_75t_L g1375 ( .A(n_758), .Y(n_1375) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_759), .A2(n_874), .B1(n_982), .B2(n_988), .Y(n_981) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
XNOR2x1_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_824), .Y(n_765) );
NOR3xp33_ASAP7_75t_SL g766 ( .A(n_767), .B(n_782), .C(n_793), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_776), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B1(n_773), .B2(n_774), .Y(n_768) );
BUFx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
BUFx2_ASAP7_75t_L g1079 ( .A(n_771), .Y(n_1079) );
BUFx2_ASAP7_75t_L g1239 ( .A(n_771), .Y(n_1239) );
AND2x6_ASAP7_75t_L g774 ( .A(n_772), .B(n_775), .Y(n_774) );
AND2x2_ASAP7_75t_L g780 ( .A(n_772), .B(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_772), .B(n_781), .Y(n_1084) );
OAI211xp5_ASAP7_75t_L g840 ( .A1(n_773), .A2(n_841), .B(n_843), .C(n_844), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_774), .A2(n_1078), .B1(n_1079), .B2(n_1080), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_774), .A2(n_1238), .B1(n_1239), .B2(n_1240), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1926 ( .A1(n_774), .A2(n_1239), .B1(n_1927), .B2(n_1928), .Y(n_1926) );
NAND2x1p5_ASAP7_75t_L g792 ( .A(n_775), .B(n_786), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_778), .A2(n_1082), .B1(n_1083), .B2(n_1084), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_778), .A2(n_1084), .B1(n_1242), .B2(n_1243), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g1929 ( .A1(n_778), .A2(n_1084), .B1(n_1930), .B2(n_1931), .Y(n_1929) );
INVx2_ASAP7_75t_SL g1363 ( .A(n_781), .Y(n_1363) );
INVx2_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NAND2x1p5_ASAP7_75t_L g789 ( .A(n_786), .B(n_790), .Y(n_789) );
INVx3_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
BUFx4f_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
BUFx4f_ASAP7_75t_L g1086 ( .A(n_789), .Y(n_1086) );
BUFx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx2_ASAP7_75t_L g1087 ( .A(n_792), .Y(n_1087) );
OAI33xp33_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_797), .A3(n_804), .B1(n_812), .B2(n_817), .B3(n_821), .Y(n_793) );
OAI33xp33_ASAP7_75t_L g1245 ( .A1(n_794), .A2(n_821), .A3(n_1246), .B1(n_1250), .B2(n_1255), .B3(n_1256), .Y(n_1245) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OAI33xp33_ASAP7_75t_L g1088 ( .A1(n_796), .A2(n_821), .A3(n_1089), .B1(n_1096), .B2(n_1102), .B3(n_1107), .Y(n_1088) );
OAI33xp33_ASAP7_75t_L g1523 ( .A1(n_796), .A2(n_1524), .A3(n_1525), .B1(n_1526), .B2(n_1528), .B3(n_1531), .Y(n_1523) );
OAI33xp33_ASAP7_75t_L g1933 ( .A1(n_796), .A2(n_821), .A3(n_1934), .B1(n_1939), .B2(n_1944), .B3(n_1947), .Y(n_1933) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_800), .B1(n_801), .B2(n_803), .Y(n_797) );
INVx3_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g817 ( .A1(n_801), .A2(n_818), .B1(n_819), .B2(n_820), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g1301 ( .A1(n_801), .A2(n_1059), .B1(n_1152), .B2(n_1302), .C(n_1303), .Y(n_1301) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_809), .B2(n_810), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_806), .A2(n_813), .B1(n_814), .B2(n_816), .Y(n_812) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx2_ASAP7_75t_L g1165 ( .A(n_808), .Y(n_1165) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g831 ( .A1(n_813), .A2(n_832), .B(n_834), .Y(n_831) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_816), .A2(n_819), .B1(n_861), .B2(n_863), .Y(n_860) );
AOI221xp5_ASAP7_75t_L g847 ( .A1(n_820), .A2(n_848), .B1(n_854), .B2(n_855), .C(n_857), .Y(n_847) );
CKINVDCx8_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
NAND3xp33_ASAP7_75t_L g1401 ( .A(n_822), .B(n_1402), .C(n_1406), .Y(n_1401) );
NAND3xp33_ASAP7_75t_L g1656 ( .A(n_822), .B(n_1657), .C(n_1658), .Y(n_1656) );
INVx5_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx6_ASAP7_75t_L g1367 ( .A(n_823), .Y(n_1367) );
AOI21xp33_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_829), .B(n_830), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_825), .A2(n_1113), .B1(n_1115), .B2(n_1137), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_825), .A2(n_1208), .B1(n_1209), .B2(n_1234), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1950 ( .A1(n_825), .A2(n_1113), .B1(n_1951), .B2(n_1963), .Y(n_1950) );
INVx5_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AND2x4_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
AOI31xp33_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_847), .A3(n_860), .B(n_866), .Y(n_830) );
AOI221xp5_ASAP7_75t_L g1116 ( .A1(n_832), .A2(n_1103), .B1(n_1117), .B2(n_1121), .C(n_1126), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1210 ( .A1(n_832), .A2(n_1211), .B1(n_1216), .B2(n_1219), .C(n_1220), .Y(n_1210) );
AOI221xp5_ASAP7_75t_L g1952 ( .A1(n_832), .A2(n_1945), .B1(n_1953), .B2(n_1955), .C(n_1958), .Y(n_1952) );
INVx1_ASAP7_75t_SL g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_SL g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g890 ( .A(n_842), .Y(n_890) );
INVx1_ASAP7_75t_L g985 ( .A(n_842), .Y(n_985) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
AND2x4_ASAP7_75t_L g857 ( .A(n_851), .B(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g1224 ( .A(n_851), .Y(n_1224) );
BUFx6f_ASAP7_75t_L g1468 ( .A(n_851), .Y(n_1468) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
AOI221xp5_ASAP7_75t_L g1130 ( .A1(n_855), .A2(n_857), .B1(n_1111), .B2(n_1131), .C(n_1134), .Y(n_1130) );
AOI221xp5_ASAP7_75t_L g1221 ( .A1(n_855), .A2(n_857), .B1(n_1222), .B2(n_1228), .C(n_1230), .Y(n_1221) );
AOI221xp5_ASAP7_75t_L g1959 ( .A1(n_855), .A2(n_857), .B1(n_1949), .B2(n_1960), .C(n_1961), .Y(n_1959) );
BUFx6f_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_SL g858 ( .A(n_859), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_861), .A2(n_863), .B1(n_1106), .B2(n_1108), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_861), .A2(n_863), .B1(n_1232), .B2(n_1233), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g1962 ( .A1(n_861), .A2(n_863), .B1(n_1946), .B2(n_1948), .Y(n_1962) );
INVx6_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx4_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g1125 ( .A(n_865), .Y(n_1125) );
INVx1_ASAP7_75t_L g1512 ( .A(n_865), .Y(n_1512) );
OAI31xp33_ASAP7_75t_L g1047 ( .A1(n_866), .A2(n_1048), .A3(n_1049), .B(n_1062), .Y(n_1047) );
OAI31xp33_ASAP7_75t_L g1288 ( .A1(n_866), .A2(n_1289), .A3(n_1300), .B(n_1309), .Y(n_1288) );
XNOR2xp5_ASAP7_75t_L g868 ( .A(n_869), .B(n_975), .Y(n_868) );
XOR2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_931), .Y(n_869) );
AND4x1_ASAP7_75t_L g871 ( .A(n_872), .B(n_901), .C(n_903), .D(n_923), .Y(n_871) );
OAI33xp33_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_875), .A3(n_881), .B1(n_888), .B2(n_892), .B3(n_898), .Y(n_873) );
OAI33xp33_ASAP7_75t_L g934 ( .A1(n_874), .A2(n_898), .A3(n_935), .B1(n_939), .B2(n_942), .B3(n_946), .Y(n_934) );
OAI33xp33_ASAP7_75t_L g1025 ( .A1(n_874), .A2(n_1026), .A3(n_1031), .B1(n_1034), .B2(n_1037), .B3(n_1040), .Y(n_1025) );
OAI33xp33_ASAP7_75t_L g1506 ( .A1(n_874), .A2(n_1040), .A3(n_1507), .B1(n_1513), .B2(n_1516), .B3(n_1519), .Y(n_1506) );
INVx1_ASAP7_75t_SL g1602 ( .A(n_874), .Y(n_1602) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_875) );
INVx2_ASAP7_75t_SL g876 ( .A(n_877), .Y(n_876) );
BUFx3_ASAP7_75t_L g2011 ( .A(n_877), .Y(n_2011) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_879), .A2(n_893), .B1(n_947), .B2(n_948), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_884), .B1(n_885), .B2(n_887), .Y(n_881) );
OAI22xp33_ASAP7_75t_L g888 ( .A1(n_882), .A2(n_889), .B1(n_890), .B2(n_891), .Y(n_888) );
OAI22xp33_ASAP7_75t_L g939 ( .A1(n_882), .A2(n_885), .B1(n_940), .B2(n_941), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g1034 ( .A1(n_882), .A2(n_985), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
OAI22xp33_ASAP7_75t_SL g1513 ( .A1(n_882), .A2(n_990), .B1(n_1514), .B2(n_1515), .Y(n_1513) );
OAI22xp33_ASAP7_75t_L g1516 ( .A1(n_882), .A2(n_1480), .B1(n_1517), .B2(n_1518), .Y(n_1516) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g928 ( .A(n_883), .Y(n_928) );
INVx2_ASAP7_75t_L g943 ( .A(n_883), .Y(n_943) );
INVx2_ASAP7_75t_SL g885 ( .A(n_886), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_894), .B1(n_895), .B2(n_897), .Y(n_892) );
INVx2_ASAP7_75t_SL g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g1199 ( .A(n_899), .Y(n_1199) );
AOI33xp33_ASAP7_75t_L g1275 ( .A1(n_899), .A2(n_1276), .A3(n_1277), .B1(n_1280), .B2(n_1283), .B3(n_1284), .Y(n_1275) );
NAND3xp33_ASAP7_75t_L g1413 ( .A(n_899), .B(n_1414), .C(n_1416), .Y(n_1413) );
AOI33xp33_ASAP7_75t_L g1601 ( .A1(n_899), .A2(n_1602), .A3(n_1603), .B1(n_1605), .B2(n_1606), .B3(n_1609), .Y(n_1601) );
NAND3xp33_ASAP7_75t_L g1662 ( .A(n_899), .B(n_1663), .C(n_1665), .Y(n_1662) );
OAI22xp33_ASAP7_75t_L g1246 ( .A1(n_910), .A2(n_1247), .B1(n_1248), .B2(n_1249), .Y(n_1246) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g1936 ( .A(n_911), .Y(n_1936) );
OAI221xp5_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_915), .B1(n_916), .B2(n_917), .C(n_918), .Y(n_913) );
OAI221xp5_ASAP7_75t_L g964 ( .A1(n_914), .A2(n_965), .B1(n_966), .B2(n_967), .C(n_968), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g1155 ( .A1(n_916), .A2(n_1156), .B1(n_1158), .B2(n_1159), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_916), .A2(n_1251), .B1(n_1253), .B2(n_1254), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1944 ( .A1(n_916), .A2(n_1251), .B1(n_1945), .B2(n_1946), .Y(n_1944) );
NOR2xp33_ASAP7_75t_L g923 ( .A(n_924), .B(n_926), .Y(n_923) );
AND4x1_ASAP7_75t_L g932 ( .A(n_933), .B(n_950), .C(n_952), .D(n_972), .Y(n_932) );
OAI21xp33_ASAP7_75t_SL g958 ( .A1(n_941), .A2(n_959), .B(n_960), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g1525 ( .A1(n_956), .A2(n_1294), .B1(n_1508), .B2(n_1510), .Y(n_1525) );
INVx2_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
OAI21xp33_ASAP7_75t_L g1007 ( .A1(n_959), .A2(n_986), .B(n_1008), .Y(n_1007) );
OAI22xp33_ASAP7_75t_L g1256 ( .A1(n_959), .A2(n_1091), .B1(n_1230), .B2(n_1232), .Y(n_1256) );
INVx2_ASAP7_75t_SL g961 ( .A(n_962), .Y(n_961) );
INVx2_ASAP7_75t_L g1298 ( .A(n_962), .Y(n_1298) );
INVx2_ASAP7_75t_L g1488 ( .A(n_962), .Y(n_1488) );
NOR2xp33_ASAP7_75t_L g972 ( .A(n_973), .B(n_974), .Y(n_972) );
AO22x2_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_1021), .B1(n_1022), .B2(n_1071), .Y(n_975) );
INVx1_ASAP7_75t_L g1071 ( .A(n_976), .Y(n_1071) );
AND4x1_ASAP7_75t_L g977 ( .A(n_978), .B(n_980), .C(n_998), .D(n_1018), .Y(n_977) );
OAI221xp5_ASAP7_75t_L g982 ( .A1(n_983), .A2(n_984), .B1(n_985), .B2(n_986), .C(n_987), .Y(n_982) );
OAI221xp5_ASAP7_75t_L g988 ( .A1(n_983), .A2(n_989), .B1(n_990), .B2(n_991), .C(n_992), .Y(n_988) );
INVx1_ASAP7_75t_L g2013 ( .A(n_993), .Y(n_2013) );
INVx2_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1003), .B1(n_1004), .B2(n_1006), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_1002), .A2(n_1028), .B1(n_1030), .B2(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1011), .Y(n_1252) );
NOR2xp33_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1020), .Y(n_1018) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
AND4x1_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1042), .C(n_1045), .D(n_1047), .Y(n_1023) );
OAI22xp33_ASAP7_75t_L g1026 ( .A1(n_1027), .A2(n_1028), .B1(n_1029), .B2(n_1030), .Y(n_1026) );
NOR2xp33_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1044), .Y(n_1042) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx2_ASAP7_75t_L g1405 ( .A(n_1053), .Y(n_1405) );
OAI22xp5_ASAP7_75t_L g1545 ( .A1(n_1053), .A2(n_1157), .B1(n_1546), .B2(n_1547), .Y(n_1545) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1053), .Y(n_1596) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1054), .Y(n_1101) );
INVx2_ASAP7_75t_L g1540 ( .A(n_1054), .Y(n_1540) );
INVx2_ASAP7_75t_SL g1056 ( .A(n_1057), .Y(n_1056) );
INVx2_ASAP7_75t_SL g1057 ( .A(n_1058), .Y(n_1057) );
OAI221xp5_ASAP7_75t_L g1170 ( .A1(n_1059), .A2(n_1171), .B1(n_1173), .B2(n_1174), .C(n_1176), .Y(n_1170) );
INVx2_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_1064), .A2(n_1097), .B1(n_1098), .B2(n_1099), .Y(n_1096) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1072), .Y(n_1138) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1112), .Y(n_1074) );
NOR3xp33_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1085), .C(n_1088), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1081), .Y(n_1076) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_1090), .A2(n_1091), .B1(n_1094), .B2(n_1095), .Y(n_1089) );
OAI22xp33_ASAP7_75t_L g1107 ( .A1(n_1091), .A2(n_1108), .B1(n_1109), .B2(n_1111), .Y(n_1107) );
BUFx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx2_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx2_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1110), .Y(n_1150) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1110), .Y(n_1248) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
OAI31xp33_ASAP7_75t_L g1536 ( .A1(n_1114), .A2(n_1537), .A3(n_1558), .B(n_1559), .Y(n_1536) );
NAND3xp33_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1130), .C(n_1136), .Y(n_1115) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1218 ( .A(n_1124), .Y(n_1218) );
BUFx2_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1125), .Y(n_1187) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
XOR2xp5_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1257), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
AOI22x1_ASAP7_75t_L g1142 ( .A1(n_1143), .A2(n_1144), .B1(n_1203), .B2(n_1204), .Y(n_1142) );
INVx2_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
NAND3xp33_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1177), .C(n_1179), .Y(n_1145) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
BUFx2_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g1304 ( .A1(n_1157), .A2(n_1305), .B1(n_1306), .B2(n_1307), .Y(n_1304) );
OAI22xp5_ASAP7_75t_L g1538 ( .A1(n_1157), .A2(n_1539), .B1(n_1540), .B2(n_1541), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_1165), .A2(n_1166), .B1(n_1167), .B2(n_1169), .Y(n_1164) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
NOR2xp33_ASAP7_75t_SL g1179 ( .A(n_1180), .B(n_1200), .Y(n_1179) );
INVx2_ASAP7_75t_SL g1186 ( .A(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1187), .Y(n_1279) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1187), .Y(n_1285) );
BUFx6f_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g2016 ( .A(n_1190), .Y(n_2016) );
INVx4_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1194), .Y(n_1213) );
INVx2_ASAP7_75t_L g1415 ( .A(n_1194), .Y(n_1415) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1196), .Y(n_1509) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1202), .Y(n_1200) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
XNOR2x1_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1206), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1235), .Y(n_1206) );
NAND3xp33_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1221), .C(n_1231), .Y(n_1209) );
BUFx2_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
NOR3xp33_ASAP7_75t_SL g1235 ( .A(n_1236), .B(n_1244), .C(n_1245), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1241), .Y(n_1236) );
OAI22xp5_ASAP7_75t_L g1939 ( .A1(n_1251), .A2(n_1940), .B1(n_1941), .B2(n_1942), .Y(n_1939) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
AO22x2_ASAP7_75t_L g1257 ( .A1(n_1258), .A2(n_1472), .B1(n_1473), .B2(n_1669), .Y(n_1257) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1258), .Y(n_1669) );
XOR2xp5_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1310), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
NAND3xp33_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1286), .C(n_1288), .Y(n_1262) );
NOR2xp33_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1271), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1268), .Y(n_1264) );
OAI221xp5_ASAP7_75t_L g1290 ( .A1(n_1266), .A2(n_1270), .B1(n_1291), .B2(n_1292), .C(n_1295), .Y(n_1290) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1294), .Y(n_1410) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1943 ( .A(n_1307), .Y(n_1943) );
HB1xp67_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1308), .Y(n_1346) );
XNOR2xp5_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1376), .Y(n_1310) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_1319), .A2(n_1349), .B1(n_1350), .B2(n_1351), .Y(n_1348) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
AOI31xp33_ASAP7_75t_L g1327 ( .A1(n_1328), .A2(n_1341), .A3(n_1348), .B(n_1353), .Y(n_1327) );
AOI211xp5_ASAP7_75t_L g1328 ( .A1(n_1329), .A2(n_1332), .B(n_1333), .C(n_1336), .Y(n_1328) );
AOI222xp33_ASAP7_75t_L g1997 ( .A1(n_1329), .A2(n_1338), .B1(n_1991), .B2(n_1992), .C1(n_1998), .C2(n_1999), .Y(n_1997) );
INVx2_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
INVx2_ASAP7_75t_SL g1330 ( .A(n_1331), .Y(n_1330) );
HB1xp67_ASAP7_75t_L g1412 ( .A(n_1331), .Y(n_1412) );
BUFx2_ASAP7_75t_L g1600 ( .A(n_1331), .Y(n_1600) );
NOR3xp33_ASAP7_75t_L g1449 ( .A(n_1333), .B(n_1450), .C(n_1453), .Y(n_1449) );
CKINVDCx11_ASAP7_75t_R g1486 ( .A(n_1333), .Y(n_1486) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVxp67_ASAP7_75t_L g1493 ( .A(n_1335), .Y(n_1493) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx2_ASAP7_75t_L g1422 ( .A(n_1338), .Y(n_1422) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1338), .Y(n_1451) );
AOI322xp5_ASAP7_75t_L g1487 ( .A1(n_1338), .A2(n_1483), .A3(n_1488), .B1(n_1489), .B2(n_1490), .C1(n_1491), .C2(n_1494), .Y(n_1487) );
AOI222xp33_ASAP7_75t_L g1642 ( .A1(n_1338), .A2(n_1491), .B1(n_1643), .B2(n_1644), .C1(n_1645), .C2(n_1646), .Y(n_1642) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1340), .Y(n_1492) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1344), .B1(n_1345), .B2(n_1347), .Y(n_1341) );
AOI22xp33_ASAP7_75t_SL g1423 ( .A1(n_1342), .A2(n_1424), .B1(n_1425), .B2(n_1426), .Y(n_1423) );
AOI22xp5_ASAP7_75t_L g1454 ( .A1(n_1342), .A2(n_1425), .B1(n_1455), .B2(n_1456), .Y(n_1454) );
AOI22xp5_ASAP7_75t_L g1580 ( .A1(n_1342), .A2(n_1345), .B1(n_1581), .B2(n_1582), .Y(n_1580) );
AOI22xp33_ASAP7_75t_L g1639 ( .A1(n_1342), .A2(n_1345), .B1(n_1640), .B2(n_1641), .Y(n_1639) );
AOI22xp33_ASAP7_75t_L g1994 ( .A1(n_1342), .A2(n_1425), .B1(n_1995), .B2(n_1996), .Y(n_1994) );
AND2x4_ASAP7_75t_L g1345 ( .A(n_1343), .B(n_1346), .Y(n_1345) );
AND2x4_ASAP7_75t_L g1425 ( .A(n_1343), .B(n_1346), .Y(n_1425) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1343), .Y(n_1483) );
AOI22xp33_ASAP7_75t_SL g1427 ( .A1(n_1349), .A2(n_1388), .B1(n_1428), .B2(n_1429), .Y(n_1427) );
AOI211xp5_ASAP7_75t_L g1479 ( .A1(n_1349), .A2(n_1480), .B(n_1481), .C(n_1485), .Y(n_1479) );
AOI22xp33_ASAP7_75t_L g1583 ( .A1(n_1349), .A2(n_1351), .B1(n_1584), .B2(n_1585), .Y(n_1583) );
AOI22xp33_ASAP7_75t_L g1649 ( .A1(n_1349), .A2(n_1351), .B1(n_1632), .B2(n_1650), .Y(n_1649) );
AOI22xp33_ASAP7_75t_L g2000 ( .A1(n_1349), .A2(n_1429), .B1(n_1987), .B2(n_2001), .Y(n_2000) );
INVx4_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVx5_ASAP7_75t_L g1429 ( .A(n_1352), .Y(n_1429) );
AOI31xp33_ASAP7_75t_L g1418 ( .A1(n_1353), .A2(n_1419), .A3(n_1423), .B(n_1427), .Y(n_1418) );
AO21x1_ASAP7_75t_SL g1448 ( .A1(n_1353), .A2(n_1449), .B(n_1454), .Y(n_1448) );
CKINVDCx16_ASAP7_75t_R g1578 ( .A(n_1353), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1368), .Y(n_1354) );
AOI33xp33_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1358), .A3(n_1360), .B1(n_1361), .B2(n_1364), .B3(n_1367), .Y(n_1355) );
AOI33xp33_ASAP7_75t_L g2003 ( .A1(n_1356), .A2(n_1367), .A3(n_2004), .B1(n_2006), .B2(n_2007), .B3(n_2008), .Y(n_2003) );
BUFx3_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
NAND3xp33_ASAP7_75t_L g1408 ( .A(n_1357), .B(n_1409), .C(n_1411), .Y(n_1408) );
INVx3_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
AOI33xp33_ASAP7_75t_L g1457 ( .A1(n_1367), .A2(n_1458), .A3(n_1459), .B1(n_1460), .B2(n_1461), .B3(n_1462), .Y(n_1457) );
INVx2_ASAP7_75t_L g1531 ( .A(n_1367), .Y(n_1531) );
AOI33xp33_ASAP7_75t_L g1592 ( .A1(n_1367), .A2(n_1458), .A3(n_1593), .B1(n_1595), .B2(n_1597), .B3(n_1599), .Y(n_1592) );
XNOR2x1_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1430), .Y(n_1376) );
NAND3xp33_ASAP7_75t_L g1379 ( .A(n_1380), .B(n_1386), .C(n_1389), .Y(n_1379) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
HB1xp67_ASAP7_75t_L g1954 ( .A(n_1383), .Y(n_1954) );
NAND4xp25_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1401), .C(n_1408), .D(n_1413), .Y(n_1392) );
NAND3xp33_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1397), .C(n_1398), .Y(n_1393) );
INVx3_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
NAND3xp33_ASAP7_75t_L g1659 ( .A(n_1398), .B(n_1660), .C(n_1661), .Y(n_1659) );
INVx3_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
INVx2_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1422), .Y(n_1589) );
INVx5_ASAP7_75t_SL g1484 ( .A(n_1425), .Y(n_1484) );
AND4x1_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1448), .C(n_1457), .D(n_1463), .Y(n_1431) );
NAND4xp25_ASAP7_75t_L g1471 ( .A(n_1432), .B(n_1448), .C(n_1457), .D(n_1463), .Y(n_1471) );
OAI31xp33_ASAP7_75t_L g1432 ( .A1(n_1433), .A2(n_1440), .A3(n_1443), .B(n_1447), .Y(n_1432) );
NAND3xp33_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1436), .C(n_1439), .Y(n_1433) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1445), .Y(n_1502) );
OAI31xp33_ASAP7_75t_SL g1495 ( .A1(n_1447), .A2(n_1496), .A3(n_1497), .B(n_1498), .Y(n_1495) );
INVx1_ASAP7_75t_SL g1623 ( .A(n_1447), .Y(n_1623) );
NAND3xp33_ASAP7_75t_L g1652 ( .A(n_1458), .B(n_1653), .C(n_1655), .Y(n_1652) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
XNOR2x1_ASAP7_75t_L g1474 ( .A(n_1475), .B(n_1574), .Y(n_1474) );
XNOR2x1_ASAP7_75t_L g1475 ( .A(n_1476), .B(n_1534), .Y(n_1475) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1477), .Y(n_1532) );
OAI211xp5_ASAP7_75t_L g1477 ( .A1(n_1478), .A2(n_1479), .B(n_1495), .C(n_1505), .Y(n_1477) );
NAND4xp25_ASAP7_75t_SL g1579 ( .A(n_1486), .B(n_1580), .C(n_1583), .D(n_1586), .Y(n_1579) );
NAND4xp25_ASAP7_75t_SL g1638 ( .A(n_1486), .B(n_1639), .C(n_1642), .D(n_1649), .Y(n_1638) );
NAND4xp25_ASAP7_75t_SL g1993 ( .A(n_1486), .B(n_1994), .C(n_1997), .D(n_2000), .Y(n_1993) );
AND2x4_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1493), .Y(n_1491) );
AND2x4_ASAP7_75t_L g1999 ( .A(n_1492), .B(n_1493), .Y(n_1999) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
NOR2xp33_ASAP7_75t_L g1505 ( .A(n_1506), .B(n_1523), .Y(n_1505) );
OAI22xp5_ASAP7_75t_L g1507 ( .A1(n_1508), .A2(n_1509), .B1(n_1510), .B2(n_1511), .Y(n_1507) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
NAND4xp25_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1560), .C(n_1571), .D(n_1573), .Y(n_1535) );
OAI221xp5_ASAP7_75t_L g1537 ( .A1(n_1538), .A2(n_1542), .B1(n_1545), .B2(n_1548), .C(n_1551), .Y(n_1537) );
INVx2_ASAP7_75t_L g1598 ( .A(n_1540), .Y(n_1598) );
INVx2_ASAP7_75t_SL g1654 ( .A(n_1540), .Y(n_1654) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
OA22x2_ASAP7_75t_L g1574 ( .A1(n_1575), .A2(n_1624), .B1(n_1625), .B2(n_1668), .Y(n_1574) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1575), .Y(n_1668) );
XNOR2xp5_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1577), .Y(n_1575) );
AOI211xp5_ASAP7_75t_L g1577 ( .A1(n_1578), .A2(n_1579), .B(n_1591), .C(n_1610), .Y(n_1577) );
NAND2xp5_ASAP7_75t_SL g1591 ( .A(n_1592), .B(n_1601), .Y(n_1591) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
AOI31xp33_ASAP7_75t_SL g1610 ( .A1(n_1611), .A2(n_1617), .A3(n_1620), .B(n_1623), .Y(n_1610) );
INVx2_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1615), .Y(n_1635) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1626), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1631), .Y(n_1627) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
NAND4xp25_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1656), .C(n_1659), .D(n_1662), .Y(n_1651) );
OAI221xp5_ASAP7_75t_L g1670 ( .A1(n_1671), .A2(n_1917), .B1(n_1921), .B2(n_1966), .C(n_1971), .Y(n_1670) );
AOI21xp5_ASAP7_75t_L g1671 ( .A1(n_1672), .A2(n_1839), .B(n_1890), .Y(n_1671) );
NAND5xp2_ASAP7_75t_L g1672 ( .A(n_1673), .B(n_1761), .C(n_1803), .D(n_1820), .E(n_1835), .Y(n_1672) );
AOI211xp5_ASAP7_75t_L g1673 ( .A1(n_1674), .A2(n_1707), .B(n_1734), .C(n_1753), .Y(n_1673) );
AOI221xp5_ASAP7_75t_L g1903 ( .A1(n_1674), .A2(n_1783), .B1(n_1904), .B2(n_1905), .C(n_1906), .Y(n_1903) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
NOR2xp33_ASAP7_75t_L g1892 ( .A(n_1675), .B(n_1784), .Y(n_1892) );
OR2x2_ASAP7_75t_L g1675 ( .A(n_1676), .B(n_1700), .Y(n_1675) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1676), .Y(n_1827) );
INVx2_ASAP7_75t_L g1859 ( .A(n_1676), .Y(n_1859) );
NAND2xp5_ASAP7_75t_L g1676 ( .A(n_1677), .B(n_1697), .Y(n_1676) );
AND2x2_ASAP7_75t_L g1802 ( .A(n_1677), .B(n_1757), .Y(n_1802) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1678), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1752 ( .A(n_1678), .B(n_1700), .Y(n_1752) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1678), .Y(n_1768) );
AND2x2_ASAP7_75t_L g1775 ( .A(n_1678), .B(n_1757), .Y(n_1775) );
BUFx6f_ASAP7_75t_L g1778 ( .A(n_1678), .Y(n_1778) );
AND2x2_ASAP7_75t_L g1830 ( .A(n_1678), .B(n_1697), .Y(n_1830) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1679), .B(n_1691), .Y(n_1678) );
AND2x4_ASAP7_75t_L g1680 ( .A(n_1681), .B(n_1686), .Y(n_1680) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
OR2x2_ASAP7_75t_L g1721 ( .A(n_1682), .B(n_1687), .Y(n_1721) );
NAND2xp5_ASAP7_75t_L g1682 ( .A(n_1683), .B(n_1685), .Y(n_1682) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1685), .Y(n_1694) );
AND2x4_ASAP7_75t_L g1688 ( .A(n_1686), .B(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
OR2x2_ASAP7_75t_L g1724 ( .A(n_1687), .B(n_1690), .Y(n_1724) );
HB1xp67_ASAP7_75t_L g2025 ( .A(n_1689), .Y(n_2025) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1692), .Y(n_1703) );
BUFx3_ASAP7_75t_L g1791 ( .A(n_1692), .Y(n_1791) );
AND2x4_ASAP7_75t_L g1692 ( .A(n_1693), .B(n_1695), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_1693), .B(n_1695), .Y(n_1712) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
AND2x4_ASAP7_75t_L g1696 ( .A(n_1694), .B(n_1695), .Y(n_1696) );
INVx2_ASAP7_75t_L g1705 ( .A(n_1696), .Y(n_1705) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1697), .Y(n_1757) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1697), .Y(n_1765) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1697), .Y(n_1781) );
AND2x2_ASAP7_75t_L g1846 ( .A(n_1697), .B(n_1772), .Y(n_1846) );
NAND2xp5_ASAP7_75t_L g1866 ( .A(n_1697), .B(n_1715), .Y(n_1866) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1698), .B(n_1699), .Y(n_1697) );
AND2x2_ASAP7_75t_L g1767 ( .A(n_1700), .B(n_1768), .Y(n_1767) );
CKINVDCx6p67_ASAP7_75t_R g1772 ( .A(n_1700), .Y(n_1772) );
OR2x2_ASAP7_75t_L g1818 ( .A(n_1700), .B(n_1768), .Y(n_1818) );
NAND2xp5_ASAP7_75t_L g1834 ( .A(n_1700), .B(n_1814), .Y(n_1834) );
OAI322xp33_ASAP7_75t_L g1847 ( .A1(n_1700), .A2(n_1848), .A3(n_1849), .B1(n_1850), .B2(n_1851), .C1(n_1853), .C2(n_1854), .Y(n_1847) );
AND2x2_ASAP7_75t_L g1876 ( .A(n_1700), .B(n_1802), .Y(n_1876) );
NAND2xp5_ASAP7_75t_L g1884 ( .A(n_1700), .B(n_1885), .Y(n_1884) );
OR2x6_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1702), .Y(n_1700) );
OR2x2_ASAP7_75t_L g1754 ( .A(n_1701), .B(n_1702), .Y(n_1754) );
OAI22xp5_ASAP7_75t_SL g1702 ( .A1(n_1703), .A2(n_1704), .B1(n_1705), .B2(n_1706), .Y(n_1702) );
INVx2_ASAP7_75t_L g1717 ( .A(n_1705), .Y(n_1717) );
INVx1_ASAP7_75t_L g1792 ( .A(n_1705), .Y(n_1792) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1708), .B(n_1713), .Y(n_1707) );
AND2x2_ASAP7_75t_L g1738 ( .A(n_1708), .B(n_1739), .Y(n_1738) );
AND2x2_ASAP7_75t_L g1749 ( .A(n_1708), .B(n_1750), .Y(n_1749) );
AND2x2_ASAP7_75t_L g1758 ( .A(n_1708), .B(n_1759), .Y(n_1758) );
AND2x2_ASAP7_75t_L g1829 ( .A(n_1708), .B(n_1716), .Y(n_1829) );
OR2x2_ASAP7_75t_L g1873 ( .A(n_1708), .B(n_1874), .Y(n_1873) );
AND2x2_ASAP7_75t_L g1904 ( .A(n_1708), .B(n_1762), .Y(n_1904) );
AND2x2_ASAP7_75t_L g1913 ( .A(n_1708), .B(n_1726), .Y(n_1913) );
CKINVDCx5p33_ASAP7_75t_R g1708 ( .A(n_1709), .Y(n_1708) );
AND2x2_ASAP7_75t_L g1742 ( .A(n_1709), .B(n_1743), .Y(n_1742) );
AND2x2_ASAP7_75t_L g1773 ( .A(n_1709), .B(n_1726), .Y(n_1773) );
AND2x2_ASAP7_75t_L g1780 ( .A(n_1709), .B(n_1715), .Y(n_1780) );
OR2x2_ASAP7_75t_L g1805 ( .A(n_1709), .B(n_1806), .Y(n_1805) );
AND2x2_ASAP7_75t_L g1809 ( .A(n_1709), .B(n_1739), .Y(n_1809) );
AND2x2_ASAP7_75t_L g1819 ( .A(n_1709), .B(n_1750), .Y(n_1819) );
NAND2xp5_ASAP7_75t_L g1824 ( .A(n_1709), .B(n_1731), .Y(n_1824) );
AND2x2_ASAP7_75t_L g1844 ( .A(n_1709), .B(n_1759), .Y(n_1844) );
HB1xp67_ASAP7_75t_L g1849 ( .A(n_1709), .Y(n_1849) );
AND2x2_ASAP7_75t_L g1852 ( .A(n_1709), .B(n_1807), .Y(n_1852) );
NOR2xp33_ASAP7_75t_L g1878 ( .A(n_1709), .B(n_1879), .Y(n_1878) );
NOR2xp33_ASAP7_75t_L g1902 ( .A(n_1709), .B(n_1807), .Y(n_1902) );
AND2x4_ASAP7_75t_SL g1709 ( .A(n_1710), .B(n_1711), .Y(n_1709) );
INVxp67_ASAP7_75t_SL g1853 ( .A(n_1713), .Y(n_1853) );
NOR2xp33_ASAP7_75t_L g1713 ( .A(n_1714), .B(n_1725), .Y(n_1713) );
NOR2x1p5_ASAP7_75t_L g1762 ( .A(n_1714), .B(n_1763), .Y(n_1762) );
AND2x2_ASAP7_75t_L g1801 ( .A(n_1714), .B(n_1802), .Y(n_1801) );
HB1xp67_ASAP7_75t_L g1843 ( .A(n_1714), .Y(n_1843) );
NAND2xp5_ASAP7_75t_L g1874 ( .A(n_1714), .B(n_1739), .Y(n_1874) );
INVxp67_ASAP7_75t_L g1885 ( .A(n_1714), .Y(n_1885) );
INVx2_ASAP7_75t_SL g1714 ( .A(n_1715), .Y(n_1714) );
BUFx2_ASAP7_75t_L g1746 ( .A(n_1715), .Y(n_1746) );
BUFx3_ASAP7_75t_L g1748 ( .A(n_1715), .Y(n_1748) );
NOR2xp33_ASAP7_75t_L g1756 ( .A(n_1715), .B(n_1757), .Y(n_1756) );
AND2x2_ASAP7_75t_L g1868 ( .A(n_1715), .B(n_1765), .Y(n_1868) );
INVx2_ASAP7_75t_SL g1715 ( .A(n_1716), .Y(n_1715) );
OAI22xp33_ASAP7_75t_L g1718 ( .A1(n_1719), .A2(n_1720), .B1(n_1722), .B2(n_1723), .Y(n_1718) );
BUFx3_ASAP7_75t_L g1795 ( .A(n_1720), .Y(n_1795) );
BUFx6f_ASAP7_75t_L g1720 ( .A(n_1721), .Y(n_1720) );
HB1xp67_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
INVx1_ASAP7_75t_L g1798 ( .A(n_1724), .Y(n_1798) );
NOR2xp33_ASAP7_75t_L g1799 ( .A(n_1725), .B(n_1800), .Y(n_1799) );
OR2x2_ASAP7_75t_L g1832 ( .A(n_1725), .B(n_1746), .Y(n_1832) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1726), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1845 ( .A(n_1726), .B(n_1829), .Y(n_1845) );
NAND3xp33_ASAP7_75t_L g1867 ( .A(n_1726), .B(n_1868), .C(n_1869), .Y(n_1867) );
AND2x2_ASAP7_75t_L g1910 ( .A(n_1726), .B(n_1780), .Y(n_1910) );
AND2x2_ASAP7_75t_L g1726 ( .A(n_1727), .B(n_1730), .Y(n_1726) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1727), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1727), .B(n_1731), .Y(n_1750) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1728), .B(n_1729), .Y(n_1727) );
INVxp67_ASAP7_75t_SL g1730 ( .A(n_1731), .Y(n_1730) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1731), .B(n_1740), .Y(n_1739) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1731), .Y(n_1743) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1731), .Y(n_1760) );
AND2x2_ASAP7_75t_L g1731 ( .A(n_1732), .B(n_1733), .Y(n_1731) );
O2A1O1Ixp33_ASAP7_75t_L g1734 ( .A1(n_1735), .A2(n_1744), .B(n_1747), .C(n_1751), .Y(n_1734) );
INVxp67_ASAP7_75t_SL g1735 ( .A(n_1736), .Y(n_1735) );
NAND2xp5_ASAP7_75t_L g1736 ( .A(n_1737), .B(n_1741), .Y(n_1736) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
AOI221xp5_ASAP7_75t_L g1875 ( .A1(n_1738), .A2(n_1771), .B1(n_1876), .B2(n_1877), .C(n_1880), .Y(n_1875) );
INVx2_ASAP7_75t_L g1763 ( .A(n_1739), .Y(n_1763) );
AND2x2_ASAP7_75t_L g1779 ( .A(n_1739), .B(n_1780), .Y(n_1779) );
AND2x2_ASAP7_75t_L g1828 ( .A(n_1739), .B(n_1829), .Y(n_1828) );
AND2x2_ASAP7_75t_L g1759 ( .A(n_1740), .B(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1740), .Y(n_1807) );
NOR2xp33_ASAP7_75t_L g1810 ( .A(n_1741), .B(n_1800), .Y(n_1810) );
O2A1O1Ixp33_ASAP7_75t_SL g1906 ( .A1(n_1741), .A2(n_1754), .B(n_1907), .C(n_1909), .Y(n_1906) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1743), .Y(n_1879) );
A2O1A1Ixp33_ASAP7_75t_L g1916 ( .A1(n_1744), .A2(n_1759), .B(n_1785), .C(n_1844), .Y(n_1916) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
AND2x2_ASAP7_75t_L g1877 ( .A(n_1745), .B(n_1878), .Y(n_1877) );
INVx2_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
AND2x2_ASAP7_75t_L g1888 ( .A(n_1746), .B(n_1750), .Y(n_1888) );
AND2x2_ASAP7_75t_L g1908 ( .A(n_1746), .B(n_1864), .Y(n_1908) );
INVx1_ASAP7_75t_L g1893 ( .A(n_1747), .Y(n_1893) );
NAND2xp5_ASAP7_75t_L g1747 ( .A(n_1748), .B(n_1749), .Y(n_1747) );
INVx1_ASAP7_75t_L g1784 ( .A(n_1748), .Y(n_1784) );
AND2x2_ASAP7_75t_L g1838 ( .A(n_1748), .B(n_1758), .Y(n_1838) );
NAND2xp5_ASAP7_75t_L g1848 ( .A(n_1748), .B(n_1802), .Y(n_1848) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1750), .Y(n_1861) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
NAND2xp5_ASAP7_75t_L g1786 ( .A(n_1752), .B(n_1781), .Y(n_1786) );
AOI22xp5_ASAP7_75t_L g1870 ( .A1(n_1752), .A2(n_1778), .B1(n_1871), .B2(n_1872), .Y(n_1870) );
AOI221xp5_ASAP7_75t_L g1912 ( .A1(n_1752), .A2(n_1865), .B1(n_1876), .B2(n_1913), .C(n_1914), .Y(n_1912) );
NOR2xp33_ASAP7_75t_L g1753 ( .A(n_1754), .B(n_1755), .Y(n_1753) );
AOI211xp5_ASAP7_75t_L g1803 ( .A1(n_1754), .A2(n_1804), .B(n_1810), .C(n_1811), .Y(n_1803) );
A2O1A1Ixp33_ASAP7_75t_L g1911 ( .A1(n_1754), .A2(n_1809), .B(n_1836), .C(n_1859), .Y(n_1911) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1755), .Y(n_1871) );
NAND2xp5_ASAP7_75t_L g1755 ( .A(n_1756), .B(n_1758), .Y(n_1755) );
OAI21xp33_ASAP7_75t_L g1816 ( .A1(n_1756), .A2(n_1817), .B(n_1819), .Y(n_1816) );
AND2x2_ASAP7_75t_L g1855 ( .A(n_1757), .B(n_1772), .Y(n_1855) );
NOR2xp33_ASAP7_75t_L g1822 ( .A(n_1758), .B(n_1823), .Y(n_1822) );
AOI221xp5_ASAP7_75t_L g1782 ( .A1(n_1759), .A2(n_1771), .B1(n_1783), .B2(n_1785), .C(n_1787), .Y(n_1782) );
AND2x2_ASAP7_75t_L g1783 ( .A(n_1759), .B(n_1784), .Y(n_1783) );
INVx1_ASAP7_75t_L g1887 ( .A(n_1759), .Y(n_1887) );
AOI211xp5_ASAP7_75t_L g1761 ( .A1(n_1762), .A2(n_1764), .B(n_1776), .C(n_1799), .Y(n_1761) );
A2O1A1Ixp33_ASAP7_75t_L g1895 ( .A1(n_1762), .A2(n_1817), .B(n_1845), .C(n_1896), .Y(n_1895) );
OAI211xp5_ASAP7_75t_L g1764 ( .A1(n_1765), .A2(n_1766), .B(n_1769), .C(n_1774), .Y(n_1764) );
NAND2xp67_ASAP7_75t_L g1909 ( .A(n_1765), .B(n_1910), .Y(n_1909) );
INVx1_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1768), .B(n_1772), .Y(n_1771) );
INVx1_ASAP7_75t_L g1864 ( .A(n_1768), .Y(n_1864) );
A2O1A1Ixp33_ASAP7_75t_L g1776 ( .A1(n_1769), .A2(n_1777), .B(n_1781), .C(n_1782), .Y(n_1776) );
NAND2xp5_ASAP7_75t_L g1769 ( .A(n_1770), .B(n_1773), .Y(n_1769) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1771), .Y(n_1770) );
NOR2xp33_ASAP7_75t_L g1836 ( .A(n_1772), .B(n_1837), .Y(n_1836) );
NAND2xp5_ASAP7_75t_SL g1850 ( .A(n_1772), .B(n_1802), .Y(n_1850) );
AND2x2_ASAP7_75t_L g1899 ( .A(n_1772), .B(n_1775), .Y(n_1899) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1773), .Y(n_1881) );
INVx1_ASAP7_75t_L g1774 ( .A(n_1775), .Y(n_1774) );
AOI21xp5_ASAP7_75t_L g1856 ( .A1(n_1775), .A2(n_1845), .B(n_1857), .Y(n_1856) );
NAND2xp5_ASAP7_75t_L g1777 ( .A(n_1778), .B(n_1779), .Y(n_1777) );
OAI22xp33_ASAP7_75t_L g1804 ( .A1(n_1778), .A2(n_1800), .B1(n_1805), .B2(n_1808), .Y(n_1804) );
CKINVDCx14_ASAP7_75t_R g1869 ( .A(n_1778), .Y(n_1869) );
INVx1_ASAP7_75t_L g1815 ( .A(n_1779), .Y(n_1815) );
INVx3_ASAP7_75t_L g1814 ( .A(n_1781), .Y(n_1814) );
NAND2xp5_ASAP7_75t_L g1826 ( .A(n_1784), .B(n_1827), .Y(n_1826) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
INVx3_ASAP7_75t_L g1889 ( .A(n_1787), .Y(n_1889) );
INVx2_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
INVx1_ASAP7_75t_L g1788 ( .A(n_1789), .Y(n_1788) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
OAI22xp33_ASAP7_75t_L g1793 ( .A1(n_1794), .A2(n_1795), .B1(n_1796), .B2(n_1797), .Y(n_1793) );
HB1xp67_ASAP7_75t_L g1920 ( .A(n_1797), .Y(n_1920) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
INVx1_ASAP7_75t_L g1800 ( .A(n_1801), .Y(n_1800) );
NAND3xp33_ASAP7_75t_L g1915 ( .A(n_1802), .B(n_1823), .C(n_1883), .Y(n_1915) );
NOR2xp33_ASAP7_75t_L g1865 ( .A(n_1805), .B(n_1866), .Y(n_1865) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1807), .Y(n_1806) );
INVx1_ASAP7_75t_L g1808 ( .A(n_1809), .Y(n_1808) );
OAI21xp33_ASAP7_75t_L g1811 ( .A1(n_1812), .A2(n_1815), .B(n_1816), .Y(n_1811) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
INVx1_ASAP7_75t_L g1896 ( .A(n_1813), .Y(n_1896) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1814), .Y(n_1813) );
INVx1_ASAP7_75t_L g1817 ( .A(n_1818), .Y(n_1817) );
AOI221xp5_ASAP7_75t_L g1891 ( .A1(n_1819), .A2(n_1830), .B1(n_1892), .B2(n_1893), .C(n_1894), .Y(n_1891) );
AOI222xp33_ASAP7_75t_L g1820 ( .A1(n_1821), .A2(n_1825), .B1(n_1828), .B2(n_1830), .C1(n_1831), .C2(n_1833), .Y(n_1820) );
INVxp67_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
INVx1_ASAP7_75t_L g1823 ( .A(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g1825 ( .A(n_1826), .Y(n_1825) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1829), .Y(n_1862) );
OAI211xp5_ASAP7_75t_L g1897 ( .A1(n_1829), .A2(n_1898), .B(n_1899), .C(n_1900), .Y(n_1897) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1832), .Y(n_1831) );
AOI321xp33_ASAP7_75t_L g1882 ( .A1(n_1833), .A2(n_1849), .A3(n_1883), .B1(n_1886), .B2(n_1888), .C(n_1889), .Y(n_1882) );
INVx1_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
INVxp67_ASAP7_75t_SL g1835 ( .A(n_1836), .Y(n_1835) );
INVx1_ASAP7_75t_L g1837 ( .A(n_1838), .Y(n_1837) );
NAND5xp2_ASAP7_75t_L g1839 ( .A(n_1840), .B(n_1856), .C(n_1870), .D(n_1875), .E(n_1882), .Y(n_1839) );
O2A1O1Ixp33_ASAP7_75t_L g1840 ( .A1(n_1841), .A2(n_1845), .B(n_1846), .C(n_1847), .Y(n_1840) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
NAND2xp5_ASAP7_75t_L g1842 ( .A(n_1843), .B(n_1844), .Y(n_1842) );
INVx1_ASAP7_75t_L g1905 ( .A(n_1850), .Y(n_1905) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1852), .Y(n_1851) );
NOR2xp33_ASAP7_75t_L g1880 ( .A(n_1854), .B(n_1881), .Y(n_1880) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1855), .Y(n_1854) );
OAI211xp5_ASAP7_75t_SL g1857 ( .A1(n_1858), .A2(n_1860), .B(n_1863), .C(n_1867), .Y(n_1857) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
OR2x2_ASAP7_75t_L g1860 ( .A(n_1861), .B(n_1862), .Y(n_1860) );
NAND2xp5_ASAP7_75t_L g1886 ( .A(n_1861), .B(n_1887), .Y(n_1886) );
NAND2xp5_ASAP7_75t_L g1863 ( .A(n_1864), .B(n_1865), .Y(n_1863) );
INVx2_ASAP7_75t_L g1872 ( .A(n_1873), .Y(n_1872) );
INVx1_ASAP7_75t_L g1898 ( .A(n_1874), .Y(n_1898) );
INVx1_ASAP7_75t_L g1883 ( .A(n_1884), .Y(n_1883) );
NAND5xp2_ASAP7_75t_L g1890 ( .A(n_1891), .B(n_1903), .C(n_1911), .D(n_1912), .E(n_1916), .Y(n_1890) );
NAND2xp5_ASAP7_75t_SL g1894 ( .A(n_1895), .B(n_1897), .Y(n_1894) );
INVx1_ASAP7_75t_L g1900 ( .A(n_1901), .Y(n_1900) );
HB1xp67_ASAP7_75t_L g1901 ( .A(n_1902), .Y(n_1901) );
INVx1_ASAP7_75t_L g1907 ( .A(n_1908), .Y(n_1907) );
INVxp67_ASAP7_75t_SL g1914 ( .A(n_1915), .Y(n_1914) );
CKINVDCx5p33_ASAP7_75t_R g1917 ( .A(n_1918), .Y(n_1917) );
INVx1_ASAP7_75t_SL g1918 ( .A(n_1919), .Y(n_1918) );
BUFx2_ASAP7_75t_SL g1919 ( .A(n_1920), .Y(n_1919) );
INVx1_ASAP7_75t_L g1965 ( .A(n_1922), .Y(n_1965) );
INVx1_ASAP7_75t_L g1922 ( .A(n_1923), .Y(n_1922) );
NAND2xp5_ASAP7_75t_L g1923 ( .A(n_1924), .B(n_1950), .Y(n_1923) );
NOR3xp33_ASAP7_75t_L g1924 ( .A(n_1925), .B(n_1932), .C(n_1933), .Y(n_1924) );
NAND2xp5_ASAP7_75t_L g1925 ( .A(n_1926), .B(n_1929), .Y(n_1925) );
OAI22xp33_ASAP7_75t_L g1934 ( .A1(n_1935), .A2(n_1936), .B1(n_1937), .B2(n_1938), .Y(n_1934) );
INVx1_ASAP7_75t_L g1942 ( .A(n_1943), .Y(n_1942) );
NAND3xp33_ASAP7_75t_L g1951 ( .A(n_1952), .B(n_1959), .C(n_1962), .Y(n_1951) );
BUFx2_ASAP7_75t_L g1956 ( .A(n_1957), .Y(n_1956) );
CKINVDCx14_ASAP7_75t_R g1966 ( .A(n_1967), .Y(n_1966) );
INVx2_ASAP7_75t_L g1967 ( .A(n_1968), .Y(n_1967) );
CKINVDCx5p33_ASAP7_75t_R g1968 ( .A(n_1969), .Y(n_1968) );
OAI21xp5_ASAP7_75t_L g2024 ( .A1(n_1970), .A2(n_2025), .B(n_2026), .Y(n_2024) );
INVx1_ASAP7_75t_L g1972 ( .A(n_1973), .Y(n_1972) );
INVx1_ASAP7_75t_L g1973 ( .A(n_1974), .Y(n_1973) );
INVx1_ASAP7_75t_L g1974 ( .A(n_1975), .Y(n_1974) );
INVx1_ASAP7_75t_L g1975 ( .A(n_1976), .Y(n_1975) );
INVx1_ASAP7_75t_L g1977 ( .A(n_1978), .Y(n_1977) );
HB1xp67_ASAP7_75t_L g1978 ( .A(n_1979), .Y(n_1978) );
INVx1_ASAP7_75t_L g1979 ( .A(n_1980), .Y(n_1979) );
INVx1_ASAP7_75t_L g2022 ( .A(n_1981), .Y(n_2022) );
NAND2xp5_ASAP7_75t_L g2002 ( .A(n_2003), .B(n_2009), .Y(n_2002) );
INVx1_ASAP7_75t_L g2012 ( .A(n_2013), .Y(n_2012) );
INVx2_ASAP7_75t_L g2015 ( .A(n_2016), .Y(n_2015) );
INVx1_ASAP7_75t_L g2017 ( .A(n_2018), .Y(n_2017) );
HB1xp67_ASAP7_75t_L g2023 ( .A(n_2024), .Y(n_2023) );
endmodule