module real_jpeg_10306_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_345, n_6, n_346, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_345;
input n_6;
input n_346;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_1),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_1),
.A2(n_65),
.B1(n_68),
.B2(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_90),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_90),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_2),
.A2(n_15),
.B(n_32),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_3),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_3),
.A2(n_22),
.B1(n_65),
.B2(n_68),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_3),
.A2(n_22),
.B1(n_47),
.B2(n_48),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_4),
.A2(n_23),
.B1(n_25),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_4),
.A2(n_55),
.B1(n_65),
.B2(n_68),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_5),
.A2(n_57),
.B1(n_65),
.B2(n_68),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_8),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_8),
.A2(n_34),
.B1(n_65),
.B2(n_68),
.Y(n_232)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_11),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_11),
.A2(n_65),
.B1(n_68),
.B2(n_102),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_102),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_102),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_12),
.A2(n_65),
.B1(n_68),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_12),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_107),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_107),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_107),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_13),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

A2O1A1O1Ixp25_ASAP7_75t_L g86 ( 
.A1(n_15),
.A2(n_48),
.B(n_60),
.C(n_87),
.D(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_15),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_15),
.B(n_46),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_15),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_15),
.A2(n_108),
.B(n_111),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_15),
.A2(n_31),
.B(n_42),
.C(n_143),
.D(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_15),
.B(n_31),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_15),
.B(n_35),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_15),
.A2(n_23),
.B1(n_25),
.B2(n_124),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_16),
.A2(n_65),
.B1(n_68),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_16),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_155),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_155),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_16),
.A2(n_23),
.B1(n_25),
.B2(n_155),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_338),
.B(n_341),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_76),
.B(n_337),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_20),
.B(n_36),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_20),
.B(n_339),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_20),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_21),
.A2(n_26),
.B1(n_35),
.B2(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_23),
.A2(n_28),
.B(n_124),
.C(n_186),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_26),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_26),
.B(n_206),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_26),
.A2(n_33),
.B(n_35),
.Y(n_340)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_27),
.A2(n_30),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_27),
.A2(n_30),
.B1(n_214),
.B2(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_27),
.A2(n_205),
.B(n_243),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_27),
.A2(n_30),
.B1(n_54),
.B2(n_287),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_30),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_30),
.A2(n_215),
.B(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_35),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_71),
.C(n_73),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_37),
.A2(n_38),
.B1(n_332),
.B2(n_334),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_52),
.C(n_58),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_39),
.A2(n_40),
.B1(n_58),
.B2(n_312),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_41),
.A2(n_50),
.B1(n_164),
.B2(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_41),
.A2(n_200),
.B(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_46),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_42),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_42),
.A2(n_46),
.B1(n_240),
.B2(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_42),
.A2(n_46),
.B1(n_259),
.B2(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_43),
.B(n_48),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_45),
.A2(n_47),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_61),
.B(n_63),
.C(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_50),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_50),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_50),
.A2(n_165),
.B(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_52),
.A2(n_53),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_58),
.A2(n_310),
.B1(n_312),
.B2(n_313),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_58),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_69),
.B(n_70),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_59),
.A2(n_69),
.B1(n_101),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_59),
.A2(n_141),
.B(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_59),
.A2(n_69),
.B1(n_197),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_59),
.A2(n_69),
.B1(n_225),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_59),
.A2(n_69),
.B1(n_234),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_60),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_60),
.A2(n_64),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_68),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_68),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_65),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_68),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_68),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_69),
.A2(n_103),
.B(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_70),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_71),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_330),
.B(n_336),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_303),
.A3(n_323),
.B1(n_328),
.B2(n_329),
.C(n_345),
.Y(n_77)
);

AOI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_251),
.A3(n_291),
.B1(n_297),
.B2(n_302),
.C(n_346),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_208),
.C(n_247),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_179),
.B(n_207),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_158),
.B(n_178),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_135),
.B(n_157),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_113),
.B(n_134),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_95),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_85),
.B(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_86),
.A2(n_91),
.B1(n_92),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_88),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_100),
.C(n_105),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_111),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_106),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_108),
.A2(n_126),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_108),
.A2(n_126),
.B1(n_190),
.B2(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_108),
.A2(n_126),
.B1(n_223),
.B2(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_108),
.A2(n_126),
.B(n_232),
.Y(n_264)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_109),
.A2(n_110),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_112),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_109),
.A2(n_110),
.B1(n_154),
.B2(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_121),
.B(n_133),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_119),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_128),
.B(n_132),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_126),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_127),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_136),
.B(n_137),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_148),
.B2(n_156),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_147),
.C(n_156),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_144),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_148),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_152),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_160),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_172),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_174),
.C(n_176),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_167),
.B2(n_171),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_168),
.C(n_169),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_174),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_181),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_194),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_183),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_183),
.B(n_193),
.C(n_194),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_188),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_191),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_196),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_209),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_227),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_210),
.B(n_227),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_221),
.C(n_226),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_220),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_219),
.C(n_220),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_226),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_224),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_245),
.B2(n_246),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_230),
.B(n_235),
.C(n_246),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_233),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_241),
.C(n_244),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_238),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_249),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_269),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_252),
.B(n_269),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_262),
.C(n_268),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_253),
.A2(n_254),
.B1(n_262),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_258),
.C(n_260),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_262),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_264),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_263),
.A2(n_282),
.B(n_286),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_265),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_265),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_266),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_289),
.B2(n_290),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_280),
.B2(n_281),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_281),
.C(n_290),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_277),
.B(n_279),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_277),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_278),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_279),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_279),
.A2(n_305),
.B1(n_314),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_288),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_284),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_298),
.B(n_301),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_293),
.B(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_316),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_316),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_314),
.C(n_315),
.Y(n_304)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_305),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_307),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_312),
.C(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_318),
.C(n_322),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_310),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_335),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_332),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_340),
.B(n_343),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);


endmodule