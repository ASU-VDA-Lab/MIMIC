module fake_jpeg_21962_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_37),
.CON(n_47),
.SN(n_47)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_42),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_22),
.C(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_30),
.Y(n_75)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_18),
.B1(n_24),
.B2(n_29),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_48),
.A2(n_49),
.B1(n_54),
.B2(n_66),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_18),
.B1(n_24),
.B2(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_52),
.Y(n_86)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_59),
.Y(n_99)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

CKINVDCx6p67_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_67),
.Y(n_101)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_73),
.Y(n_80)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_36),
.A2(n_27),
.B1(n_23),
.B2(n_34),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_25),
.B1(n_30),
.B2(n_20),
.Y(n_106)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_19),
.Y(n_73)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_32),
.B1(n_17),
.B2(n_31),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_44),
.B1(n_28),
.B2(n_22),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_82),
.A2(n_85),
.B1(n_96),
.B2(n_105),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_44),
.B1(n_37),
.B2(n_43),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_100),
.B1(n_107),
.B2(n_53),
.Y(n_112)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_44),
.B1(n_28),
.B2(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_97),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_43),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_32),
.C(n_33),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_45),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_78),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_28),
.B1(n_21),
.B2(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_45),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_74),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_50),
.A2(n_41),
.B1(n_27),
.B2(n_25),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_27),
.Y(n_103)
);

NOR2xp67_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_64),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_50),
.A2(n_25),
.B1(n_20),
.B2(n_30),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_108),
.B1(n_33),
.B2(n_56),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_61),
.A2(n_17),
.B1(n_16),
.B2(n_20),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_68),
.B(n_59),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_124),
.B(n_135),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_66),
.B1(n_53),
.B2(n_55),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_110),
.A2(n_134),
.B1(n_89),
.B2(n_104),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_132),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_112),
.A2(n_116),
.B1(n_96),
.B2(n_90),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_72),
.C(n_54),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_100),
.C(n_88),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_117),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_55),
.B1(n_52),
.B2(n_67),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_72),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_74),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_122),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_94),
.B1(n_90),
.B2(n_107),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_95),
.Y(n_121)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_130),
.B1(n_133),
.B2(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_102),
.B(n_10),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_70),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_9),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_1),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_82),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_82),
.A2(n_63),
.B1(n_9),
.B2(n_3),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_8),
.A3(n_14),
.B1(n_3),
.B2(n_5),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_1),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

BUFx6f_ASAP7_75t_SL g138 ( 
.A(n_123),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_SL g141 ( 
.A(n_124),
.B(n_96),
.C(n_103),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_147),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_103),
.B1(n_88),
.B2(n_106),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_155),
.B1(n_110),
.B2(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_146),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_161),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_160),
.B1(n_128),
.B2(n_122),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_96),
.B(n_86),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_157),
.B(n_158),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_131),
.B1(n_113),
.B2(n_123),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_114),
.A2(n_101),
.B(n_83),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_104),
.B(n_83),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_166),
.Y(n_181)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_167),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_169),
.B1(n_174),
.B2(n_178),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_121),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_159),
.C(n_156),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_129),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_180),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_112),
.B1(n_135),
.B2(n_129),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_148),
.Y(n_185)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_148),
.A3(n_141),
.B1(n_159),
.B2(n_142),
.C1(n_156),
.C2(n_157),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_173),
.B(n_172),
.C(n_180),
.D(n_162),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_113),
.B(n_136),
.C(n_125),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_133),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_185),
.A2(n_152),
.B(n_139),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_188),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_190),
.B(n_170),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_155),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_194),
.Y(n_208)
);

OAI322xp33_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_149),
.A3(n_154),
.B1(n_144),
.B2(n_143),
.C1(n_161),
.C2(n_137),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_111),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_192),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_137),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_154),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_195),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_125),
.C(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_147),
.C(n_130),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_139),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_164),
.B1(n_163),
.B2(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_197),
.B(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_169),
.B1(n_178),
.B2(n_175),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_204),
.B(n_209),
.Y(n_210)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_167),
.C(n_180),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_204),
.C(n_200),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_178),
.B1(n_175),
.B2(n_166),
.Y(n_204)
);

AOI211xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_207),
.B(n_193),
.C(n_152),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_184),
.A2(n_188),
.B1(n_192),
.B2(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_179),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_209),
.A2(n_186),
.B(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_216),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_202),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_191),
.B(n_153),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_218),
.B(n_198),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_217),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_126),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_165),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_15),
.B(n_8),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_206),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_222),
.B(n_224),
.Y(n_230)
);

NAND4xp25_ASAP7_75t_SL g221 ( 
.A(n_219),
.B(n_211),
.C(n_210),
.D(n_1),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_226),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_224),
.B(n_11),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_201),
.B1(n_3),
.B2(n_5),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_221),
.A2(n_214),
.B1(n_201),
.B2(n_7),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_10),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_12),
.Y(n_235)
);

AOI21x1_ASAP7_75t_L g233 ( 
.A1(n_230),
.A2(n_231),
.B(n_10),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_225),
.A2(n_6),
.B(n_8),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_234),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_13),
.C(n_14),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_225),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_13),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_234),
.C(n_2),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_238),
.A2(n_2),
.B(n_236),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);


endmodule