module real_aes_8407_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_L g435 ( .A1(n_0), .A2(n_7), .B1(n_436), .B2(n_708), .C1(n_713), .C2(n_714), .Y(n_435) );
INVx1_ASAP7_75t_L g104 ( .A(n_1), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_2), .A2(n_137), .B(n_142), .C(n_179), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_3), .A2(n_132), .B(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g448 ( .A(n_4), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_5), .B(n_156), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_6), .B(n_432), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_7), .Y(n_713) );
AOI21xp33_ASAP7_75t_L g465 ( .A1(n_8), .A2(n_132), .B(n_466), .Y(n_465) );
AND2x6_ASAP7_75t_L g137 ( .A(n_9), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g166 ( .A(n_10), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_11), .B(n_43), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_11), .B(n_43), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_12), .A2(n_244), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_13), .B(n_147), .Y(n_183) );
INVx1_ASAP7_75t_L g470 ( .A(n_14), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_15), .B(n_146), .Y(n_518) );
INVx1_ASAP7_75t_L g130 ( .A(n_16), .Y(n_130) );
INVx1_ASAP7_75t_L g530 ( .A(n_17), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_18), .A2(n_167), .B(n_192), .C(n_194), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_19), .B(n_156), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_20), .B(n_459), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_21), .B(n_132), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_22), .B(n_252), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_23), .A2(n_146), .B(n_148), .C(n_152), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_24), .B(n_156), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_25), .B(n_147), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_26), .A2(n_150), .B(n_194), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_27), .B(n_147), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g212 ( .A(n_28), .Y(n_212) );
INVx1_ASAP7_75t_L g226 ( .A(n_29), .Y(n_226) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_30), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_31), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_32), .B(n_147), .Y(n_449) );
INVx1_ASAP7_75t_L g249 ( .A(n_33), .Y(n_249) );
INVx1_ASAP7_75t_L g483 ( .A(n_34), .Y(n_483) );
INVx2_ASAP7_75t_L g135 ( .A(n_35), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_36), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_37), .A2(n_146), .B(n_205), .C(n_207), .Y(n_204) );
INVxp67_ASAP7_75t_L g250 ( .A(n_38), .Y(n_250) );
CKINVDCx14_ASAP7_75t_R g203 ( .A(n_39), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_40), .A2(n_142), .B(n_225), .C(n_231), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_41), .A2(n_137), .B(n_142), .C(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g114 ( .A1(n_42), .A2(n_115), .B1(n_116), .B2(n_423), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_42), .Y(n_423) );
INVx1_ASAP7_75t_L g482 ( .A(n_44), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_45), .A2(n_164), .B(n_165), .C(n_168), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_46), .B(n_147), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_47), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_48), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_49), .A2(n_100), .B1(n_108), .B2(n_719), .Y(n_99) );
INVx1_ASAP7_75t_L g140 ( .A(n_50), .Y(n_140) );
CKINVDCx16_ASAP7_75t_R g484 ( .A(n_51), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_52), .B(n_132), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_53), .A2(n_142), .B1(n_152), .B2(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_54), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g445 ( .A(n_55), .Y(n_445) );
CKINVDCx14_ASAP7_75t_R g162 ( .A(n_56), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_57), .A2(n_164), .B(n_207), .C(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_58), .Y(n_511) );
INVx1_ASAP7_75t_L g467 ( .A(n_59), .Y(n_467) );
INVx1_ASAP7_75t_L g138 ( .A(n_60), .Y(n_138) );
INVx1_ASAP7_75t_L g129 ( .A(n_61), .Y(n_129) );
INVx1_ASAP7_75t_SL g206 ( .A(n_62), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_63), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_64), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g215 ( .A(n_65), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_SL g458 ( .A1(n_66), .A2(n_207), .B(n_459), .C(n_460), .Y(n_458) );
INVxp67_ASAP7_75t_L g461 ( .A(n_67), .Y(n_461) );
INVx1_ASAP7_75t_L g107 ( .A(n_68), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_69), .A2(n_132), .B(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_70), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_71), .A2(n_132), .B(n_189), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_72), .Y(n_486) );
INVx1_ASAP7_75t_L g505 ( .A(n_73), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_74), .A2(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g190 ( .A(n_75), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_76), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_77), .A2(n_137), .B(n_142), .C(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_78), .A2(n_132), .B(n_139), .Y(n_131) );
INVx1_ASAP7_75t_L g193 ( .A(n_79), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_80), .B(n_227), .Y(n_499) );
INVx2_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
INVx1_ASAP7_75t_L g180 ( .A(n_82), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_83), .B(n_459), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_84), .A2(n_137), .B(n_142), .C(n_447), .Y(n_446) );
NAND3xp33_ASAP7_75t_SL g103 ( .A(n_85), .B(n_104), .C(n_105), .Y(n_103) );
OR2x2_ASAP7_75t_L g427 ( .A(n_85), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g706 ( .A(n_85), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_85), .B(n_429), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_86), .A2(n_142), .B(n_214), .C(n_217), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_87), .B(n_159), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_88), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_89), .A2(n_137), .B(n_142), .C(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_90), .Y(n_522) );
INVx1_ASAP7_75t_L g457 ( .A(n_91), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g527 ( .A(n_92), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_93), .B(n_227), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_94), .B(n_125), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_95), .B(n_125), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_96), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g149 ( .A(n_97), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_98), .A2(n_132), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
BUFx2_ASAP7_75t_L g719 ( .A(n_101), .Y(n_719) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_103), .Y(n_101) );
AND2x2_ASAP7_75t_L g429 ( .A(n_104), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AO21x2_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_113), .B(n_434), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g718 ( .A(n_112), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_424), .B(n_431), .Y(n_113) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI22xp5_ASAP7_75t_SL g436 ( .A1(n_117), .A2(n_437), .B1(n_705), .B2(n_707), .Y(n_436) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g712 ( .A(n_118), .Y(n_712) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_349), .Y(n_118) );
NOR4xp25_ASAP7_75t_L g119 ( .A(n_120), .B(n_291), .C(n_321), .D(n_331), .Y(n_119) );
OAI211xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_196), .B(n_254), .C(n_281), .Y(n_120) );
OAI222xp33_ASAP7_75t_L g376 ( .A1(n_121), .A2(n_296), .B1(n_377), .B2(n_378), .C1(n_379), .C2(n_380), .Y(n_376) );
OR2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_171), .Y(n_121) );
AOI33xp33_ASAP7_75t_L g302 ( .A1(n_122), .A2(n_289), .A3(n_290), .B1(n_303), .B2(n_308), .B3(n_310), .Y(n_302) );
OAI211xp5_ASAP7_75t_SL g359 ( .A1(n_122), .A2(n_360), .B(n_362), .C(n_364), .Y(n_359) );
OR2x2_ASAP7_75t_L g375 ( .A(n_122), .B(n_361), .Y(n_375) );
INVx1_ASAP7_75t_L g408 ( .A(n_122), .Y(n_408) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_158), .Y(n_122) );
INVx2_ASAP7_75t_L g285 ( .A(n_123), .Y(n_285) );
AND2x2_ASAP7_75t_L g301 ( .A(n_123), .B(n_187), .Y(n_301) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_123), .Y(n_336) );
AND2x2_ASAP7_75t_L g365 ( .A(n_123), .B(n_158), .Y(n_365) );
OA21x2_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_131), .B(n_155), .Y(n_123) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_124), .A2(n_188), .B(n_195), .Y(n_187) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_124), .A2(n_201), .B(n_209), .Y(n_200) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx4_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_125), .A2(n_455), .B(n_462), .Y(n_454) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g242 ( .A(n_126), .Y(n_242) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_127), .B(n_128), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
BUFx2_ASAP7_75t_L g244 ( .A(n_132), .Y(n_244) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NAND2x1p5_ASAP7_75t_L g177 ( .A(n_133), .B(n_137), .Y(n_177) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g230 ( .A(n_134), .Y(n_230) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
INVx1_ASAP7_75t_L g153 ( .A(n_135), .Y(n_153) );
INVx1_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_136), .Y(n_151) );
INVx3_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
INVx1_ASAP7_75t_L g459 ( .A(n_136), .Y(n_459) );
INVx4_ASAP7_75t_SL g154 ( .A(n_137), .Y(n_154) );
BUFx3_ASAP7_75t_L g231 ( .A(n_137), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_SL g139 ( .A1(n_140), .A2(n_141), .B(n_145), .C(n_154), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_SL g161 ( .A1(n_141), .A2(n_154), .B(n_162), .C(n_163), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_SL g189 ( .A1(n_141), .A2(n_154), .B(n_190), .C(n_191), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_141), .A2(n_154), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_SL g245 ( .A1(n_141), .A2(n_154), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_141), .A2(n_154), .B(n_457), .C(n_458), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_141), .A2(n_154), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_141), .A2(n_154), .B(n_527), .C(n_528), .Y(n_526) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx3_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_143), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_146), .B(n_206), .Y(n_205) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g164 ( .A(n_147), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_150), .B(n_193), .Y(n_192) );
OAI22xp33_ASAP7_75t_L g248 ( .A1(n_150), .A2(n_227), .B1(n_249), .B2(n_250), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_150), .B(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g182 ( .A(n_151), .Y(n_182) );
OAI22xp5_ASAP7_75t_SL g481 ( .A1(n_151), .A2(n_182), .B1(n_482), .B2(n_483), .Y(n_481) );
INVx2_ASAP7_75t_L g450 ( .A(n_152), .Y(n_450) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g217 ( .A(n_154), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g479 ( .A1(n_154), .A2(n_177), .B1(n_480), .B2(n_484), .Y(n_479) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_156), .A2(n_465), .B(n_471), .Y(n_464) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_157), .B(n_186), .Y(n_185) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_157), .A2(n_211), .B(n_218), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_157), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_SL g501 ( .A(n_157), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g265 ( .A(n_158), .Y(n_265) );
BUFx3_ASAP7_75t_L g273 ( .A(n_158), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_158), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g284 ( .A(n_158), .B(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_158), .B(n_172), .Y(n_313) );
AND2x2_ASAP7_75t_L g382 ( .A(n_158), .B(n_316), .Y(n_382) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_170), .Y(n_158) );
INVx1_ASAP7_75t_L g174 ( .A(n_159), .Y(n_174) );
INVx2_ASAP7_75t_L g220 ( .A(n_159), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_159), .A2(n_177), .B(n_223), .C(n_224), .Y(n_222) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_159), .A2(n_525), .B(n_531), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx5_ASAP7_75t_L g227 ( .A(n_167), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_167), .B(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_167), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g184 ( .A(n_168), .Y(n_184) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g194 ( .A(n_169), .Y(n_194) );
INVx2_ASAP7_75t_SL g276 ( .A(n_171), .Y(n_276) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_187), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_172), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g318 ( .A(n_172), .Y(n_318) );
AND2x2_ASAP7_75t_L g329 ( .A(n_172), .B(n_285), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_172), .B(n_314), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_172), .B(n_316), .Y(n_361) );
AND2x2_ASAP7_75t_L g420 ( .A(n_172), .B(n_365), .Y(n_420) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g290 ( .A(n_173), .B(n_187), .Y(n_290) );
AND2x2_ASAP7_75t_L g300 ( .A(n_173), .B(n_301), .Y(n_300) );
BUFx3_ASAP7_75t_L g322 ( .A(n_173), .Y(n_322) );
AND3x2_ASAP7_75t_L g381 ( .A(n_173), .B(n_382), .C(n_383), .Y(n_381) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_185), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_174), .B(n_452), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_174), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_174), .B(n_522), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_178), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_177), .A2(n_212), .B(n_213), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g444 ( .A1(n_177), .A2(n_445), .B(n_446), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_177), .A2(n_505), .B(n_506), .Y(n_504) );
O2A1O1Ixp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_183), .C(n_184), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_181), .A2(n_184), .B(n_215), .C(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_184), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_184), .A2(n_508), .B(n_509), .Y(n_507) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_187), .Y(n_272) );
INVx1_ASAP7_75t_SL g316 ( .A(n_187), .Y(n_316) );
NAND3xp33_ASAP7_75t_L g328 ( .A(n_187), .B(n_265), .C(n_329), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_234), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g351 ( .A1(n_197), .A2(n_300), .B(n_352), .C(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_199), .B(n_221), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_199), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_SL g368 ( .A(n_199), .Y(n_368) );
AND2x2_ASAP7_75t_L g389 ( .A(n_199), .B(n_236), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_199), .B(n_298), .Y(n_417) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_210), .Y(n_199) );
AND2x2_ASAP7_75t_L g262 ( .A(n_200), .B(n_253), .Y(n_262) );
INVx2_ASAP7_75t_L g269 ( .A(n_200), .Y(n_269) );
AND2x2_ASAP7_75t_L g289 ( .A(n_200), .B(n_236), .Y(n_289) );
AND2x2_ASAP7_75t_L g339 ( .A(n_200), .B(n_221), .Y(n_339) );
INVx1_ASAP7_75t_L g343 ( .A(n_200), .Y(n_343) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_208), .Y(n_519) );
INVx2_ASAP7_75t_SL g253 ( .A(n_210), .Y(n_253) );
BUFx2_ASAP7_75t_L g279 ( .A(n_210), .Y(n_279) );
AND2x2_ASAP7_75t_L g406 ( .A(n_210), .B(n_221), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx1_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_220), .A2(n_514), .B(n_521), .Y(n_513) );
INVx3_ASAP7_75t_SL g236 ( .A(n_221), .Y(n_236) );
AND2x2_ASAP7_75t_L g261 ( .A(n_221), .B(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g268 ( .A(n_221), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g298 ( .A(n_221), .B(n_258), .Y(n_298) );
OR2x2_ASAP7_75t_L g307 ( .A(n_221), .B(n_253), .Y(n_307) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_221), .Y(n_325) );
AND2x2_ASAP7_75t_L g330 ( .A(n_221), .B(n_283), .Y(n_330) );
AND2x2_ASAP7_75t_L g358 ( .A(n_221), .B(n_238), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_221), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g396 ( .A(n_221), .B(n_237), .Y(n_396) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_232), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_228), .C(n_229), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g447 ( .A1(n_227), .A2(n_448), .B(n_449), .C(n_450), .Y(n_447) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_230), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
AND2x2_ASAP7_75t_L g320 ( .A(n_236), .B(n_269), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_236), .B(n_262), .Y(n_348) );
AND2x2_ASAP7_75t_L g366 ( .A(n_236), .B(n_283), .Y(n_366) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_253), .Y(n_237) );
AND2x2_ASAP7_75t_L g267 ( .A(n_238), .B(n_253), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_238), .B(n_296), .Y(n_295) );
BUFx3_ASAP7_75t_L g305 ( .A(n_238), .Y(n_305) );
OR2x2_ASAP7_75t_L g353 ( .A(n_238), .B(n_273), .Y(n_353) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_243), .B(n_251), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_240), .A2(n_259), .B(n_260), .Y(n_258) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_240), .A2(n_504), .B(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AOI21xp5_ASAP7_75t_SL g495 ( .A1(n_241), .A2(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_242), .A2(n_444), .B(n_451), .Y(n_443) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_242), .A2(n_479), .B(n_485), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_242), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g259 ( .A(n_243), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_251), .Y(n_260) );
AND2x2_ASAP7_75t_L g288 ( .A(n_253), .B(n_258), .Y(n_288) );
INVx1_ASAP7_75t_L g296 ( .A(n_253), .Y(n_296) );
AND2x2_ASAP7_75t_L g391 ( .A(n_253), .B(n_269), .Y(n_391) );
AOI222xp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_263), .B1(n_266), .B2(n_270), .C1(n_274), .C2(n_277), .Y(n_254) );
INVx1_ASAP7_75t_L g386 ( .A(n_255), .Y(n_386) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_261), .Y(n_255) );
AND2x2_ASAP7_75t_L g282 ( .A(n_256), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g293 ( .A(n_256), .B(n_262), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_256), .B(n_284), .Y(n_309) );
OAI222xp33_ASAP7_75t_L g331 ( .A1(n_256), .A2(n_332), .B1(n_337), .B2(n_338), .C1(n_346), .C2(n_348), .Y(n_331) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g319 ( .A(n_258), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_258), .B(n_339), .Y(n_379) );
AND2x2_ASAP7_75t_L g390 ( .A(n_258), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g398 ( .A(n_261), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_263), .B(n_314), .Y(n_377) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_265), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g335 ( .A(n_265), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx3_ASAP7_75t_L g280 ( .A(n_268), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g370 ( .A1(n_268), .A2(n_371), .B(n_374), .C(n_376), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_268), .B(n_305), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_268), .B(n_288), .Y(n_410) );
AND2x2_ASAP7_75t_L g283 ( .A(n_269), .B(n_279), .Y(n_283) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g310 ( .A(n_272), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_273), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g362 ( .A(n_273), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g401 ( .A(n_273), .B(n_301), .Y(n_401) );
INVx1_ASAP7_75t_L g413 ( .A(n_273), .Y(n_413) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_276), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g394 ( .A(n_279), .Y(n_394) );
A2O1A1Ixp33_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_284), .B(n_286), .C(n_290), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_282), .A2(n_312), .B1(n_327), .B2(n_330), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_283), .B(n_297), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_283), .B(n_305), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_284), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g347 ( .A(n_284), .Y(n_347) );
AND2x2_ASAP7_75t_L g354 ( .A(n_284), .B(n_334), .Y(n_354) );
INVx2_ASAP7_75t_L g315 ( .A(n_285), .Y(n_315) );
INVxp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NOR4xp25_ASAP7_75t_L g292 ( .A(n_289), .B(n_293), .C(n_294), .D(n_297), .Y(n_292) );
INVx1_ASAP7_75t_SL g363 ( .A(n_290), .Y(n_363) );
AND2x2_ASAP7_75t_L g407 ( .A(n_290), .B(n_408), .Y(n_407) );
OAI211xp5_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_299), .B(n_302), .C(n_311), .Y(n_291) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_298), .B(n_368), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_300), .A2(n_419), .B1(n_420), .B2(n_421), .Y(n_418) );
INVx1_ASAP7_75t_SL g373 ( .A(n_301), .Y(n_373) );
AND2x2_ASAP7_75t_L g412 ( .A(n_301), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_305), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_309), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_310), .B(n_335), .Y(n_395) );
OAI21xp5_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_317), .B(n_319), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g387 ( .A(n_314), .Y(n_387) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g415 ( .A(n_315), .Y(n_415) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_316), .Y(n_342) );
OAI21xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B(n_326), .Y(n_321) );
CKINVDCx16_ASAP7_75t_R g334 ( .A(n_322), .Y(n_334) );
OR2x2_ASAP7_75t_L g372 ( .A(n_322), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI21xp33_ASAP7_75t_SL g367 ( .A1(n_325), .A2(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_329), .A2(n_356), .B1(n_359), .B2(n_366), .C(n_367), .Y(n_355) );
INVx1_ASAP7_75t_SL g399 ( .A(n_330), .Y(n_399) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OR2x2_ASAP7_75t_L g346 ( .A(n_334), .B(n_347), .Y(n_346) );
INVxp67_ASAP7_75t_L g383 ( .A(n_336), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_343), .B2(n_344), .Y(n_338) );
INVx1_ASAP7_75t_L g378 ( .A(n_339), .Y(n_378) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_342), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR4xp25_ASAP7_75t_L g349 ( .A(n_350), .B(n_384), .C(n_397), .D(n_409), .Y(n_349) );
NAND3xp33_ASAP7_75t_SL g350 ( .A(n_351), .B(n_355), .C(n_370), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_353), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_360), .B(n_365), .Y(n_369) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI221xp5_ASAP7_75t_SL g397 ( .A1(n_372), .A2(n_398), .B1(n_399), .B2(n_400), .C(n_402), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_374), .A2(n_389), .B(n_390), .C(n_392), .Y(n_388) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_375), .A2(n_393), .B1(n_395), .B2(n_396), .Y(n_392) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
A2O1A1Ixp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B(n_387), .C(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g403 ( .A(n_396), .Y(n_403) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI21xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_404), .B(n_407), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI221xp5_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_411), .B1(n_414), .B2(n_416), .C(n_418), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_427), .Y(n_433) );
NOR2x2_ASAP7_75t_L g716 ( .A(n_428), .B(n_706), .Y(n_716) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g705 ( .A(n_429), .B(n_706), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_431), .A2(n_435), .B(n_717), .Y(n_434) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g709 ( .A(n_437), .Y(n_709) );
NAND2x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_621), .Y(n_437) );
NOR5xp2_ASAP7_75t_L g438 ( .A(n_439), .B(n_544), .C(n_576), .D(n_591), .E(n_608), .Y(n_438) );
A2O1A1Ixp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_472), .B(n_491), .C(n_532), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_453), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_441), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_441), .B(n_596), .Y(n_659) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_442), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_442), .B(n_488), .Y(n_545) );
AND2x2_ASAP7_75t_L g586 ( .A(n_442), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_442), .B(n_555), .Y(n_590) );
OR2x2_ASAP7_75t_L g627 ( .A(n_442), .B(n_478), .Y(n_627) );
INVx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g477 ( .A(n_443), .B(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g535 ( .A(n_443), .Y(n_535) );
OR2x2_ASAP7_75t_L g698 ( .A(n_443), .B(n_538), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_453), .A2(n_601), .B1(n_602), .B2(n_605), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_453), .B(n_535), .Y(n_684) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_463), .Y(n_453) );
AND2x2_ASAP7_75t_L g490 ( .A(n_454), .B(n_478), .Y(n_490) );
AND2x2_ASAP7_75t_L g537 ( .A(n_454), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g542 ( .A(n_454), .Y(n_542) );
INVx3_ASAP7_75t_L g555 ( .A(n_454), .Y(n_555) );
OR2x2_ASAP7_75t_L g575 ( .A(n_454), .B(n_538), .Y(n_575) );
AND2x2_ASAP7_75t_L g594 ( .A(n_454), .B(n_464), .Y(n_594) );
BUFx2_ASAP7_75t_L g626 ( .A(n_454), .Y(n_626) );
AND2x4_ASAP7_75t_L g541 ( .A(n_463), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
BUFx2_ASAP7_75t_L g476 ( .A(n_464), .Y(n_476) );
INVx2_ASAP7_75t_L g489 ( .A(n_464), .Y(n_489) );
OR2x2_ASAP7_75t_L g557 ( .A(n_464), .B(n_538), .Y(n_557) );
AND2x2_ASAP7_75t_L g587 ( .A(n_464), .B(n_478), .Y(n_587) );
AND2x2_ASAP7_75t_L g604 ( .A(n_464), .B(n_535), .Y(n_604) );
AND2x2_ASAP7_75t_L g644 ( .A(n_464), .B(n_555), .Y(n_644) );
AND2x2_ASAP7_75t_SL g680 ( .A(n_464), .B(n_490), .Y(n_680) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp33_ASAP7_75t_SL g473 ( .A(n_474), .B(n_487), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_475), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_476), .A2(n_490), .B(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_476), .B(n_478), .Y(n_674) );
AND2x2_ASAP7_75t_L g610 ( .A(n_477), .B(n_611), .Y(n_610) );
INVx3_ASAP7_75t_L g538 ( .A(n_478), .Y(n_538) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_478), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_487), .B(n_535), .Y(n_703) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_488), .A2(n_646), .B1(n_647), .B2(n_652), .Y(n_645) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
AND2x2_ASAP7_75t_L g536 ( .A(n_489), .B(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g574 ( .A(n_489), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_SL g611 ( .A(n_489), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_490), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g665 ( .A(n_490), .Y(n_665) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_512), .Y(n_492) );
INVx4_ASAP7_75t_L g551 ( .A(n_493), .Y(n_551) );
AND2x2_ASAP7_75t_L g629 ( .A(n_493), .B(n_596), .Y(n_629) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
INVx3_ASAP7_75t_L g548 ( .A(n_494), .Y(n_548) );
AND2x2_ASAP7_75t_L g562 ( .A(n_494), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g566 ( .A(n_494), .Y(n_566) );
INVx2_ASAP7_75t_L g580 ( .A(n_494), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_494), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g637 ( .A(n_494), .B(n_632), .Y(n_637) );
AND2x2_ASAP7_75t_L g702 ( .A(n_494), .B(n_672), .Y(n_702) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_501), .Y(n_494) );
AND2x2_ASAP7_75t_L g543 ( .A(n_503), .B(n_524), .Y(n_543) );
INVx2_ASAP7_75t_L g563 ( .A(n_503), .Y(n_563) );
INVx1_ASAP7_75t_L g568 ( .A(n_512), .Y(n_568) );
AND2x2_ASAP7_75t_L g614 ( .A(n_512), .B(n_562), .Y(n_614) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_523), .Y(n_512) );
INVx2_ASAP7_75t_L g553 ( .A(n_513), .Y(n_553) );
INVx1_ASAP7_75t_L g561 ( .A(n_513), .Y(n_561) );
AND2x2_ASAP7_75t_L g579 ( .A(n_513), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_513), .B(n_563), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_520), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_519), .Y(n_516) );
AND2x2_ASAP7_75t_L g596 ( .A(n_523), .B(n_553), .Y(n_596) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g549 ( .A(n_524), .Y(n_549) );
AND2x2_ASAP7_75t_L g632 ( .A(n_524), .B(n_563), .Y(n_632) );
OAI21xp5_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_539), .B(n_543), .Y(n_532) );
INVx1_ASAP7_75t_SL g577 ( .A(n_533), .Y(n_577) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_534), .B(n_541), .Y(n_634) );
INVx1_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g583 ( .A(n_535), .B(n_538), .Y(n_583) );
AND2x2_ASAP7_75t_L g612 ( .A(n_535), .B(n_556), .Y(n_612) );
OR2x2_ASAP7_75t_L g615 ( .A(n_535), .B(n_575), .Y(n_615) );
AOI222xp33_ASAP7_75t_L g679 ( .A1(n_536), .A2(n_628), .B1(n_680), .B2(n_681), .C1(n_683), .C2(n_685), .Y(n_679) );
BUFx2_ASAP7_75t_L g593 ( .A(n_538), .Y(n_593) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g582 ( .A(n_541), .B(n_583), .Y(n_582) );
INVx3_ASAP7_75t_SL g599 ( .A(n_541), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_541), .B(n_593), .Y(n_653) );
AND2x2_ASAP7_75t_L g588 ( .A(n_543), .B(n_548), .Y(n_588) );
INVx1_ASAP7_75t_L g607 ( .A(n_543), .Y(n_607) );
OAI221xp5_ASAP7_75t_SL g544 ( .A1(n_545), .A2(n_546), .B1(n_550), .B2(n_554), .C(n_558), .Y(n_544) );
OR2x2_ASAP7_75t_L g616 ( .A(n_546), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AND2x2_ASAP7_75t_L g601 ( .A(n_548), .B(n_571), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_548), .B(n_561), .Y(n_641) );
AND2x2_ASAP7_75t_L g646 ( .A(n_548), .B(n_596), .Y(n_646) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_548), .Y(n_656) );
NAND2x1_ASAP7_75t_SL g667 ( .A(n_548), .B(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g552 ( .A(n_549), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g572 ( .A(n_549), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_549), .B(n_567), .Y(n_598) );
INVx1_ASAP7_75t_L g664 ( .A(n_549), .Y(n_664) );
INVx1_ASAP7_75t_L g639 ( .A(n_550), .Y(n_639) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g651 ( .A(n_551), .Y(n_651) );
NOR2xp67_ASAP7_75t_L g663 ( .A(n_551), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g668 ( .A(n_552), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_552), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g571 ( .A(n_553), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_553), .B(n_563), .Y(n_584) );
INVx1_ASAP7_75t_L g650 ( .A(n_553), .Y(n_650) );
INVx1_ASAP7_75t_L g671 ( .A(n_554), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI21xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_564), .B(n_573), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
AND2x2_ASAP7_75t_L g704 ( .A(n_560), .B(n_637), .Y(n_704) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g672 ( .A(n_561), .B(n_632), .Y(n_672) );
AOI32xp33_ASAP7_75t_L g585 ( .A1(n_562), .A2(n_568), .A3(n_586), .B1(n_588), .B2(n_589), .Y(n_585) );
AOI322xp5_ASAP7_75t_L g687 ( .A1(n_562), .A2(n_594), .A3(n_677), .B1(n_688), .B2(n_689), .C1(n_690), .C2(n_692), .Y(n_687) );
INVx2_ASAP7_75t_L g567 ( .A(n_563), .Y(n_567) );
INVx1_ASAP7_75t_L g677 ( .A(n_563), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .B1(n_569), .B2(n_570), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_565), .B(n_571), .Y(n_620) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_566), .B(n_632), .Y(n_682) );
INVx1_ASAP7_75t_L g569 ( .A(n_567), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_567), .B(n_596), .Y(n_686) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_575), .B(n_670), .Y(n_669) );
OAI221xp5_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_578), .B1(n_581), .B2(n_584), .C(n_585), .Y(n_576) );
OR2x2_ASAP7_75t_L g597 ( .A(n_578), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g606 ( .A(n_578), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g631 ( .A(n_579), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g635 ( .A(n_589), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_595), .B1(n_597), .B2(n_599), .C(n_600), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_593), .A2(n_624), .B1(n_628), .B2(n_629), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_594), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g699 ( .A(n_594), .Y(n_699) );
INVx1_ASAP7_75t_L g693 ( .A(n_596), .Y(n_693) );
INVx1_ASAP7_75t_SL g628 ( .A(n_597), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_599), .B(n_627), .Y(n_689) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_604), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g670 ( .A(n_604), .Y(n_670) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
OAI221xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_613), .B1(n_615), .B2(n_616), .C(n_618), .Y(n_608) );
NOR2xp33_ASAP7_75t_SL g609 ( .A(n_610), .B(n_612), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_610), .A2(n_628), .B1(n_674), .B2(n_675), .Y(n_673) );
CKINVDCx14_ASAP7_75t_R g613 ( .A(n_614), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g692 ( .A1(n_615), .A2(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR3xp33_ASAP7_75t_SL g621 ( .A(n_622), .B(n_654), .C(n_678), .Y(n_621) );
NAND4xp25_ASAP7_75t_L g622 ( .A(n_623), .B(n_630), .C(n_638), .D(n_645), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g701 ( .A(n_626), .Y(n_701) );
INVx3_ASAP7_75t_SL g695 ( .A(n_627), .Y(n_695) );
OR2x2_ASAP7_75t_L g700 ( .A(n_627), .B(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B1(n_635), .B2(n_637), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_632), .B(n_650), .Y(n_691) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_640), .B(n_642), .Y(n_638) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI211xp5_ASAP7_75t_SL g654 ( .A1(n_655), .A2(n_657), .B(n_660), .C(n_673), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g688 ( .A(n_659), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_665), .B1(n_666), .B2(n_669), .C1(n_671), .C2(n_672), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND4xp25_ASAP7_75t_SL g697 ( .A(n_670), .B(n_698), .C(n_699), .D(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND3xp33_ASAP7_75t_SL g678 ( .A(n_679), .B(n_687), .C(n_696), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_705), .A2(n_709), .B1(n_710), .B2(n_712), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_707), .Y(n_711) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
endmodule