module fake_jpeg_6087_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_30),
.B(n_33),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx12_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_1),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_28),
.B(n_29),
.C(n_15),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_50),
.Y(n_73)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_53),
.Y(n_74)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_22),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_58),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_SL g60 ( 
.A(n_53),
.B(n_37),
.C(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_63),
.B(n_65),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_39),
.B(n_36),
.C(n_34),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_72),
.B1(n_54),
.B2(n_52),
.Y(n_82)
);

FAx1_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_40),
.CI(n_25),
.CON(n_65),
.SN(n_65)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_76),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_28),
.B(n_29),
.C(n_26),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_28),
.B1(n_16),
.B2(n_24),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_17),
.B1(n_56),
.B2(n_59),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_51),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_39),
.B1(n_26),
.B2(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_25),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_82),
.B1(n_62),
.B2(n_75),
.Y(n_110)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_86),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_48),
.B1(n_46),
.B2(n_16),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_94),
.B1(n_64),
.B2(n_62),
.Y(n_104)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_17),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_64),
.B(n_71),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_16),
.B1(n_59),
.B2(n_51),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_65),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_109),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_76),
.C(n_65),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_106),
.C(n_108),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_110),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_82),
.B1(n_84),
.B2(n_94),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_68),
.C(n_67),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_68),
.C(n_63),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_64),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_64),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_85),
.C(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_81),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_116),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_86),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_121),
.C(n_108),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_78),
.C(n_77),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_75),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVxp67_ASAP7_75t_SL g134 ( 
.A(n_126),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_103),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_64),
.B1(n_89),
.B2(n_18),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_95),
.B1(n_23),
.B2(n_18),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_23),
.B1(n_27),
.B2(n_21),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_112),
.B(n_97),
.C(n_98),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_126),
.A2(n_115),
.B(n_97),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_141),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_142),
.C(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_121),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_119),
.B1(n_113),
.B2(n_122),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_142),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_117),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_117),
.C(n_127),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_154),
.C(n_155),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_23),
.C(n_21),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_159),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_134),
.B1(n_133),
.B2(n_136),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_157),
.A2(n_135),
.B1(n_21),
.B2(n_23),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_2),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_27),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_154),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_162),
.A2(n_170),
.B(n_167),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_135),
.B1(n_145),
.B2(n_132),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_172),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_146),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_143),
.C(n_135),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_159),
.C(n_147),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_171),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_175),
.C(n_179),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_163),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_153),
.B1(n_158),
.B2(n_4),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_162),
.A3(n_166),
.B1(n_165),
.B2(n_163),
.C1(n_14),
.C2(n_13),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_2),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_181),
.B(n_3),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_176),
.B(n_181),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_186),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_183),
.A2(n_185),
.B(n_174),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_162),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_6),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_13),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_187),
.B(n_5),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_194),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_173),
.B1(n_179),
.B2(n_7),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_193),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_27),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_189),
.C(n_193),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_198),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_6),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_8),
.B(n_9),
.C(n_10),
.D(n_11),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_195),
.C(n_10),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_9),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);


endmodule