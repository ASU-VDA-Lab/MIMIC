module fake_jpeg_25828_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_46),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_56),
.Y(n_73)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_19),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_27),
.B1(n_22),
.B2(n_25),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_22),
.B1(n_36),
.B2(n_25),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_68),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_22),
.B1(n_25),
.B2(n_30),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_30),
.B1(n_40),
.B2(n_21),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_17),
.B(n_33),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_44),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_70),
.A2(n_78),
.B1(n_94),
.B2(n_32),
.Y(n_119)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_22),
.B1(n_53),
.B2(n_55),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_60),
.B1(n_53),
.B2(n_49),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_36),
.B1(n_40),
.B2(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_81),
.B(n_88),
.Y(n_128)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_99),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_93),
.B1(n_96),
.B2(n_60),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_50),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_86),
.Y(n_123)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_90),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_97),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_30),
.B1(n_34),
.B2(n_21),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_34),
.B1(n_32),
.B2(n_26),
.Y(n_110)
);

BUFx12f_ASAP7_75t_SL g93 ( 
.A(n_54),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_30),
.B1(n_19),
.B2(n_34),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_88),
.B(n_73),
.Y(n_120)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_20),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_55),
.C(n_41),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_105),
.C(n_38),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

AOI22x1_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_43),
.B1(n_44),
.B2(n_41),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_103),
.A2(n_80),
.B1(n_87),
.B2(n_38),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_21),
.Y(n_105)
);

NOR2x1p5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_109),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_53),
.B1(n_17),
.B2(n_33),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_119),
.B1(n_129),
.B2(n_71),
.Y(n_135)
);

AND2x4_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_49),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_122),
.B1(n_94),
.B2(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_35),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_76),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_20),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_32),
.B1(n_18),
.B2(n_26),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_78),
.A2(n_70),
.B1(n_97),
.B2(n_90),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_23),
.B1(n_18),
.B2(n_35),
.Y(n_154)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_69),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_18),
.B1(n_23),
.B2(n_26),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_135),
.B1(n_111),
.B2(n_125),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_114),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_72),
.Y(n_137)
);

OR2x2_ASAP7_75t_SL g138 ( 
.A(n_101),
.B(n_86),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_138),
.A2(n_139),
.B(n_148),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_98),
.C(n_76),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_109),
.C(n_123),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_142),
.Y(n_171)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_89),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_145),
.Y(n_162)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

AOI21x1_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_52),
.B(n_115),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_144),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_85),
.B(n_31),
.C(n_52),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_105),
.B(n_12),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_85),
.B1(n_26),
.B2(n_23),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_151),
.A2(n_152),
.B1(n_124),
.B2(n_125),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_23),
.B1(n_18),
.B2(n_35),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_111),
.B(n_109),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_155),
.B1(n_122),
.B2(n_110),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_119),
.B1(n_103),
.B2(n_109),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_101),
.A2(n_20),
.B1(n_31),
.B2(n_24),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_160),
.A2(n_172),
.B(n_177),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_163),
.A2(n_190),
.B1(n_31),
.B2(n_7),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_170),
.C(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_167),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_176),
.B1(n_180),
.B2(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_123),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_12),
.C(n_15),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_168),
.B(n_182),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_113),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_114),
.B(n_121),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_121),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_181),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_113),
.C(n_115),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_130),
.B1(n_155),
.B2(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_8),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_183),
.Y(n_195)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_31),
.B(n_24),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_156),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_189),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_52),
.B1(n_31),
.B2(n_2),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_146),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_206),
.B(n_174),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_193),
.A2(n_221),
.B1(n_175),
.B2(n_188),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_157),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_196),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_203),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_183),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_201),
.B(n_202),
.Y(n_248)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_131),
.C(n_158),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_209),
.C(n_199),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_146),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_131),
.C(n_141),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_142),
.B1(n_31),
.B2(n_24),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_210),
.A2(n_185),
.B1(n_186),
.B2(n_188),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_24),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_191),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_161),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_184),
.B1(n_192),
.B2(n_217),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_187),
.Y(n_228)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_187),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_7),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_11),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_222),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_15),
.B1(n_13),
.B2(n_11),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_223),
.A2(n_242),
.B1(n_244),
.B2(n_208),
.Y(n_269)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_224),
.B(n_227),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_231),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_232),
.B(n_236),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_207),
.A2(n_191),
.B(n_169),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_239),
.B1(n_246),
.B2(n_247),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_238),
.C(n_211),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_169),
.C(n_174),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_163),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_193),
.Y(n_251)
);

OAI21x1_ASAP7_75t_R g243 ( 
.A1(n_195),
.A2(n_172),
.B(n_1),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_243),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_194),
.B(n_173),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_0),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_250),
.C(n_261),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_206),
.C(n_212),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_254),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_219),
.B1(n_213),
.B2(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_232),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_206),
.B1(n_222),
.B2(n_231),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_263),
.B1(n_260),
.B2(n_266),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_207),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_13),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_201),
.C(n_202),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_203),
.C(n_213),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_210),
.C(n_195),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_208),
.C(n_220),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_269),
.A2(n_233),
.B(n_245),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_274),
.B(n_281),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_223),
.B1(n_224),
.B2(n_227),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_277),
.B1(n_288),
.B2(n_261),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_252),
.A2(n_243),
.B1(n_245),
.B2(n_240),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_286),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_226),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_280),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_257),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_248),
.C(n_243),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_251),
.C(n_255),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_248),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_270),
.A2(n_13),
.B(n_11),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_258),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_262),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_259),
.C(n_254),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_289),
.A2(n_283),
.B(n_271),
.Y(n_310)
);

BUFx12_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_267),
.C(n_264),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_292),
.A2(n_278),
.B(n_275),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_282),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_300),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_250),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_271),
.C(n_300),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_283),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_310),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_311),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_R g306 ( 
.A(n_293),
.B(n_274),
.C(n_295),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_306),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_276),
.B(n_284),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_10),
.B(n_9),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_299),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_10),
.C(n_8),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_1),
.C(n_2),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_298),
.B(n_294),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_4),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_291),
.B1(n_290),
.B2(n_10),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_317),
.B(n_319),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_291),
.Y(n_319)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_1),
.C(n_3),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_304),
.C(n_5),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_314),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_5),
.Y(n_332)
);

AOI31xp67_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_307),
.A3(n_313),
.B(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_328),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_4),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_332),
.C(n_321),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_330),
.B(n_331),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_333),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_334),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_326),
.C(n_320),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_323),
.B(n_322),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_323),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_5),
.B(n_6),
.Y(n_342)
);


endmodule