module fake_jpeg_7644_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_35),
.B(n_41),
.Y(n_66)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_44),
.B1(n_28),
.B2(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_3),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_27),
.B1(n_26),
.B2(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_27),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_67),
.Y(n_89)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_18),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_65),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_16),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_16),
.B(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_66),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_36),
.B1(n_28),
.B2(n_34),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_69),
.A2(n_80),
.B1(n_26),
.B2(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_91),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_36),
.C(n_34),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_78),
.C(n_81),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_22),
.C(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_84),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_22),
.C(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_17),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_21),
.Y(n_110)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_51),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVxp33_ASAP7_75t_SL g113 ( 
.A(n_96),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_111),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_88),
.B1(n_85),
.B2(n_70),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_66),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_76),
.C(n_69),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_55),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_46),
.B(n_53),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_108),
.B(n_110),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_56),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_58),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_71),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_118),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_74),
.B(n_85),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_100),
.B(n_105),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_100),
.C(n_97),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_128),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_108),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_135),
.B(n_138),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_126),
.C(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

NOR4xp25_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_104),
.C(n_110),
.D(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_103),
.C(n_89),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_108),
.B(n_109),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_101),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_131),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_148),
.C(n_151),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_125),
.C(n_121),
.Y(n_148)
);

AOI321xp33_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_131),
.A3(n_133),
.B1(n_120),
.B2(n_92),
.C(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_150),
.B(n_145),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_122),
.C(n_123),
.Y(n_151)
);

XOR2x2_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_142),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_155),
.B1(n_149),
.B2(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_159),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_139),
.B(n_116),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_154),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_137),
.A3(n_70),
.B1(n_90),
.B2(n_62),
.C1(n_84),
.C2(n_79),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_161),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_147),
.A2(n_90),
.B1(n_74),
.B2(n_106),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_144),
.C(n_148),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_166),
.B(n_62),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_167),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_158),
.B(n_153),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_168),
.B(n_163),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_155),
.B(n_6),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_169),
.A2(n_171),
.B(n_172),
.Y(n_174)
);

OAI31xp33_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_62),
.A3(n_7),
.B(n_8),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_175),
.C(n_10),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_58),
.A3(n_10),
.B1(n_12),
.B2(n_15),
.C1(n_25),
.C2(n_21),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_177),
.C(n_15),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_58),
.C(n_12),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_5),
.Y(n_179)
);


endmodule