module real_aes_17065_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_1638;
wire n_495;
wire n_1072;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1679;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1647;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_0), .A2(n_79), .B1(n_927), .B2(n_932), .Y(n_931) );
INVxp33_ASAP7_75t_SL g965 ( .A(n_0), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g1433 ( .A1(n_1), .A2(n_230), .B1(n_1406), .B2(n_1410), .Y(n_1433) );
AOI221xp5_ASAP7_75t_L g1172 ( .A1(n_2), .A2(n_62), .B1(n_821), .B2(n_1153), .C(n_1173), .Y(n_1172) );
AOI22xp33_ASAP7_75t_SL g1186 ( .A1(n_2), .A2(n_205), .B1(n_1187), .B2(n_1189), .Y(n_1186) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_3), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g1269 ( .A1(n_4), .A2(n_235), .B1(n_476), .B2(n_945), .C(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1296 ( .A(n_4), .Y(n_1296) );
OAI22xp5_ASAP7_75t_L g1177 ( .A1(n_5), .A2(n_112), .B1(n_737), .B2(n_765), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1442 ( .A1(n_6), .A2(n_243), .B1(n_1406), .B2(n_1410), .Y(n_1442) );
INVx1_ASAP7_75t_L g1271 ( .A(n_7), .Y(n_1271) );
AOI221xp5_ASAP7_75t_L g1298 ( .A1(n_7), .A2(n_171), .B1(n_805), .B2(n_1154), .C(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g878 ( .A(n_8), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_8), .A2(n_130), .B1(n_628), .B2(n_724), .Y(n_910) );
AOI221xp5_ASAP7_75t_L g1152 ( .A1(n_9), .A2(n_66), .B1(n_1022), .B2(n_1153), .C(n_1155), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_9), .A2(n_34), .B1(n_772), .B2(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1235 ( .A(n_10), .Y(n_1235) );
OAI221xp5_ASAP7_75t_L g868 ( .A1(n_11), .A2(n_245), .B1(n_461), .B2(n_582), .C(n_761), .Y(n_868) );
OA222x2_ASAP7_75t_L g912 ( .A1(n_11), .A2(n_53), .B1(n_248), .B2(n_797), .C1(n_913), .C2(n_914), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_12), .A2(n_20), .B1(n_639), .B2(n_642), .Y(n_638) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_12), .A2(n_20), .B1(n_672), .B2(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g1160 ( .A(n_13), .Y(n_1160) );
OAI22xp33_ASAP7_75t_L g1196 ( .A1(n_13), .A2(n_33), .B1(n_1197), .B2(n_1200), .Y(n_1196) );
INVx1_ASAP7_75t_L g312 ( .A(n_14), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_14), .B(n_322), .Y(n_340) );
AND2x2_ASAP7_75t_L g387 ( .A(n_14), .B(n_255), .Y(n_387) );
AND2x2_ASAP7_75t_L g411 ( .A(n_14), .B(n_412), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g1371 ( .A1(n_15), .A2(n_221), .B1(n_476), .B2(n_1005), .C(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1397 ( .A(n_15), .Y(n_1397) );
INVx1_ASAP7_75t_L g599 ( .A(n_16), .Y(n_599) );
INVx1_ASAP7_75t_L g811 ( .A(n_17), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_17), .A2(n_282), .B1(n_458), .B2(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g1118 ( .A(n_18), .Y(n_1118) );
AOI22xp5_ASAP7_75t_L g1136 ( .A1(n_18), .A2(n_38), .B1(n_1137), .B2(n_1138), .Y(n_1136) );
INVx2_ASAP7_75t_L g1409 ( .A(n_19), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_19), .B(n_123), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_19), .B(n_1415), .Y(n_1417) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_21), .Y(n_707) );
AOI22xp33_ASAP7_75t_SL g780 ( .A1(n_21), .A2(n_194), .B1(n_781), .B2(n_782), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g1427 ( .A1(n_22), .A2(n_32), .B1(n_1413), .B2(n_1416), .Y(n_1427) );
XOR2xp5_ASAP7_75t_L g1264 ( .A(n_23), .B(n_1265), .Y(n_1264) );
CKINVDCx5p33_ASAP7_75t_R g1001 ( .A(n_24), .Y(n_1001) );
XNOR2xp5_ASAP7_75t_L g1308 ( .A(n_25), .B(n_1309), .Y(n_1308) );
AOI22xp5_ASAP7_75t_L g1432 ( .A1(n_26), .A2(n_144), .B1(n_1413), .B2(n_1416), .Y(n_1432) );
INVx1_ASAP7_75t_L g1076 ( .A(n_27), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g934 ( .A1(n_28), .A2(n_86), .B1(n_833), .B2(n_836), .C(n_935), .Y(n_934) );
AOI22xp33_ASAP7_75t_SL g971 ( .A1(n_28), .A2(n_30), .B1(n_557), .B2(n_808), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g1638 ( .A(n_29), .Y(n_1638) );
AOI22xp33_ASAP7_75t_SL g924 ( .A1(n_30), .A2(n_159), .B1(n_925), .B2(n_927), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_31), .Y(n_369) );
XOR2x2_ASAP7_75t_L g684 ( .A(n_32), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g1162 ( .A(n_33), .Y(n_1162) );
INVxp67_ASAP7_75t_SL g1169 ( .A(n_34), .Y(n_1169) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_35), .A2(n_134), .B1(n_765), .B2(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g794 ( .A(n_36), .Y(n_794) );
INVx1_ASAP7_75t_L g938 ( .A(n_37), .Y(n_938) );
OA222x2_ASAP7_75t_L g952 ( .A1(n_37), .A2(n_190), .B1(n_294), .B2(n_797), .C1(n_914), .C2(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g1126 ( .A(n_38), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1491 ( .A1(n_39), .A2(n_117), .B1(n_1406), .B2(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_L g1123 ( .A(n_40), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_40), .A2(n_199), .B1(n_805), .B2(n_1137), .Y(n_1142) );
INVx1_ASAP7_75t_L g1272 ( .A(n_41), .Y(n_1272) );
AOI221xp5_ASAP7_75t_L g1290 ( .A1(n_41), .A2(n_84), .B1(n_1291), .B2(n_1293), .C(n_1295), .Y(n_1290) );
AOI221xp5_ASAP7_75t_L g928 ( .A1(n_42), .A2(n_234), .B1(n_834), .B2(n_929), .C(n_930), .Y(n_928) );
INVx1_ASAP7_75t_L g968 ( .A(n_42), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g1419 ( .A1(n_43), .A2(n_105), .B1(n_1406), .B2(n_1420), .Y(n_1419) );
AOI211xp5_ASAP7_75t_L g1363 ( .A1(n_44), .A2(n_833), .B(n_1364), .C(n_1366), .Y(n_1363) );
INVx1_ASAP7_75t_L g1393 ( .A(n_44), .Y(n_1393) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_45), .A2(n_205), .B1(n_816), .B2(n_1158), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_45), .A2(n_62), .B1(n_1191), .B2(n_1192), .Y(n_1190) );
INVx1_ASAP7_75t_L g1146 ( .A(n_46), .Y(n_1146) );
OAI221xp5_ASAP7_75t_L g1281 ( .A1(n_47), .A2(n_72), .B1(n_458), .B2(n_462), .C(n_469), .Y(n_1281) );
INVxp67_ASAP7_75t_SL g1286 ( .A(n_47), .Y(n_1286) );
OAI21xp33_ASAP7_75t_L g796 ( .A1(n_48), .A2(n_797), .B(n_799), .Y(n_796) );
OAI221xp5_ASAP7_75t_L g841 ( .A1(n_48), .A2(n_59), .B1(n_842), .B2(n_843), .C(n_844), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g541 ( .A1(n_49), .A2(n_187), .B1(n_458), .B2(n_462), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_49), .A2(n_89), .B1(n_382), .B2(n_391), .Y(n_566) );
INVxp67_ASAP7_75t_SL g701 ( .A(n_50), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g770 ( .A1(n_50), .A2(n_52), .B1(n_771), .B2(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g434 ( .A(n_51), .Y(n_434) );
INVx1_ASAP7_75t_L g448 ( .A(n_51), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_52), .A2(n_194), .B1(n_717), .B2(n_718), .C(n_722), .Y(n_716) );
INVx1_ASAP7_75t_L g867 ( .A(n_53), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g1438 ( .A1(n_54), .A2(n_153), .B1(n_1406), .B2(n_1420), .Y(n_1438) );
OAI221xp5_ASAP7_75t_L g1360 ( .A1(n_55), .A2(n_274), .B1(n_458), .B2(n_462), .C(n_469), .Y(n_1360) );
OAI22xp5_ASAP7_75t_L g1383 ( .A1(n_55), .A2(n_148), .B1(n_384), .B2(n_738), .Y(n_1383) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_56), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_57), .Y(n_374) );
INVx1_ASAP7_75t_L g813 ( .A(n_58), .Y(n_813) );
INVxp67_ASAP7_75t_SL g848 ( .A(n_59), .Y(n_848) );
INVx1_ASAP7_75t_L g1067 ( .A(n_60), .Y(n_1067) );
OAI221xp5_ASAP7_75t_L g1107 ( .A1(n_61), .A2(n_124), .B1(n_497), .B2(n_990), .C(n_1108), .Y(n_1107) );
INVxp67_ASAP7_75t_SL g1131 ( .A(n_61), .Y(n_1131) );
INVx1_ASAP7_75t_L g631 ( .A(n_63), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g1493 ( .A1(n_64), .A2(n_251), .B1(n_1413), .B2(n_1416), .Y(n_1493) );
INVx1_ASAP7_75t_L g305 ( .A(n_65), .Y(n_305) );
AOI22xp33_ASAP7_75t_SL g1195 ( .A1(n_66), .A2(n_99), .B1(n_771), .B2(n_772), .Y(n_1195) );
INVx2_ASAP7_75t_L g437 ( .A(n_67), .Y(n_437) );
INVx1_ASAP7_75t_L g1234 ( .A(n_68), .Y(n_1234) );
OAI322xp33_ASAP7_75t_L g1238 ( .A1(n_68), .A2(n_1239), .A3(n_1244), .B1(n_1245), .B2(n_1248), .C1(n_1253), .C2(n_1255), .Y(n_1238) );
OAI22xp5_ASAP7_75t_L g1280 ( .A1(n_69), .A2(n_242), .B1(n_497), .B2(n_990), .Y(n_1280) );
INVx1_ASAP7_75t_L g1289 ( .A(n_69), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1268 ( .A1(n_70), .A2(n_215), .B1(n_1078), .B2(n_1079), .Y(n_1268) );
INVx1_ASAP7_75t_L g1287 ( .A(n_70), .Y(n_1287) );
INVx1_ASAP7_75t_L g526 ( .A(n_71), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_71), .A2(n_250), .B1(n_413), .B2(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g1307 ( .A(n_72), .Y(n_1307) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_73), .Y(n_539) );
OAI21xp5_ASAP7_75t_SL g987 ( .A1(n_74), .A2(n_950), .B(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g1014 ( .A(n_74), .Y(n_1014) );
INVx1_ASAP7_75t_L g581 ( .A(n_75), .Y(n_581) );
INVx1_ASAP7_75t_L g589 ( .A(n_76), .Y(n_589) );
INVx1_ASAP7_75t_L g578 ( .A(n_77), .Y(n_578) );
INVx1_ASAP7_75t_L g416 ( .A(n_78), .Y(n_416) );
INVxp67_ASAP7_75t_SL g970 ( .A(n_79), .Y(n_970) );
AOI21xp33_ASAP7_75t_L g1071 ( .A1(n_80), .A2(n_529), .B(n_834), .Y(n_1071) );
INVxp67_ASAP7_75t_L g1093 ( .A(n_80), .Y(n_1093) );
AOI221xp5_ASAP7_75t_L g1228 ( .A1(n_81), .A2(n_198), .B1(n_960), .B2(n_1155), .C(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1247 ( .A(n_81), .Y(n_1247) );
INVx1_ASAP7_75t_L g1315 ( .A(n_82), .Y(n_1315) );
OAI211xp5_ASAP7_75t_L g624 ( .A1(n_83), .A2(n_563), .B(n_625), .C(n_630), .Y(n_624) );
INVx1_ASAP7_75t_L g670 ( .A(n_83), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_84), .A2(n_236), .B1(n_476), .B2(n_1274), .C(n_1275), .Y(n_1273) );
INVx1_ASAP7_75t_L g1643 ( .A(n_85), .Y(n_1643) );
AOI22xp5_ASAP7_75t_L g1657 ( .A1(n_85), .A2(n_119), .B1(n_808), .B2(n_1658), .Y(n_1657) );
AOI221xp5_ASAP7_75t_L g958 ( .A1(n_86), .A2(n_234), .B1(n_959), .B2(n_960), .C(n_961), .Y(n_958) );
CKINVDCx5p33_ASAP7_75t_R g872 ( .A(n_87), .Y(n_872) );
INVx1_ASAP7_75t_L g881 ( .A(n_88), .Y(n_881) );
AOI221x1_ASAP7_75t_SL g901 ( .A1(n_88), .A2(n_108), .B1(n_413), .B2(n_718), .C(n_902), .Y(n_901) );
OAI221xp5_ASAP7_75t_L g535 ( .A1(n_89), .A2(n_186), .B1(n_536), .B2(n_537), .C(n_538), .Y(n_535) );
OAI222xp33_ASAP7_75t_L g440 ( .A1(n_90), .A2(n_147), .B1(n_267), .B2(n_441), .C1(n_443), .C2(n_450), .Y(n_440) );
INVx1_ASAP7_75t_L g503 ( .A(n_90), .Y(n_503) );
INVx1_ASAP7_75t_L g584 ( .A(n_91), .Y(n_584) );
INVx1_ASAP7_75t_L g944 ( .A(n_92), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g949 ( .A(n_92), .B(n_950), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_93), .A2(n_200), .B1(n_497), .B2(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g1039 ( .A(n_93), .Y(n_1039) );
INVx1_ASAP7_75t_L g1124 ( .A(n_94), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_94), .A2(n_257), .B1(n_413), .B2(n_557), .Y(n_1139) );
OAI221xp5_ASAP7_75t_L g1321 ( .A1(n_95), .A2(n_172), .B1(n_1167), .B2(n_1322), .C(n_1323), .Y(n_1321) );
OAI22xp33_ASAP7_75t_L g1343 ( .A1(n_95), .A2(n_172), .B1(n_1344), .B2(n_1346), .Y(n_1343) );
XOR2x2_ASAP7_75t_L g1355 ( .A(n_96), .B(n_1356), .Y(n_1355) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_97), .A2(n_128), .B1(n_1406), .B2(n_1410), .Y(n_1405) );
AOI22xp5_ASAP7_75t_L g1458 ( .A1(n_98), .A2(n_145), .B1(n_1413), .B2(n_1416), .Y(n_1458) );
INVxp67_ASAP7_75t_SL g1171 ( .A(n_99), .Y(n_1171) );
CKINVDCx5p33_ASAP7_75t_R g1114 ( .A(n_100), .Y(n_1114) );
INVx1_ASAP7_75t_L g734 ( .A(n_101), .Y(n_734) );
INVx1_ASAP7_75t_L g863 ( .A(n_102), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_102), .A2(n_245), .B1(n_382), .B2(n_391), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_103), .A2(n_207), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
INVxp67_ASAP7_75t_SL g1082 ( .A(n_103), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g1370 ( .A1(n_104), .A2(n_148), .B1(n_1078), .B2(n_1079), .Y(n_1370) );
OAI211xp5_ASAP7_75t_L g1376 ( .A1(n_104), .A2(n_950), .B(n_1377), .C(n_1380), .Y(n_1376) );
INVx1_ASAP7_75t_L g373 ( .A(n_106), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_106), .A2(n_170), .B1(n_473), .B2(n_476), .C(n_478), .Y(n_472) );
INVx1_ASAP7_75t_L g946 ( .A(n_107), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_107), .A2(n_210), .B1(n_384), .B2(n_738), .Y(n_974) );
INVx1_ASAP7_75t_L g896 ( .A(n_108), .Y(n_896) );
INVx1_ASAP7_75t_L g1369 ( .A(n_109), .Y(n_1369) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_110), .Y(n_307) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_110), .B(n_305), .Y(n_1407) );
INVx1_ASAP7_75t_L g592 ( .A(n_111), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g1150 ( .A1(n_112), .A2(n_713), .B(n_1151), .C(n_1159), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_113), .A2(n_141), .B1(n_724), .B2(n_726), .Y(n_1218) );
INVxp33_ASAP7_75t_L g1246 ( .A(n_113), .Y(n_1246) );
CKINVDCx5p33_ASAP7_75t_R g1324 ( .A(n_114), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_115), .A2(n_118), .B1(n_724), .B2(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1251 ( .A(n_115), .Y(n_1251) );
INVx1_ASAP7_75t_L g1374 ( .A(n_116), .Y(n_1374) );
INVxp67_ASAP7_75t_L g1243 ( .A(n_118), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1633 ( .A1(n_119), .A2(n_181), .B1(n_935), .B2(n_1192), .Y(n_1633) );
CKINVDCx5p33_ASAP7_75t_R g1642 ( .A(n_120), .Y(n_1642) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_121), .A2(n_209), .B1(n_720), .B2(n_805), .Y(n_804) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_121), .A2(n_193), .B1(n_775), .B2(n_833), .C(n_834), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g1320 ( .A1(n_122), .A2(n_211), .B1(n_808), .B2(n_1144), .Y(n_1320) );
INVx1_ASAP7_75t_L g1336 ( .A(n_122), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_123), .B(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1415 ( .A(n_123), .Y(n_1415) );
INVx1_ASAP7_75t_L g1145 ( .A(n_124), .Y(n_1145) );
AOI22xp5_ASAP7_75t_L g1437 ( .A1(n_125), .A2(n_191), .B1(n_1413), .B2(n_1416), .Y(n_1437) );
AOI22xp5_ASAP7_75t_L g1611 ( .A1(n_125), .A2(n_1612), .B1(n_1613), .B2(n_1665), .Y(n_1611) );
INVx1_ASAP7_75t_L g1665 ( .A(n_125), .Y(n_1665) );
AOI22xp5_ASAP7_75t_L g1671 ( .A1(n_125), .A2(n_1672), .B1(n_1677), .B2(n_1680), .Y(n_1671) );
OAI221xp5_ASAP7_75t_SL g1165 ( .A1(n_126), .A2(n_152), .B1(n_688), .B2(n_1166), .C(n_1168), .Y(n_1165) );
INVx1_ASAP7_75t_L g1182 ( .A(n_126), .Y(n_1182) );
CKINVDCx5p33_ASAP7_75t_R g752 ( .A(n_127), .Y(n_752) );
INVx1_ASAP7_75t_L g1373 ( .A(n_129), .Y(n_1373) );
INVx1_ASAP7_75t_L g887 ( .A(n_130), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_131), .A2(n_291), .B1(n_724), .B2(n_726), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_131), .A2(n_176), .B1(n_775), .B2(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g994 ( .A(n_132), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_132), .A2(n_208), .B1(n_391), .B2(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1207 ( .A(n_133), .Y(n_1207) );
OAI211xp5_ASAP7_75t_SL g1311 ( .A1(n_134), .A2(n_1312), .B(n_1314), .C(n_1317), .Y(n_1311) );
INVx2_ASAP7_75t_L g439 ( .A(n_135), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_135), .B(n_437), .Y(n_456) );
INVx1_ASAP7_75t_L g489 ( .A(n_135), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_136), .Y(n_519) );
INVx1_ASAP7_75t_L g419 ( .A(n_137), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_137), .A2(n_177), .B1(n_458), .B2(n_462), .Y(n_457) );
OAI211xp5_ASAP7_75t_L g992 ( .A1(n_138), .A2(n_469), .B(n_846), .C(n_993), .Y(n_992) );
CKINVDCx5p33_ASAP7_75t_R g1044 ( .A(n_138), .Y(n_1044) );
INVx1_ASAP7_75t_L g1069 ( .A(n_139), .Y(n_1069) );
AOI221xp5_ASAP7_75t_L g1214 ( .A1(n_140), .A2(n_202), .B1(n_698), .B2(n_717), .C(n_1215), .Y(n_1214) );
INVxp67_ASAP7_75t_L g1250 ( .A(n_140), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_141), .A2(n_198), .B1(n_771), .B2(n_929), .Y(n_1252) );
INVx1_ASAP7_75t_L g1349 ( .A(n_142), .Y(n_1349) );
AOI221xp5_ASAP7_75t_L g1003 ( .A1(n_143), .A2(n_281), .B1(n_834), .B2(n_1004), .C(n_1005), .Y(n_1003) );
AOI221xp5_ASAP7_75t_SL g1030 ( .A1(n_143), .A2(n_146), .B1(n_1022), .B2(n_1031), .C(n_1032), .Y(n_1030) );
XOR2xp5_ASAP7_75t_L g854 ( .A(n_144), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g1009 ( .A(n_146), .Y(n_1009) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_147), .A2(n_177), .B1(n_382), .B2(n_391), .C(n_396), .Y(n_381) );
INVx1_ASAP7_75t_L g331 ( .A(n_149), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g806 ( .A1(n_150), .A2(n_284), .B1(n_807), .B2(n_808), .Y(n_806) );
AOI221xp5_ASAP7_75t_L g835 ( .A1(n_150), .A2(n_241), .B1(n_771), .B2(n_833), .C(n_836), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_151), .A2(n_985), .B1(n_986), .B2(n_1048), .Y(n_984) );
INVx1_ASAP7_75t_L g1048 ( .A(n_151), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1412 ( .A1(n_151), .A2(n_268), .B1(n_1413), .B2(n_1416), .Y(n_1412) );
INVx1_ASAP7_75t_L g1181 ( .A(n_152), .Y(n_1181) );
AOI22xp5_ASAP7_75t_L g1457 ( .A1(n_154), .A2(n_157), .B1(n_1406), .B2(n_1410), .Y(n_1457) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_155), .Y(n_883) );
INVx1_ASAP7_75t_L g1127 ( .A(n_156), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_156), .A2(n_214), .B1(n_727), .B2(n_1144), .Y(n_1143) );
OAI22xp33_ASAP7_75t_L g645 ( .A1(n_158), .A2(n_201), .B1(n_646), .B2(n_647), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_158), .A2(n_201), .B1(n_654), .B2(n_655), .Y(n_653) );
INVxp67_ASAP7_75t_SL g962 ( .A(n_159), .Y(n_962) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_160), .A2(n_167), .B1(n_486), .B2(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g917 ( .A(n_160), .Y(n_917) );
INVx1_ASAP7_75t_L g1221 ( .A(n_161), .Y(n_1221) );
INVx1_ASAP7_75t_L g586 ( .A(n_162), .Y(n_586) );
INVx1_ASAP7_75t_L g1279 ( .A(n_163), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1441 ( .A1(n_164), .A2(n_165), .B1(n_1413), .B2(n_1416), .Y(n_1441) );
XOR2x2_ASAP7_75t_L g1052 ( .A(n_165), .B(n_1053), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_166), .A2(n_497), .B1(n_523), .B2(n_527), .Y(n_522) );
INVx1_ASAP7_75t_L g549 ( .A(n_166), .Y(n_549) );
INVx1_ASAP7_75t_L g916 ( .A(n_167), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g1361 ( .A1(n_168), .A2(n_174), .B1(n_497), .B2(n_990), .Y(n_1361) );
INVxp67_ASAP7_75t_SL g1381 ( .A(n_168), .Y(n_1381) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_169), .A2(n_240), .B1(n_807), .B2(n_816), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_169), .A2(n_284), .B1(n_516), .B2(n_771), .Y(n_831) );
INVx1_ASAP7_75t_L g342 ( .A(n_170), .Y(n_342) );
INVx1_ASAP7_75t_L g1276 ( .A(n_171), .Y(n_1276) );
INVx1_ASAP7_75t_L g695 ( .A(n_173), .Y(n_695) );
AOI22xp33_ASAP7_75t_SL g778 ( .A1(n_173), .A2(n_291), .B1(n_777), .B2(n_779), .Y(n_778) );
INVxp67_ASAP7_75t_SL g1378 ( .A(n_174), .Y(n_1378) );
BUFx3_ASAP7_75t_L g431 ( .A(n_175), .Y(n_431) );
INVx1_ASAP7_75t_L g696 ( .A(n_176), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g1421 ( .A1(n_178), .A2(n_180), .B1(n_1413), .B2(n_1416), .Y(n_1421) );
INVx1_ASAP7_75t_L g1056 ( .A(n_179), .Y(n_1056) );
AOI22xp33_ASAP7_75t_SL g1651 ( .A1(n_181), .A2(n_263), .B1(n_1652), .B2(n_1653), .Y(n_1651) );
AOI22xp33_ASAP7_75t_SL g1327 ( .A1(n_182), .A2(n_273), .B1(n_1328), .B2(n_1329), .Y(n_1327) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_182), .A2(n_278), .B1(n_771), .B2(n_773), .Y(n_1337) );
INVx1_ASAP7_75t_L g1365 ( .A(n_183), .Y(n_1365) );
AOI22xp5_ASAP7_75t_L g1428 ( .A1(n_184), .A2(n_256), .B1(n_1406), .B2(n_1410), .Y(n_1428) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_185), .Y(n_319) );
OAI211xp5_ASAP7_75t_L g546 ( .A1(n_186), .A2(n_547), .B(n_548), .C(n_551), .Y(n_546) );
INVx1_ASAP7_75t_L g550 ( .A(n_187), .Y(n_550) );
OAI21xp5_ASAP7_75t_SL g736 ( .A1(n_188), .A2(n_737), .B(n_741), .Y(n_736) );
INVx1_ASAP7_75t_L g800 ( .A(n_189), .Y(n_800) );
INVx1_ASAP7_75t_L g948 ( .A(n_190), .Y(n_948) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_192), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_193), .A2(n_241), .B1(n_820), .B2(n_821), .Y(n_819) );
AOI221xp5_ASAP7_75t_L g1011 ( .A1(n_195), .A2(n_239), .B1(n_833), .B2(n_836), .C(n_1012), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_195), .A2(n_281), .B1(n_820), .B2(n_1022), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g1061 ( .A1(n_196), .A2(n_771), .B(n_836), .Y(n_1061) );
INVxp67_ASAP7_75t_SL g1090 ( .A(n_196), .Y(n_1090) );
XOR2xp5_ASAP7_75t_L g1147 ( .A(n_197), .B(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1117 ( .A(n_199), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_200), .Y(n_1029) );
INVxp67_ASAP7_75t_L g1240 ( .A(n_202), .Y(n_1240) );
INVx1_ASAP7_75t_L g1628 ( .A(n_203), .Y(n_1628) );
OAI221xp5_ASAP7_75t_L g1654 ( .A1(n_203), .A2(n_904), .B1(n_914), .B2(n_1655), .C(n_1660), .Y(n_1654) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_204), .Y(n_366) );
INVx1_ASAP7_75t_L g532 ( .A(n_206), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_206), .A2(n_218), .B1(n_557), .B2(n_565), .Y(n_564) );
OAI221xp5_ASAP7_75t_L g1099 ( .A1(n_207), .A2(n_237), .B1(n_382), .B2(n_391), .C(n_396), .Y(n_1099) );
INVx1_ASAP7_75t_L g1017 ( .A(n_208), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_209), .A2(n_240), .B1(n_516), .B2(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g937 ( .A(n_210), .Y(n_937) );
INVx1_ASAP7_75t_L g1339 ( .A(n_211), .Y(n_1339) );
CKINVDCx5p33_ASAP7_75t_R g1176 ( .A(n_212), .Y(n_1176) );
INVx1_ASAP7_75t_L g1227 ( .A(n_213), .Y(n_1227) );
INVx1_ASAP7_75t_L g1121 ( .A(n_214), .Y(n_1121) );
INVxp67_ASAP7_75t_SL g1305 ( .A(n_215), .Y(n_1305) );
INVx1_ASAP7_75t_L g1075 ( .A(n_216), .Y(n_1075) );
AOI221xp5_ASAP7_75t_L g1318 ( .A1(n_217), .A2(n_278), .B1(n_722), .B2(n_1138), .C(n_1319), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_217), .A2(n_273), .B1(n_771), .B2(n_1341), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_218), .A2(n_250), .B1(n_475), .B2(n_516), .C(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g1002 ( .A(n_219), .Y(n_1002) );
AOI22xp33_ASAP7_75t_SL g1025 ( .A1(n_219), .A2(n_266), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
CKINVDCx5p33_ASAP7_75t_R g1619 ( .A(n_220), .Y(n_1619) );
INVx1_ASAP7_75t_L g1388 ( .A(n_221), .Y(n_1388) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_222), .Y(n_318) );
OAI222xp33_ASAP7_75t_L g687 ( .A1(n_223), .A2(n_290), .B1(n_688), .B2(n_692), .C1(n_700), .C2(n_708), .Y(n_687) );
INVx1_ASAP7_75t_L g755 ( .A(n_223), .Y(n_755) );
INVx1_ASAP7_75t_L g1064 ( .A(n_224), .Y(n_1064) );
INVx1_ASAP7_75t_L g1110 ( .A(n_225), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_225), .A2(n_226), .B1(n_384), .B2(n_738), .Y(n_1134) );
INVx1_ASAP7_75t_L g1113 ( .A(n_226), .Y(n_1113) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_227), .Y(n_875) );
INVx1_ASAP7_75t_L g1367 ( .A(n_228), .Y(n_1367) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_229), .Y(n_524) );
XNOR2xp5_ASAP7_75t_L g1678 ( .A(n_231), .B(n_1679), .Y(n_1678) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_232), .Y(n_361) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_233), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_233), .A2(n_485), .B1(n_490), .B2(n_497), .Y(n_484) );
INVx1_ASAP7_75t_L g1300 ( .A(n_235), .Y(n_1300) );
INVx1_ASAP7_75t_L g1303 ( .A(n_236), .Y(n_1303) );
OAI221xp5_ASAP7_75t_L g1057 ( .A1(n_237), .A2(n_262), .B1(n_458), .B2(n_462), .C(n_469), .Y(n_1057) );
INVx1_ASAP7_75t_L g731 ( .A(n_238), .Y(n_731) );
INVx1_ASAP7_75t_L g1035 ( .A(n_239), .Y(n_1035) );
INVxp67_ASAP7_75t_SL g1283 ( .A(n_242), .Y(n_1283) );
OAI211xp5_ASAP7_75t_L g1111 ( .A1(n_244), .A2(n_428), .B(n_469), .C(n_1112), .Y(n_1111) );
INVxp33_ASAP7_75t_SL g1133 ( .A(n_244), .Y(n_1133) );
INVx1_ASAP7_75t_L g1359 ( .A(n_246), .Y(n_1359) );
INVx1_ASAP7_75t_L g1316 ( .A(n_247), .Y(n_1316) );
INVx1_ASAP7_75t_L g860 ( .A(n_248), .Y(n_860) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_249), .Y(n_344) );
INVx1_ASAP7_75t_L g1615 ( .A(n_252), .Y(n_1615) );
INVxp67_ASAP7_75t_SL g1620 ( .A(n_253), .Y(n_1620) );
OAI221xp5_ASAP7_75t_L g1634 ( .A1(n_253), .A2(n_469), .B1(n_990), .B2(n_1635), .C(n_1640), .Y(n_1634) );
INVx1_ASAP7_75t_L g995 ( .A(n_254), .Y(n_995) );
OAI21xp33_ASAP7_75t_L g1045 ( .A1(n_254), .A2(n_396), .B(n_914), .Y(n_1045) );
BUFx3_ASAP7_75t_L g322 ( .A(n_255), .Y(n_322) );
INVx1_ASAP7_75t_L g412 ( .A(n_255), .Y(n_412) );
INVx1_ASAP7_75t_L g1120 ( .A(n_257), .Y(n_1120) );
CKINVDCx5p33_ASAP7_75t_R g1258 ( .A(n_258), .Y(n_1258) );
INVx1_ASAP7_75t_L g975 ( .A(n_259), .Y(n_975) );
INVx1_ASAP7_75t_L g1224 ( .A(n_260), .Y(n_1224) );
OAI211xp5_ASAP7_75t_L g1259 ( .A1(n_260), .A2(n_1197), .B(n_1202), .C(n_1260), .Y(n_1259) );
AOI21xp5_ASAP7_75t_L g1632 ( .A1(n_261), .A2(n_834), .B(n_1191), .Y(n_1632) );
INVx1_ASAP7_75t_L g1650 ( .A(n_261), .Y(n_1650) );
INVxp67_ASAP7_75t_SL g1101 ( .A(n_262), .Y(n_1101) );
INVx1_ASAP7_75t_L g1639 ( .A(n_263), .Y(n_1639) );
OAI211xp5_ASAP7_75t_L g712 ( .A1(n_264), .A2(n_713), .B(n_715), .C(n_729), .Y(n_712) );
INVx1_ASAP7_75t_L g763 ( .A(n_264), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g1625 ( .A(n_265), .Y(n_1625) );
INVx1_ASAP7_75t_L g1010 ( .A(n_266), .Y(n_1010) );
INVx1_ASAP7_75t_L g421 ( .A(n_267), .Y(n_421) );
INVx2_ASAP7_75t_L g339 ( .A(n_269), .Y(n_339) );
INVx1_ASAP7_75t_L g380 ( .A(n_269), .Y(n_380) );
INVx1_ASAP7_75t_L g402 ( .A(n_269), .Y(n_402) );
XOR2x2_ASAP7_75t_L g570 ( .A(n_270), .B(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_271), .A2(n_283), .B1(n_475), .B2(n_477), .Y(n_1072) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_271), .Y(n_1097) );
INVx1_ASAP7_75t_L g1277 ( .A(n_272), .Y(n_1277) );
INVxp67_ASAP7_75t_SL g1379 ( .A(n_274), .Y(n_1379) );
INVx1_ASAP7_75t_L g511 ( .A(n_275), .Y(n_511) );
AOI21xp33_ASAP7_75t_L g1326 ( .A1(n_276), .A2(n_1137), .B(n_1173), .Y(n_1326) );
INVx1_ASAP7_75t_L g1333 ( .A(n_276), .Y(n_1333) );
INVx1_ASAP7_75t_L g534 ( .A(n_277), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g1630 ( .A(n_279), .Y(n_1630) );
INVx1_ASAP7_75t_L g1060 ( .A(n_280), .Y(n_1060) );
INVx1_ASAP7_75t_L g801 ( .A(n_282), .Y(n_801) );
INVxp67_ASAP7_75t_SL g1088 ( .A(n_283), .Y(n_1088) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_285), .Y(n_1211) );
NOR2xp33_ASAP7_75t_L g1661 ( .A(n_286), .B(n_1662), .Y(n_1661) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_287), .Y(n_892) );
OAI21xp33_ASAP7_75t_SL g1105 ( .A1(n_288), .A2(n_950), .B(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1109 ( .A(n_288), .Y(n_1109) );
INVx1_ASAP7_75t_L g601 ( .A(n_289), .Y(n_601) );
INVx1_ASAP7_75t_L g758 ( .A(n_290), .Y(n_758) );
INVx1_ASAP7_75t_L g634 ( .A(n_292), .Y(n_634) );
OAI211xp5_ASAP7_75t_L g658 ( .A1(n_292), .A2(n_600), .B(n_659), .C(n_662), .Y(n_658) );
INVxp67_ASAP7_75t_SL g790 ( .A(n_293), .Y(n_790) );
OAI221xp5_ASAP7_75t_L g942 ( .A1(n_294), .A2(n_296), .B1(n_528), .B2(n_888), .C(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g1627 ( .A(n_295), .Y(n_1627) );
INVxp67_ASAP7_75t_SL g955 ( .A(n_296), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_323), .B(n_1399), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx4f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_308), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g1670 ( .A(n_302), .B(n_311), .Y(n_1670) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g1676 ( .A(n_304), .B(n_307), .Y(n_1676) );
INVx1_ASAP7_75t_L g1684 ( .A(n_304), .Y(n_1684) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g1686 ( .A(n_307), .B(n_1684), .Y(n_1686) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g650 ( .A(n_311), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g377 ( .A(n_312), .B(n_322), .Y(n_377) );
AND2x4_ASAP7_75t_L g699 ( .A(n_312), .B(n_321), .Y(n_699) );
INVx1_ASAP7_75t_L g646 ( .A(n_313), .Y(n_646) );
AND2x4_ASAP7_75t_SL g1669 ( .A(n_313), .B(n_1670), .Y(n_1669) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x6_ASAP7_75t_L g314 ( .A(n_315), .B(n_320), .Y(n_314) );
BUFx4f_ASAP7_75t_L g343 ( .A(n_315), .Y(n_343) );
INVxp67_ASAP7_75t_L g372 ( .A(n_315), .Y(n_372) );
OR2x6_ASAP7_75t_L g640 ( .A(n_315), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g1302 ( .A(n_315), .Y(n_1302) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g608 ( .A(n_316), .Y(n_608) );
BUFx4f_ASAP7_75t_L g964 ( .A(n_316), .Y(n_964) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g349 ( .A(n_318), .Y(n_349) );
NAND2x1_ASAP7_75t_L g355 ( .A(n_318), .B(n_319), .Y(n_355) );
INVx2_ASAP7_75t_L g360 ( .A(n_318), .Y(n_360) );
INVx1_ASAP7_75t_L g394 ( .A(n_318), .Y(n_394) );
AND2x2_ASAP7_75t_L g507 ( .A(n_318), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g629 ( .A(n_318), .B(n_319), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_319), .B(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g359 ( .A(n_319), .B(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g390 ( .A(n_319), .Y(n_390) );
INVx1_ASAP7_75t_L g406 ( .A(n_319), .Y(n_406) );
AND2x2_ASAP7_75t_L g415 ( .A(n_319), .B(n_349), .Y(n_415) );
INVx2_ASAP7_75t_L g508 ( .A(n_319), .Y(n_508) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g627 ( .A(n_321), .Y(n_627) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g633 ( .A(n_322), .Y(n_633) );
AND2x4_ASAP7_75t_L g637 ( .A(n_322), .B(n_393), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B1(n_980), .B2(n_981), .Y(n_323) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B1(n_786), .B2(n_979), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_568), .B1(n_569), .B2(n_785), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g785 ( .A(n_329), .Y(n_785) );
XNOR2x1_ASAP7_75t_L g329 ( .A(n_330), .B(n_509), .Y(n_329) );
XNOR2x1_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NOR2x1_ASAP7_75t_L g332 ( .A(n_333), .B(n_425), .Y(n_332) );
NAND3xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_398), .C(n_420), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_381), .Y(n_334) );
OAI33xp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_341), .A3(n_350), .B1(n_362), .B2(n_370), .B3(n_375), .Y(n_335) );
OAI22xp5_ASAP7_75t_SL g552 ( .A1(n_336), .A2(n_553), .B1(n_558), .B2(n_561), .Y(n_552) );
OAI33xp33_ASAP7_75t_L g1086 ( .A1(n_336), .A2(n_1087), .A3(n_1092), .B1(n_1094), .B2(n_1096), .B3(n_1098), .Y(n_1086) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g603 ( .A(n_337), .Y(n_603) );
AOI31xp33_ASAP7_75t_L g803 ( .A1(n_337), .A2(n_567), .A3(n_804), .B(n_806), .Y(n_803) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_337), .Y(n_900) );
INVx2_ASAP7_75t_L g973 ( .A(n_337), .Y(n_973) );
INVx4_ASAP7_75t_L g1141 ( .A(n_337), .Y(n_1141) );
AOI222xp33_ASAP7_75t_L g1288 ( .A1(n_337), .A2(n_399), .B1(n_818), .B2(n_1289), .C1(n_1290), .C2(n_1298), .Y(n_1288) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx1_ASAP7_75t_L g501 ( .A(n_338), .Y(n_501) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_339), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g544 ( .A(n_339), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_344), .B2(n_345), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g485 ( .A1(n_344), .A2(n_369), .B1(n_479), .B2(n_486), .C(n_487), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_345), .A2(n_371), .B1(n_373), .B2(n_374), .Y(n_370) );
HB1xp67_ASAP7_75t_L g1036 ( .A(n_345), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_345), .A2(n_1300), .B1(n_1301), .B2(n_1303), .Y(n_1299) );
OAI22xp5_ASAP7_75t_L g1395 ( .A1(n_345), .A2(n_1369), .B1(n_1396), .B2(n_1397), .Y(n_1395) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx4_ASAP7_75t_L g610 ( .A(n_346), .Y(n_610) );
INVx2_ASAP7_75t_L g706 ( .A(n_346), .Y(n_706) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_346), .Y(n_909) );
INVx1_ASAP7_75t_L g1170 ( .A(n_346), .Y(n_1170) );
INVx2_ASAP7_75t_L g1391 ( .A(n_346), .Y(n_1391) );
INVx8_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g644 ( .A(n_347), .B(n_633), .Y(n_644) );
BUFx2_ASAP7_75t_L g1091 ( .A(n_347), .Y(n_1091) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_356), .B2(n_361), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_351), .A2(n_374), .B1(n_491), .B2(n_493), .Y(n_490) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_352), .Y(n_613) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g969 ( .A(n_353), .Y(n_969) );
INVx1_ASAP7_75t_L g1394 ( .A(n_353), .Y(n_1394) );
INVx4_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x6_ASAP7_75t_L g396 ( .A(n_354), .B(n_397), .Y(n_396) );
BUFx4f_ASAP7_75t_L g555 ( .A(n_354), .Y(n_555) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_354), .Y(n_563) );
BUFx4f_ASAP7_75t_L g617 ( .A(n_354), .Y(n_617) );
BUFx4f_ASAP7_75t_L g1325 ( .A(n_354), .Y(n_1325) );
BUFx4f_ASAP7_75t_L g1387 ( .A(n_354), .Y(n_1387) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx3_ASAP7_75t_L g368 ( .A(n_355), .Y(n_368) );
INVx4_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g1386 ( .A(n_357), .Y(n_1386) );
INVx2_ASAP7_75t_L g1656 ( .A(n_357), .Y(n_1656) );
INVx4_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g365 ( .A(n_359), .Y(n_365) );
BUFx3_ASAP7_75t_L g554 ( .A(n_359), .Y(n_554) );
INVx1_ASAP7_75t_L g907 ( .A(n_359), .Y(n_907) );
BUFx2_ASAP7_75t_L g1095 ( .A(n_359), .Y(n_1095) );
AND2x2_ASAP7_75t_L g405 ( .A(n_360), .B(n_406), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g478 ( .A1(n_361), .A2(n_366), .B1(n_479), .B2(n_480), .C(n_482), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B1(n_367), .B2(n_369), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g1392 ( .A1(n_363), .A2(n_1373), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
INVx4_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g562 ( .A(n_365), .Y(n_562) );
INVx2_ASAP7_75t_L g612 ( .A(n_365), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_367), .A2(n_607), .B1(n_872), .B2(n_883), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_367), .A2(n_906), .B1(n_1064), .B2(n_1093), .Y(n_1092) );
BUFx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g418 ( .A(n_368), .B(n_410), .Y(n_418) );
INVx2_ASAP7_75t_SL g694 ( .A(n_368), .Y(n_694) );
OR2x2_ASAP7_75t_L g914 ( .A(n_368), .B(n_410), .Y(n_914) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI33xp33_ASAP7_75t_L g1384 ( .A1(n_375), .A2(n_603), .A3(n_1385), .B1(n_1389), .B2(n_1392), .B3(n_1395), .Y(n_1384) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g1098 ( .A(n_376), .Y(n_1098) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_377), .B(n_378), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_377), .B(n_559), .Y(n_558) );
INVx4_ASAP7_75t_L g722 ( .A(n_377), .Y(n_722) );
AND2x4_ASAP7_75t_L g818 ( .A(n_377), .B(n_559), .Y(n_818) );
INVx4_ASAP7_75t_L g1156 ( .A(n_377), .Y(n_1156) );
INVx1_ASAP7_75t_L g560 ( .A(n_378), .Y(n_560) );
OR2x2_ASAP7_75t_L g575 ( .A(n_378), .B(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_378), .Y(n_683) );
OR2x2_ASAP7_75t_L g740 ( .A(n_378), .B(n_456), .Y(n_740) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx2_ASAP7_75t_L g395 ( .A(n_379), .Y(n_395) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g810 ( .A(n_384), .Y(n_810) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_384), .Y(n_1047) );
NAND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g397 ( .A(n_385), .Y(n_397) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_387), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_387), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g711 ( .A(n_387), .Y(n_711) );
AND2x6_ASAP7_75t_L g728 ( .A(n_387), .B(n_628), .Y(n_728) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_387), .B(n_1220), .Y(n_1219) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g632 ( .A(n_390), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g710 ( .A(n_390), .Y(n_710) );
BUFx2_ASAP7_75t_L g1220 ( .A(n_390), .Y(n_1220) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_395), .Y(n_391) );
OR2x2_ASAP7_75t_L g738 ( .A(n_392), .B(n_395), .Y(n_738) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g423 ( .A(n_395), .Y(n_423) );
INVx1_ASAP7_75t_L g651 ( .A(n_395), .Y(n_651) );
INVxp67_ASAP7_75t_L g766 ( .A(n_395), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_396), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g903 ( .A1(n_396), .A2(n_904), .B(n_905), .Y(n_903) );
OAI21xp5_ASAP7_75t_L g966 ( .A1(n_396), .A2(n_967), .B(n_972), .Y(n_966) );
OAI21xp5_ASAP7_75t_SL g1646 ( .A1(n_396), .A2(n_1647), .B(n_1649), .Y(n_1646) );
AOI222xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_407), .B1(n_408), .B2(n_416), .C1(n_417), .C2(n_419), .Y(n_398) );
AOI322xp5_ASAP7_75t_L g1020 ( .A1(n_399), .A2(n_818), .A3(n_1021), .B1(n_1025), .B2(n_1029), .C1(n_1030), .C2(n_1037), .Y(n_1020) );
AOI222xp33_ASAP7_75t_L g1100 ( .A1(n_399), .A2(n_408), .B1(n_417), .B2(n_1056), .C1(n_1076), .C2(n_1101), .Y(n_1100) );
AOI332xp33_ASAP7_75t_L g1135 ( .A1(n_399), .A2(n_818), .A3(n_1136), .B1(n_1139), .B2(n_1140), .B3(n_1142), .C1(n_1143), .C2(n_1145), .Y(n_1135) );
AOI222xp33_ASAP7_75t_L g1377 ( .A1(n_399), .A2(n_408), .B1(n_417), .B2(n_1359), .C1(n_1378), .C2(n_1379), .Y(n_1377) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_403), .Y(n_399) );
AOI332xp33_ASAP7_75t_L g548 ( .A1(n_400), .A2(n_403), .A3(n_409), .B1(n_413), .B2(n_417), .B3(n_534), .C1(n_549), .C2(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g751 ( .A(n_401), .B(n_404), .Y(n_751) );
AND2x4_ASAP7_75t_L g757 ( .A(n_401), .B(n_435), .Y(n_757) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_402), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g597 ( .A(n_402), .Y(n_597) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g424 ( .A(n_405), .B(n_411), .Y(n_424) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_405), .Y(n_557) );
INVx3_ASAP7_75t_L g725 ( .A(n_405), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_408), .A2(n_417), .B1(n_800), .B2(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g913 ( .A(n_408), .Y(n_913) );
INVxp67_ASAP7_75t_L g953 ( .A(n_408), .Y(n_953) );
AOI211xp5_ASAP7_75t_L g1043 ( .A1(n_408), .A2(n_1044), .B(n_1045), .C(n_1046), .Y(n_1043) );
AOI21xp33_ASAP7_75t_L g1132 ( .A1(n_408), .A2(n_1133), .B(n_1134), .Y(n_1132) );
AOI222xp33_ASAP7_75t_L g1285 ( .A1(n_408), .A2(n_810), .B1(n_812), .B2(n_1279), .C1(n_1286), .C2(n_1287), .Y(n_1285) );
INVx1_ASAP7_75t_L g1618 ( .A(n_408), .Y(n_1618) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_413), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g505 ( .A(n_411), .B(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_SL g691 ( .A(n_411), .B(n_628), .Y(n_691) );
AND2x4_ASAP7_75t_L g714 ( .A(n_411), .B(n_565), .Y(n_714) );
AND2x4_ASAP7_75t_L g733 ( .A(n_411), .B(n_506), .Y(n_733) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_411), .B(n_413), .Y(n_1313) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_412), .Y(n_641) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g1329 ( .A(n_414), .Y(n_1329) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_415), .Y(n_565) );
BUFx3_ASAP7_75t_L g727 ( .A(n_415), .Y(n_727) );
BUFx3_ASAP7_75t_L g808 ( .A(n_415), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_416), .A2(n_427), .B1(n_440), .B2(n_453), .C(n_457), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g1129 ( .A1(n_417), .A2(n_567), .B(n_1114), .Y(n_1129) );
AOI21xp5_ASAP7_75t_L g1306 ( .A1(n_417), .A2(n_567), .B(n_1307), .Y(n_1306) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_422), .B(n_539), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_422), .B(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g915 ( .A1(n_422), .A2(n_504), .B1(n_916), .B2(n_917), .Y(n_915) );
INVx3_ASAP7_75t_L g950 ( .A(n_422), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_422), .B(n_1305), .Y(n_1304) );
AOI222xp33_ASAP7_75t_L g1614 ( .A1(n_422), .A2(n_504), .B1(n_1615), .B2(n_1616), .C1(n_1619), .C2(n_1620), .Y(n_1614) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
AND2x4_ASAP7_75t_L g504 ( .A(n_423), .B(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_424), .Y(n_730) );
INVx1_ASAP7_75t_L g1223 ( .A(n_424), .Y(n_1223) );
A2O1A1Ixp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_467), .B(n_499), .C(n_502), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g533 ( .A1(n_427), .A2(n_453), .B1(n_534), .B2(n_535), .C(n_541), .Y(n_533) );
INVx2_ASAP7_75t_L g846 ( .A(n_427), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_427), .A2(n_940), .B1(n_942), .B2(n_948), .Y(n_939) );
AOI211xp5_ASAP7_75t_L g1055 ( .A1(n_427), .A2(n_1056), .B(n_1057), .C(n_1058), .Y(n_1055) );
AOI211xp5_ASAP7_75t_SL g1278 ( .A1(n_427), .A2(n_1279), .B(n_1280), .C(n_1281), .Y(n_1278) );
AOI211xp5_ASAP7_75t_L g1358 ( .A1(n_427), .A2(n_1359), .B(n_1360), .C(n_1361), .Y(n_1358) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x6_ASAP7_75t_L g765 ( .A(n_428), .B(n_766), .Y(n_765) );
OR2x2_ASAP7_75t_L g1617 ( .A(n_428), .B(n_766), .Y(n_1617) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_429), .B(n_435), .Y(n_428) );
BUFx3_ASAP7_75t_L g475 ( .A(n_429), .Y(n_475) );
BUFx3_ASAP7_75t_L g540 ( .A(n_429), .Y(n_540) );
INVx8_ASAP7_75t_L g744 ( .A(n_429), .Y(n_744) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_429), .B(n_1016), .Y(n_1015) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
AND2x4_ASAP7_75t_L g451 ( .A(n_430), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g442 ( .A(n_431), .B(n_433), .Y(n_442) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_431), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_431), .B(n_448), .Y(n_496) );
AND2x4_ASAP7_75t_L g661 ( .A(n_431), .B(n_466), .Y(n_661) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g452 ( .A(n_434), .Y(n_452) );
AND2x6_ASAP7_75t_L g459 ( .A(n_435), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g463 ( .A(n_435), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g471 ( .A(n_435), .Y(n_471) );
AND2x4_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g488 ( .A(n_436), .B(n_489), .Y(n_488) );
NAND3x1_ASAP7_75t_L g596 ( .A(n_436), .B(n_489), .C(n_597), .Y(n_596) );
OR2x4_ASAP7_75t_L g654 ( .A(n_436), .B(n_442), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_436), .Y(n_657) );
AND2x4_ASAP7_75t_L g660 ( .A(n_436), .B(n_661), .Y(n_660) );
OR2x6_ASAP7_75t_L g676 ( .A(n_436), .B(n_677), .Y(n_676) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g483 ( .A(n_437), .Y(n_483) );
NAND2xp33_ASAP7_75t_SL g576 ( .A(n_437), .B(n_439), .Y(n_576) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g482 ( .A(n_439), .B(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_439), .Y(n_681) );
AND3x4_ASAP7_75t_L g769 ( .A(n_439), .B(n_483), .C(n_544), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g877 ( .A1(n_441), .A2(n_487), .B1(n_878), .B2(n_879), .C(n_881), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_441), .A2(n_1367), .B1(n_1368), .B2(n_1369), .Y(n_1366) );
BUFx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx3_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
BUFx4f_ASAP7_75t_L g525 ( .A(n_442), .Y(n_525) );
OR2x4_ASAP7_75t_L g674 ( .A(n_442), .B(n_657), .Y(n_674) );
INVx2_ASAP7_75t_L g886 ( .A(n_442), .Y(n_886) );
OAI22xp33_ASAP7_75t_L g1245 ( .A1(n_443), .A2(n_579), .B1(n_1246), .B2(n_1247), .Y(n_1245) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g537 ( .A(n_444), .Y(n_537) );
INVx3_ASAP7_75t_L g1070 ( .A(n_444), .Y(n_1070) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_445), .A2(n_482), .B1(n_518), .B2(n_519), .C(n_520), .Y(n_517) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_445), .Y(n_582) );
OR2x2_ASAP7_75t_L g739 ( .A(n_445), .B(n_740), .Y(n_739) );
INVx4_ASAP7_75t_L g880 ( .A(n_445), .Y(n_880) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g470 ( .A(n_446), .Y(n_470) );
BUFx3_ASAP7_75t_L g479 ( .A(n_446), .Y(n_479) );
NAND2x1p5_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
BUFx2_ASAP7_75t_L g669 ( .A(n_447), .Y(n_669) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g466 ( .A(n_448), .Y(n_466) );
INVx2_ASAP7_75t_L g461 ( .A(n_449), .Y(n_461) );
AND2x4_ASAP7_75t_L g477 ( .A(n_449), .B(n_465), .Y(n_477) );
BUFx2_ASAP7_75t_L g666 ( .A(n_449), .Y(n_666) );
INVx3_ASAP7_75t_L g481 ( .A(n_450), .Y(n_481) );
BUFx2_ASAP7_75t_L g588 ( .A(n_450), .Y(n_588) );
OR2x6_ASAP7_75t_SL g990 ( .A(n_450), .B(n_991), .Y(n_990) );
BUFx2_ASAP7_75t_L g1188 ( .A(n_450), .Y(n_1188) );
INVx1_ASAP7_75t_L g1242 ( .A(n_450), .Y(n_1242) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx8_ASAP7_75t_L g492 ( .A(n_451), .Y(n_492) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_451), .Y(n_521) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_451), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_453), .A2(n_800), .B1(n_841), .B2(n_845), .Y(n_840) );
INVx1_ASAP7_75t_L g858 ( .A(n_453), .Y(n_858) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g941 ( .A(n_454), .Y(n_941) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g498 ( .A(n_455), .B(n_477), .Y(n_498) );
INVx2_ASAP7_75t_L g991 ( .A(n_455), .Y(n_991) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g1016 ( .A(n_456), .Y(n_1016) );
INVx4_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_459), .A2(n_463), .B1(n_468), .B2(n_937), .C(n_938), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_459), .A2(n_463), .B1(n_994), .B2(n_995), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_459), .A2(n_463), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1626 ( .A1(n_459), .A2(n_463), .B1(n_1627), .B2(n_1628), .Y(n_1626) );
AND2x2_ASAP7_75t_L g756 ( .A(n_460), .B(n_757), .Y(n_756) );
NAND2x1_ASAP7_75t_L g1262 ( .A(n_460), .B(n_757), .Y(n_1262) );
AND2x4_ASAP7_75t_SL g1345 ( .A(n_460), .B(n_757), .Y(n_1345) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_463), .Y(n_829) );
INVx1_ASAP7_75t_L g761 ( .A(n_464), .Y(n_761) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_472), .C(n_484), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_468), .B(n_515), .C(n_522), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_468), .B(n_827), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_470), .A2(n_487), .B1(n_524), .B2(n_525), .C(n_526), .Y(n_523) );
INVx1_ASAP7_75t_L g869 ( .A(n_471), .Y(n_869) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g935 ( .A(n_475), .Y(n_935) );
AOI221xp5_ASAP7_75t_SL g859 ( .A1(n_476), .A2(n_860), .B1(n_861), .B2(n_863), .C(n_864), .Y(n_859) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx12f_ASAP7_75t_L g516 ( .A(n_477), .Y(n_516) );
BUFx3_ASAP7_75t_L g777 ( .A(n_477), .Y(n_777) );
BUFx2_ASAP7_75t_L g927 ( .A(n_477), .Y(n_927) );
INVx5_ASAP7_75t_L g1193 ( .A(n_477), .Y(n_1193) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_479), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g1270 ( .A1(n_479), .A2(n_482), .B1(n_865), .B2(n_1271), .C(n_1272), .Y(n_1270) );
OAI221xp5_ASAP7_75t_L g1275 ( .A1(n_479), .A2(n_487), .B1(n_525), .B2(n_1276), .C(n_1277), .Y(n_1275) );
OAI221xp5_ASAP7_75t_L g1372 ( .A1(n_479), .A2(n_486), .B1(n_487), .B2(n_1373), .C(n_1374), .Y(n_1372) );
INVx2_ASAP7_75t_L g1637 ( .A(n_479), .Y(n_1637) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g536 ( .A(n_481), .Y(n_536) );
OAI221xp5_ASAP7_75t_L g891 ( .A1(n_482), .A2(n_892), .B1(n_893), .B2(n_894), .C(n_896), .Y(n_891) );
OAI221xp5_ASAP7_75t_L g1116 ( .A1(n_482), .A2(n_582), .B1(n_839), .B2(n_1117), .C(n_1118), .Y(n_1116) );
OAI21xp33_ASAP7_75t_L g1364 ( .A1(n_482), .A2(n_839), .B(n_1365), .Y(n_1364) );
INVx3_ASAP7_75t_L g665 ( .A(n_483), .Y(n_665) );
OAI221xp5_ASAP7_75t_L g1122 ( .A1(n_486), .A2(n_487), .B1(n_893), .B2(n_1123), .C(n_1124), .Y(n_1122) );
INVx3_ASAP7_75t_L g836 ( .A(n_487), .Y(n_836) );
OAI221xp5_ASAP7_75t_L g1635 ( .A1(n_487), .A2(n_579), .B1(n_1636), .B2(n_1638), .C(n_1639), .Y(n_1635) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g1191 ( .A(n_491), .Y(n_1191) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g746 ( .A(n_492), .B(n_745), .Y(n_746) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_492), .Y(n_779) );
INVx3_ASAP7_75t_L g839 ( .A(n_492), .Y(n_839) );
INVx2_ASAP7_75t_SL g1063 ( .A(n_492), .Y(n_1063) );
INVx2_ASAP7_75t_SL g1641 ( .A(n_492), .Y(n_1641) );
OAI22xp5_ASAP7_75t_L g1119 ( .A1(n_493), .A2(n_885), .B1(n_1120), .B2(n_1121), .Y(n_1119) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g531 ( .A(n_494), .Y(n_531) );
CKINVDCx8_ASAP7_75t_R g843 ( .A(n_494), .Y(n_843) );
INVx1_ASAP7_75t_L g1368 ( .A(n_494), .Y(n_1368) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g591 ( .A(n_495), .Y(n_591) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx2_ASAP7_75t_L g677 ( .A(n_496), .Y(n_677) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g1073 ( .A1(n_498), .A2(n_1074), .B1(n_1075), .B2(n_1076), .C(n_1077), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_498), .B(n_501), .Y(n_1664) );
A2O1A1Ixp33_ASAP7_75t_L g1266 ( .A1(n_499), .A2(n_1267), .B(n_1278), .C(n_1282), .Y(n_1266) );
INVx1_ASAP7_75t_L g1375 ( .A(n_499), .Y(n_1375) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g921 ( .A1(n_500), .A2(n_922), .B(n_949), .Y(n_921) );
OAI31xp33_ASAP7_75t_SL g988 ( .A1(n_500), .A2(n_989), .A3(n_992), .B(n_996), .Y(n_988) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g898 ( .A(n_501), .Y(n_898) );
NAND2xp33_ASAP7_75t_SL g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g547 ( .A(n_504), .Y(n_547) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_504), .Y(n_956) );
INVx1_ASAP7_75t_L g1041 ( .A(n_504), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_504), .B(n_1075), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_504), .B(n_1131), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1380 ( .A(n_504), .B(n_1381), .Y(n_1380) );
BUFx6f_ASAP7_75t_L g1137 ( .A(n_506), .Y(n_1137) );
INVx2_ASAP7_75t_L g1217 ( .A(n_506), .Y(n_1217) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g648 ( .A(n_507), .B(n_641), .Y(n_648) );
INVx2_ASAP7_75t_L g721 ( .A(n_507), .Y(n_721) );
BUFx3_ASAP7_75t_L g1154 ( .A(n_507), .Y(n_1154) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
XNOR2x1_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_546), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_533), .B(n_542), .C(n_545), .Y(n_513) );
BUFx2_ASAP7_75t_L g1189 ( .A(n_516), .Y(n_1189) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_518), .A2(n_524), .B1(n_562), .B2(n_563), .C(n_564), .Y(n_561) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_519), .A2(n_530), .B1(n_554), .B2(n_555), .C(n_556), .Y(n_553) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g585 ( .A(n_521), .Y(n_585) );
AND2x4_ASAP7_75t_L g656 ( .A(n_521), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g842 ( .A(n_521), .Y(n_842) );
BUFx6f_ASAP7_75t_L g895 ( .A(n_521), .Y(n_895) );
BUFx6f_ASAP7_75t_L g1008 ( .A(n_521), .Y(n_1008) );
INVx1_ASAP7_75t_L g580 ( .A(n_525), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_530), .B1(n_531), .B2(n_532), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx5_ASAP7_75t_L g776 ( .A(n_529), .Y(n_776) );
INVx2_ASAP7_75t_SL g865 ( .A(n_529), .Y(n_865) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_529), .Y(n_874) );
INVx2_ASAP7_75t_SL g933 ( .A(n_529), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_531), .A2(n_584), .B1(n_585), .B2(n_586), .Y(n_583) );
HB1xp67_ASAP7_75t_L g1631 ( .A(n_537), .Y(n_1631) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx2_ASAP7_75t_SL g926 ( .A(n_540), .Y(n_926) );
BUFx3_ASAP7_75t_L g1012 ( .A(n_540), .Y(n_1012) );
OAI21xp33_ASAP7_75t_L g1310 ( .A1(n_542), .A2(n_1311), .B(n_1321), .Y(n_1310) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g1080 ( .A(n_543), .Y(n_1080) );
BUFx2_ASAP7_75t_L g1174 ( .A(n_543), .Y(n_1174) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g735 ( .A(n_544), .Y(n_735) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_544), .A2(n_825), .B1(n_847), .B2(n_848), .Y(n_824) );
OAI31xp33_ASAP7_75t_SL g1106 ( .A1(n_544), .A2(n_1107), .A3(n_1111), .B(n_1115), .Y(n_1106) );
INVx1_ASAP7_75t_L g847 ( .A(n_547), .Y(n_847) );
NOR3xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_566), .C(n_567), .Y(n_551) );
INVx2_ASAP7_75t_L g616 ( .A(n_554), .Y(n_616) );
OAI221xp5_ASAP7_75t_L g1649 ( .A1(n_555), .A2(n_612), .B1(n_1642), .B2(n_1650), .C(n_1651), .Y(n_1649) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_557), .Y(n_807) );
INVx3_ASAP7_75t_L g1659 ( .A(n_557), .Y(n_1659) );
INVx1_ASAP7_75t_L g619 ( .A(n_558), .Y(n_619) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI221xp5_ASAP7_75t_L g692 ( .A1(n_562), .A2(n_693), .B1(n_695), .B2(n_696), .C(n_697), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_563), .A2(n_1060), .B1(n_1069), .B2(n_1095), .Y(n_1094) );
INVx1_ASAP7_75t_L g817 ( .A(n_565), .Y(n_817) );
BUFx2_ASAP7_75t_L g1653 ( .A(n_565), .Y(n_1653) );
OR3x1_ASAP7_75t_L g1382 ( .A(n_567), .B(n_1383), .C(n_1384), .Y(n_1382) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
XNOR2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_684), .Y(n_569) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_623), .C(n_652), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_602), .Y(n_572) );
OAI33xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_577), .A3(n_583), .B1(n_587), .B2(n_593), .B3(n_598), .Y(n_573) );
BUFx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx8_ASAP7_75t_L g1244 ( .A(n_575), .Y(n_1244) );
BUFx2_ASAP7_75t_L g834 ( .A(n_576), .Y(n_834) );
OAI22xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B1(n_581), .B2(n_582), .Y(n_577) );
OAI22xp5_ASAP7_75t_SL g604 ( .A1(n_578), .A2(n_599), .B1(n_605), .B2(n_609), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_579), .A2(n_599), .B1(n_600), .B2(n_601), .Y(n_598) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_581), .A2(n_601), .B1(n_615), .B2(n_617), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_584), .A2(n_589), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g1005 ( .A(n_585), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_586), .A2(n_592), .B1(n_605), .B2(n_621), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_590), .B2(n_592), .Y(n_587) );
OAI221xp5_ASAP7_75t_L g997 ( .A1(n_590), .A2(n_998), .B1(n_1001), .B2(n_1002), .C(n_1003), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g1006 ( .A1(n_590), .A2(n_1007), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1239 ( .A1(n_590), .A2(n_1240), .B1(n_1241), .B2(n_1243), .Y(n_1239) );
BUFx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g750 ( .A(n_591), .B(n_740), .Y(n_750) );
INVx1_ASAP7_75t_L g1066 ( .A(n_591), .Y(n_1066) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI33xp33_ASAP7_75t_L g767 ( .A1(n_594), .A2(n_768), .A3(n_770), .B1(n_774), .B2(n_778), .B3(n_780), .Y(n_767) );
BUFx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g1254 ( .A(n_595), .Y(n_1254) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx3_ASAP7_75t_L g1194 ( .A(n_596), .Y(n_1194) );
OAI33xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .A3(n_611), .B1(n_614), .B2(n_618), .B3(n_620), .Y(n_602) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_SL g703 ( .A(n_608), .Y(n_703) );
BUFx6f_ASAP7_75t_L g1089 ( .A(n_608), .Y(n_1089) );
BUFx3_ASAP7_75t_L g1396 ( .A(n_608), .Y(n_1396) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g622 ( .A(n_610), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g1295 ( .A1(n_610), .A2(n_1277), .B1(n_1296), .B2(n_1297), .Y(n_1295) );
OAI221xp5_ASAP7_75t_L g967 ( .A1(n_615), .A2(n_968), .B1(n_969), .B2(n_970), .C(n_971), .Y(n_967) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g1655 ( .A1(n_617), .A2(n_1630), .B1(n_1638), .B2(n_1656), .C(n_1657), .Y(n_1655) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI31xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_638), .A3(n_645), .B(n_649), .Y(n_623) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
BUFx3_ASAP7_75t_L g717 ( .A(n_628), .Y(n_717) );
BUFx3_ASAP7_75t_L g805 ( .A(n_628), .Y(n_805) );
BUFx3_ASAP7_75t_L g960 ( .A(n_628), .Y(n_960) );
BUFx6f_ASAP7_75t_L g1024 ( .A(n_628), .Y(n_1024) );
BUFx3_ASAP7_75t_L g1138 ( .A(n_628), .Y(n_1138) );
INVx1_ASAP7_75t_L g1292 ( .A(n_628), .Y(n_1292) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g823 ( .A(n_629), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_634), .B2(n_635), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_631), .A2(n_663), .B1(n_667), .B2(n_670), .Y(n_662) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx3_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
BUFx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI31xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_658), .A3(n_671), .B(n_678), .Y(n_652) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
CKINVDCx8_ASAP7_75t_R g659 ( .A(n_660), .Y(n_659) );
BUFx2_ASAP7_75t_L g773 ( .A(n_661), .Y(n_773) );
BUFx2_ASAP7_75t_L g782 ( .A(n_661), .Y(n_782) );
BUFx3_ASAP7_75t_L g833 ( .A(n_661), .Y(n_833) );
INVx2_ASAP7_75t_L g862 ( .A(n_661), .Y(n_862) );
BUFx2_ASAP7_75t_L g929 ( .A(n_661), .Y(n_929) );
BUFx2_ASAP7_75t_L g947 ( .A(n_661), .Y(n_947) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_661), .B(n_1016), .Y(n_1018) );
BUFx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
AND2x4_ASAP7_75t_L g668 ( .A(n_665), .B(n_669), .Y(n_668) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
BUFx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
BUFx3_ASAP7_75t_L g876 ( .A(n_677), .Y(n_876) );
INVx1_ASAP7_75t_L g890 ( .A(n_677), .Y(n_890) );
BUFx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_680), .B(n_682), .Y(n_679) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND3x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_747), .C(n_753), .Y(n_685) );
O2A1O1Ixp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_712), .B(n_735), .C(n_736), .Y(n_686) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g1322 ( .A(n_689), .Y(n_1322) );
INVx4_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx3_ASAP7_75t_L g1226 ( .A(n_691), .Y(n_1226) );
INVx5_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g1173 ( .A(n_699), .Y(n_1173) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B1(n_704), .B2(n_707), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_702), .A2(n_1067), .B1(n_1091), .B2(n_1097), .Y(n_1096) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g1167 ( .A(n_709), .Y(n_1167) );
NOR2x1_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx3_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_SL g1233 ( .A1(n_714), .A2(n_732), .B1(n_1234), .B2(n_1235), .Y(n_1233) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_723), .B(n_728), .Y(n_715) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g820 ( .A(n_719), .Y(n_820) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
HB1xp67_ASAP7_75t_L g1031 ( .A(n_720), .Y(n_1031) );
INVx1_ASAP7_75t_L g1230 ( .A(n_720), .Y(n_1230) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g959 ( .A(n_721), .Y(n_959) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g1026 ( .A(n_725), .Y(n_1026) );
INVx2_ASAP7_75t_SL g1144 ( .A(n_725), .Y(n_1144) );
INVx1_ASAP7_75t_L g1328 ( .A(n_725), .Y(n_1328) );
INVx2_ASAP7_75t_L g1652 ( .A(n_725), .Y(n_1652) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g1028 ( .A(n_727), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g1232 ( .A(n_727), .Y(n_1232) );
AOI21xp5_ASAP7_75t_L g1151 ( .A1(n_728), .A2(n_1152), .B(n_1157), .Y(n_1151) );
AOI221xp5_ASAP7_75t_L g1225 ( .A1(n_728), .A2(n_1226), .B1(n_1227), .B2(n_1228), .C(n_1231), .Y(n_1225) );
AOI21xp5_ASAP7_75t_L g1317 ( .A1(n_728), .A2(n_1318), .B(n_1320), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_732), .B2(n_734), .Y(n_729) );
HB1xp67_ASAP7_75t_L g1161 ( .A(n_730), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_730), .A2(n_733), .B1(n_1315), .B2(n_1316), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_731), .A2(n_734), .B1(n_742), .B2(n_746), .Y(n_741) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g1164 ( .A(n_733), .Y(n_1164) );
INVx2_ASAP7_75t_L g1210 ( .A(n_737), .Y(n_1210) );
AND2x4_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx2_ASAP7_75t_SL g812 ( .A(n_738), .Y(n_812) );
AND2x4_ASAP7_75t_L g1351 ( .A(n_738), .B(n_739), .Y(n_1351) );
INVx1_ASAP7_75t_L g745 ( .A(n_740), .Y(n_745) );
INVx1_ASAP7_75t_L g1199 ( .A(n_740), .Y(n_1199) );
AND2x4_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .Y(n_742) );
AND2x4_ASAP7_75t_L g1353 ( .A(n_743), .B(n_745), .Y(n_1353) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx8_ASAP7_75t_L g771 ( .A(n_744), .Y(n_771) );
INVx3_ASAP7_75t_L g781 ( .A(n_744), .Y(n_781) );
INVx2_ASAP7_75t_L g945 ( .A(n_744), .Y(n_945) );
INVx2_ASAP7_75t_L g1200 ( .A(n_746), .Y(n_1200) );
INVx2_ASAP7_75t_L g1255 ( .A(n_746), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_746), .A2(n_1315), .B1(n_1316), .B2(n_1353), .Y(n_1352) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_752), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g1175 ( .A1(n_748), .A2(n_1176), .B(n_1177), .Y(n_1175) );
AOI221xp5_ASAP7_75t_L g1256 ( .A1(n_748), .A2(n_1235), .B1(n_1257), .B2(n_1258), .C(n_1259), .Y(n_1256) );
AOI21xp5_ASAP7_75t_L g1348 ( .A1(n_748), .A2(n_1349), .B(n_1350), .Y(n_1348) );
INVx8_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g798 ( .A(n_751), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g1663 ( .A(n_751), .B(n_1664), .Y(n_1663) );
AND4x1_ASAP7_75t_SL g753 ( .A(n_754), .B(n_762), .C(n_767), .D(n_783), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_758), .B2(n_759), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_756), .A2(n_759), .B1(n_1181), .B2(n_1182), .Y(n_1180) );
AND2x4_ASAP7_75t_L g759 ( .A(n_757), .B(n_760), .Y(n_759) );
AND2x4_ASAP7_75t_L g784 ( .A(n_757), .B(n_773), .Y(n_784) );
AND2x4_ASAP7_75t_SL g1347 ( .A(n_757), .B(n_760), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_759), .A2(n_1221), .B1(n_1227), .B2(n_1261), .Y(n_1260) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx5_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx3_ASAP7_75t_L g1257 ( .A(n_765), .Y(n_1257) );
AOI33xp33_ASAP7_75t_L g1183 ( .A1(n_768), .A2(n_1184), .A3(n_1186), .B1(n_1190), .B2(n_1194), .B3(n_1195), .Y(n_1183) );
BUFx3_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g1624 ( .A1(n_771), .A2(n_929), .B1(n_1619), .B2(n_1625), .Y(n_1624) );
BUFx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_773), .A2(n_781), .B1(n_794), .B2(n_813), .Y(n_844) );
INVx8_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
A2O1A1Ixp33_ASAP7_75t_L g866 ( .A1(n_781), .A2(n_867), .B(n_868), .C(n_869), .Y(n_866) );
INVx3_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx3_ASAP7_75t_L g1202 ( .A(n_784), .Y(n_1202) );
NOR3xp33_ASAP7_75t_L g1330 ( .A(n_784), .B(n_1331), .C(n_1343), .Y(n_1330) );
INVx1_ASAP7_75t_L g979 ( .A(n_786), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .B1(n_850), .B2(n_978), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OAI21x1_ASAP7_75t_SL g789 ( .A1(n_790), .A2(n_791), .B(n_849), .Y(n_789) );
NAND4xp25_ASAP7_75t_L g849 ( .A(n_790), .B(n_793), .C(n_795), .D(n_824), .Y(n_849) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_795), .C(n_824), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_802), .Y(n_795) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND3xp33_ASAP7_75t_SL g802 ( .A(n_803), .B(n_809), .C(n_814), .Y(n_802) );
HB1xp67_ASAP7_75t_L g1158 ( .A(n_807), .Y(n_1158) );
AOI22xp33_ASAP7_75t_SL g809 ( .A1(n_810), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g1660 ( .A1(n_810), .A2(n_812), .B1(n_1625), .B2(n_1627), .Y(n_1660) );
NAND3xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_818), .C(n_819), .Y(n_814) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_818), .Y(n_904) );
AOI211xp5_ASAP7_75t_L g957 ( .A1(n_818), .A2(n_958), .B(n_966), .C(n_974), .Y(n_957) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NAND3xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_830), .C(n_840), .Y(n_825) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_832), .B1(n_835), .B2(n_837), .Y(n_830) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g1125 ( .A1(n_839), .A2(n_1065), .B1(n_1126), .B2(n_1127), .Y(n_1125) );
OAI21xp5_ASAP7_75t_L g1332 ( .A1(n_839), .A2(n_1333), .B(n_1334), .Y(n_1332) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_843), .A2(n_894), .B1(n_1324), .B2(n_1339), .C(n_1340), .Y(n_1338) );
OAI22xp5_ASAP7_75t_L g1640 ( .A1(n_843), .A2(n_1641), .B1(n_1642), .B2(n_1643), .Y(n_1640) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_847), .B(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g978 ( .A(n_850), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B1(n_918), .B2(n_977), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
NAND4xp75_ASAP7_75t_L g855 ( .A(n_856), .B(n_899), .C(n_912), .D(n_915), .Y(n_855) );
OAI21x1_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_870), .B(n_897), .Y(n_856) );
OAI21xp5_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_859), .B(n_866), .Y(n_857) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx2_ASAP7_75t_L g1341 ( .A(n_862), .Y(n_1341) );
INVx2_ASAP7_75t_L g930 ( .A(n_865), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_877), .B1(n_882), .B2(n_891), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_873), .B1(n_875), .B2(n_876), .Y(n_871) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
OAI221xp5_ASAP7_75t_L g905 ( .A1(n_875), .A2(n_892), .B1(n_906), .B2(n_908), .C(n_910), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g1248 ( .A1(n_876), .A2(n_1249), .B1(n_1250), .B2(n_1251), .C(n_1252), .Y(n_1248) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g893 ( .A(n_880), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_883), .A2(n_884), .B1(n_887), .B2(n_888), .Y(n_882) );
BUFx4f_ASAP7_75t_SL g884 ( .A(n_885), .Y(n_884) );
INVx3_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx2_ASAP7_75t_SL g1000 ( .A(n_886), .Y(n_1000) );
OAI21xp33_ASAP7_75t_L g1335 ( .A1(n_888), .A2(n_1336), .B(n_1337), .Y(n_1335) );
INVx3_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
BUFx2_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
OAI21xp33_ASAP7_75t_L g1059 ( .A1(n_893), .A2(n_1060), .B(n_1061), .Y(n_1059) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
AOI211x1_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_901), .B(n_903), .C(n_911), .Y(n_899) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
OAI22xp33_ASAP7_75t_L g961 ( .A1(n_908), .A2(n_962), .B1(n_963), .B2(n_965), .Y(n_961) );
INVx6_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g977 ( .A(n_918), .Y(n_977) );
BUFx2_ASAP7_75t_SL g918 ( .A(n_919), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g919 ( .A1(n_920), .A2(n_975), .B(n_976), .Y(n_919) );
AND3x1_ASAP7_75t_L g920 ( .A(n_921), .B(n_951), .C(n_957), .Y(n_920) );
AOI31xp33_ASAP7_75t_L g976 ( .A1(n_921), .A2(n_951), .A3(n_957), .B(n_975), .Y(n_976) );
NAND3xp33_ASAP7_75t_SL g922 ( .A(n_923), .B(n_936), .C(n_939), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g923 ( .A1(n_924), .A2(n_928), .B1(n_931), .B2(n_934), .Y(n_923) );
BUFx2_ASAP7_75t_SL g1185 ( .A(n_925), .Y(n_1185) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVxp67_ASAP7_75t_L g1623 ( .A(n_940), .Y(n_1623) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_944), .A2(n_945), .B1(n_946), .B2(n_947), .Y(n_943) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_947), .Y(n_1004) );
INVx1_ASAP7_75t_L g1083 ( .A(n_950), .Y(n_1083) );
AND2x2_ASAP7_75t_L g951 ( .A(n_952), .B(n_954), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_956), .Y(n_954) );
INVx3_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
BUFx6f_ASAP7_75t_L g1034 ( .A(n_964), .Y(n_1034) );
INVx4_ASAP7_75t_L g1297 ( .A(n_964), .Y(n_1297) );
INVx1_ASAP7_75t_L g1037 ( .A(n_972), .Y(n_1037) );
BUFx6f_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
XNOR2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_1204), .Y(n_981) );
OA22x2_ASAP7_75t_L g982 ( .A1(n_983), .A2(n_1049), .B1(n_1050), .B2(n_1203), .Y(n_982) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g1203 ( .A(n_984), .Y(n_1203) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
NOR2x1_ASAP7_75t_L g986 ( .A(n_987), .B(n_1019), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g1074 ( .A(n_990), .Y(n_1074) );
NAND3xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_1006), .C(n_1013), .Y(n_996) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx2_ASAP7_75t_SL g999 ( .A(n_1000), .Y(n_999) );
OR2x6_ASAP7_75t_L g1197 ( .A(n_1000), .B(n_1198), .Y(n_1197) );
OAI22xp5_ASAP7_75t_SL g1032 ( .A1(n_1001), .A2(n_1033), .B1(n_1035), .B2(n_1036), .Y(n_1032) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1008), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_1014), .A2(n_1015), .B1(n_1017), .B2(n_1018), .Y(n_1013) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1015), .Y(n_1078) );
AOI22xp5_ASAP7_75t_L g1108 ( .A1(n_1015), .A2(n_1018), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1018), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1038), .Y(n_1019) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_SL g1027 ( .A(n_1028), .Y(n_1027) );
OAI221xp5_ASAP7_75t_L g1168 ( .A1(n_1033), .A2(n_1169), .B1(n_1170), .B2(n_1171), .C(n_1172), .Y(n_1168) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx3_ASAP7_75t_L g1390 ( .A(n_1034), .Y(n_1390) );
AOI21xp5_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1040), .B(n_1042), .Y(n_1038) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
XNOR2xp5_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1147), .Y(n_1050) );
XNOR2xp5_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1103), .Y(n_1051) );
OR2x2_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1084), .Y(n_1053) );
A2O1A1Ixp33_ASAP7_75t_SL g1054 ( .A1(n_1055), .A2(n_1073), .B(n_1080), .C(n_1081), .Y(n_1054) );
OAI21xp33_ASAP7_75t_L g1058 ( .A1(n_1059), .A2(n_1062), .B(n_1068), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1064), .B1(n_1065), .B2(n_1067), .Y(n_1062) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1063), .Y(n_1274) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
OAI211xp5_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1070), .B(n_1071), .C(n_1072), .Y(n_1068) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1080), .Y(n_1237) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1080), .Y(n_1644) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1083), .Y(n_1081) );
NAND3xp33_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1100), .C(n_1102), .Y(n_1084) );
NOR2xp33_ASAP7_75t_SL g1085 ( .A(n_1086), .B(n_1099), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_1088), .A2(n_1089), .B1(n_1090), .B2(n_1091), .Y(n_1087) );
XOR2x2_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1146), .Y(n_1103) );
NOR2xp33_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1128), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_1116), .A2(n_1119), .B1(n_1122), .B2(n_1125), .Y(n_1115) );
NAND4xp25_ASAP7_75t_SL g1128 ( .A(n_1129), .B(n_1130), .C(n_1132), .D(n_1135), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1648 ( .A(n_1140), .Y(n_1648) );
INVx2_ASAP7_75t_SL g1140 ( .A(n_1141), .Y(n_1140) );
NAND3xp33_ASAP7_75t_SL g1148 ( .A(n_1149), .B(n_1175), .C(n_1178), .Y(n_1148) );
OAI21xp33_ASAP7_75t_L g1149 ( .A1(n_1150), .A2(n_1165), .B(n_1174), .Y(n_1149) );
BUFx2_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1154), .Y(n_1294) );
HB1xp67_ASAP7_75t_SL g1155 ( .A(n_1156), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_1160), .A2(n_1161), .B1(n_1162), .B2(n_1163), .Y(n_1159) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
BUFx2_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
NOR3xp33_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1196), .C(n_1201), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1183), .Y(n_1179) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
CKINVDCx5p33_ASAP7_75t_R g1342 ( .A(n_1194), .Y(n_1342) );
INVxp67_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_SL g1201 ( .A(n_1202), .Y(n_1201) );
AOI22xp5_ASAP7_75t_L g1204 ( .A1(n_1205), .A2(n_1354), .B1(n_1355), .B2(n_1398), .Y(n_1204) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1205), .Y(n_1398) );
XOR2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1263), .Y(n_1205) );
XNOR2x1_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1208), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1256), .Y(n_1208) );
AOI221xp5_ASAP7_75t_L g1209 ( .A1(n_1210), .A2(n_1211), .B1(n_1212), .B2(n_1236), .C(n_1238), .Y(n_1209) );
NAND3xp33_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1225), .C(n_1233), .Y(n_1212) );
AOI222xp33_ASAP7_75t_L g1213 ( .A1(n_1214), .A2(n_1218), .B1(n_1219), .B2(n_1221), .C1(n_1222), .C2(n_1224), .Y(n_1213) );
BUFx2_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx2_ASAP7_75t_L g1319 ( .A(n_1217), .Y(n_1319) );
INVx2_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
CKINVDCx20_ASAP7_75t_R g1334 ( .A(n_1244), .Y(n_1334) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
XNOR2xp5_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1308), .Y(n_1263) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1284), .Y(n_1265) );
NOR3xp33_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1269), .C(n_1273), .Y(n_1267) );
NAND4xp25_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1288), .C(n_1304), .D(n_1306), .Y(n_1284) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
AND4x1_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1330), .C(n_1348), .D(n_1352), .Y(n_1309) );
INVx2_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
OAI211xp5_ASAP7_75t_L g1323 ( .A1(n_1324), .A2(n_1325), .B(n_1326), .C(n_1327), .Y(n_1323) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_1332), .A2(n_1335), .B1(n_1338), .B2(n_1342), .Y(n_1331) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
AOI211x1_ASAP7_75t_L g1356 ( .A1(n_1357), .A2(n_1375), .B(n_1376), .C(n_1382), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1362), .Y(n_1357) );
NOR3xp33_ASAP7_75t_L g1362 ( .A(n_1363), .B(n_1370), .C(n_1371), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g1385 ( .A1(n_1365), .A2(n_1386), .B1(n_1387), .B2(n_1388), .Y(n_1385) );
OAI22xp5_ASAP7_75t_L g1389 ( .A1(n_1367), .A2(n_1374), .B1(n_1390), .B2(n_1391), .Y(n_1389) );
OAI221xp5_ASAP7_75t_L g1399 ( .A1(n_1400), .A2(n_1607), .B1(n_1610), .B2(n_1666), .C(n_1671), .Y(n_1399) );
AND4x1_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1562), .C(n_1580), .D(n_1596), .Y(n_1400) );
OAI33xp33_ASAP7_75t_L g1401 ( .A1(n_1402), .A2(n_1494), .A3(n_1512), .B1(n_1518), .B2(n_1530), .B3(n_1541), .Y(n_1401) );
OAI211xp5_ASAP7_75t_SL g1402 ( .A1(n_1403), .A2(n_1422), .B(n_1443), .C(n_1475), .Y(n_1402) );
INVx2_ASAP7_75t_L g1496 ( .A(n_1403), .Y(n_1496) );
AOI331xp33_ASAP7_75t_L g1519 ( .A1(n_1403), .A2(n_1424), .A3(n_1489), .B1(n_1517), .B2(n_1520), .B3(n_1522), .C1(n_1523), .Y(n_1519) );
NOR2xp33_ASAP7_75t_L g1554 ( .A(n_1403), .B(n_1445), .Y(n_1554) );
NOR2xp33_ASAP7_75t_L g1597 ( .A(n_1403), .B(n_1425), .Y(n_1597) );
OR2x2_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1418), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1404), .B(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1404), .Y(n_1467) );
INVx2_ASAP7_75t_SL g1488 ( .A(n_1404), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1404), .B(n_1425), .Y(n_1553) );
NAND2xp5_ASAP7_75t_L g1599 ( .A(n_1404), .B(n_1600), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1412), .Y(n_1404) );
AND2x6_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1408), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1407), .B(n_1411), .Y(n_1410) );
AND2x4_ASAP7_75t_L g1413 ( .A(n_1407), .B(n_1414), .Y(n_1413) );
AND2x6_ASAP7_75t_L g1416 ( .A(n_1407), .B(n_1417), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1407), .B(n_1411), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1407), .B(n_1411), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1409), .B(n_1415), .Y(n_1414) );
INVx2_ASAP7_75t_L g1609 ( .A(n_1416), .Y(n_1609) );
HB1xp67_ASAP7_75t_L g1683 ( .A(n_1417), .Y(n_1683) );
CKINVDCx5p33_ASAP7_75t_R g1460 ( .A(n_1418), .Y(n_1460) );
NAND2xp5_ASAP7_75t_L g1466 ( .A(n_1418), .B(n_1467), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1484 ( .A(n_1418), .B(n_1426), .Y(n_1484) );
NAND2xp5_ASAP7_75t_L g1524 ( .A(n_1418), .B(n_1525), .Y(n_1524) );
AOI22xp5_ASAP7_75t_L g1531 ( .A1(n_1418), .A2(n_1510), .B1(n_1532), .B2(n_1535), .Y(n_1531) );
OAI22xp5_ASAP7_75t_L g1571 ( .A1(n_1418), .A2(n_1504), .B1(n_1572), .B2(n_1578), .Y(n_1571) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1418), .B(n_1455), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1418), .B(n_1456), .Y(n_1606) );
AND2x4_ASAP7_75t_L g1418 ( .A(n_1419), .B(n_1421), .Y(n_1418) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1429), .Y(n_1423) );
O2A1O1Ixp33_ASAP7_75t_SL g1468 ( .A1(n_1424), .A2(n_1469), .B(n_1470), .C(n_1472), .Y(n_1468) );
NAND2xp5_ASAP7_75t_L g1582 ( .A(n_1424), .B(n_1583), .Y(n_1582) );
CKINVDCx14_ASAP7_75t_R g1424 ( .A(n_1425), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1425), .B(n_1430), .Y(n_1501) );
NOR2xp33_ASAP7_75t_L g1503 ( .A(n_1425), .B(n_1504), .Y(n_1503) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1425), .B(n_1464), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1511 ( .A(n_1425), .B(n_1496), .Y(n_1511) );
NAND2xp5_ASAP7_75t_L g1533 ( .A(n_1425), .B(n_1534), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_1425), .B(n_1429), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1568 ( .A(n_1425), .B(n_1488), .Y(n_1568) );
INVx3_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
CKINVDCx5p33_ASAP7_75t_R g1449 ( .A(n_1426), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1426), .B(n_1471), .Y(n_1470) );
OR2x2_ASAP7_75t_L g1498 ( .A(n_1426), .B(n_1499), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1426), .B(n_1431), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1528 ( .A(n_1426), .B(n_1504), .Y(n_1528) );
AND2x4_ASAP7_75t_SL g1426 ( .A(n_1427), .B(n_1428), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1430), .B(n_1434), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1451 ( .A(n_1430), .B(n_1440), .Y(n_1451) );
OR2x2_ASAP7_75t_L g1462 ( .A(n_1430), .B(n_1463), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1430), .B(n_1483), .Y(n_1482) );
NAND2xp5_ASAP7_75t_L g1521 ( .A(n_1430), .B(n_1477), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1430), .B(n_1464), .Y(n_1545) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_1430), .B(n_1435), .Y(n_1550) );
OR2x2_ASAP7_75t_L g1561 ( .A(n_1430), .B(n_1446), .Y(n_1561) );
OR2x2_ASAP7_75t_L g1590 ( .A(n_1430), .B(n_1508), .Y(n_1590) );
INVx2_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
OR2x2_ASAP7_75t_L g1445 ( .A(n_1431), .B(n_1446), .Y(n_1445) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_1431), .B(n_1440), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1431), .B(n_1477), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1431), .B(n_1447), .Y(n_1486) );
OR2x2_ASAP7_75t_L g1499 ( .A(n_1431), .B(n_1436), .Y(n_1499) );
AND2x2_ASAP7_75t_L g1516 ( .A(n_1431), .B(n_1517), .Y(n_1516) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_1431), .B(n_1478), .Y(n_1527) );
NAND2xp5_ASAP7_75t_L g1577 ( .A(n_1431), .B(n_1436), .Y(n_1577) );
NOR2xp33_ASAP7_75t_L g1592 ( .A(n_1431), .B(n_1593), .Y(n_1592) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1433), .Y(n_1431) );
NOR2xp33_ASAP7_75t_L g1593 ( .A(n_1434), .B(n_1471), .Y(n_1593) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1439), .Y(n_1435) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1436), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1436), .B(n_1440), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1438), .Y(n_1436) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
OR2x2_ASAP7_75t_L g1446 ( .A(n_1440), .B(n_1447), .Y(n_1446) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1440), .Y(n_1478) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1440), .Y(n_1483) );
NAND2x1_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1442), .Y(n_1440) );
AOI221xp5_ASAP7_75t_L g1443 ( .A1(n_1444), .A2(n_1452), .B1(n_1461), .B2(n_1465), .C(n_1468), .Y(n_1443) );
NAND2xp5_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1448), .Y(n_1444) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1445), .Y(n_1583) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1446), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1447), .B(n_1478), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1449), .B(n_1450), .Y(n_1448) );
OR2x2_ASAP7_75t_L g1514 ( .A(n_1449), .B(n_1451), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1449), .B(n_1477), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_1449), .B(n_1486), .Y(n_1535) );
OR2x2_ASAP7_75t_L g1547 ( .A(n_1449), .B(n_1466), .Y(n_1547) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1449), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1449), .B(n_1527), .Y(n_1587) );
AOI22xp5_ASAP7_75t_L g1538 ( .A1(n_1450), .A2(n_1460), .B1(n_1505), .B2(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
NAND2xp5_ASAP7_75t_L g1529 ( .A(n_1452), .B(n_1461), .Y(n_1529) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1453 ( .A(n_1454), .B(n_1459), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1455), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1455), .B(n_1473), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1594 ( .A(n_1455), .B(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1456), .Y(n_1489) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1456), .Y(n_1507) );
AND2x2_ASAP7_75t_L g1522 ( .A(n_1456), .B(n_1460), .Y(n_1522) );
NAND2xp5_ASAP7_75t_L g1552 ( .A(n_1456), .B(n_1553), .Y(n_1552) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1456), .B(n_1568), .Y(n_1567) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1457), .B(n_1458), .Y(n_1456) );
OR2x2_ASAP7_75t_L g1487 ( .A(n_1460), .B(n_1488), .Y(n_1487) );
OAI32xp33_ASAP7_75t_L g1500 ( .A1(n_1460), .A2(n_1469), .A3(n_1477), .B1(n_1501), .B2(n_1502), .Y(n_1500) );
HB1xp67_ASAP7_75t_SL g1513 ( .A(n_1460), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1460), .B(n_1507), .Y(n_1573) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
OR2x2_ASAP7_75t_L g1601 ( .A(n_1463), .B(n_1501), .Y(n_1601) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1464), .B(n_1506), .Y(n_1505) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1466), .Y(n_1595) );
INVx2_ASAP7_75t_L g1473 ( .A(n_1467), .Y(n_1473) );
AOI31xp33_ASAP7_75t_L g1584 ( .A1(n_1467), .A2(n_1544), .A3(n_1585), .B(n_1586), .Y(n_1584) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1469), .Y(n_1510) );
NAND2xp5_ASAP7_75t_L g1520 ( .A(n_1469), .B(n_1521), .Y(n_1520) );
OAI221xp5_ASAP7_75t_L g1530 ( .A1(n_1472), .A2(n_1489), .B1(n_1531), .B2(n_1536), .C(n_1538), .Y(n_1530) );
OR2x2_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1474), .Y(n_1472) );
OAI221xp5_ASAP7_75t_SL g1494 ( .A1(n_1473), .A2(n_1495), .B1(n_1507), .B2(n_1508), .C(n_1509), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1473), .B(n_1505), .Y(n_1579) );
AOI221xp5_ASAP7_75t_L g1475 ( .A1(n_1476), .A2(n_1479), .B1(n_1480), .B2(n_1489), .C(n_1490), .Y(n_1475) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1476), .Y(n_1603) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1477), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1477), .B(n_1506), .Y(n_1575) );
OAI22xp33_ASAP7_75t_L g1480 ( .A1(n_1481), .A2(n_1484), .B1(n_1485), .B2(n_1487), .Y(n_1480) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVxp33_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1487), .Y(n_1534) );
INVx2_ASAP7_75t_L g1504 ( .A(n_1488), .Y(n_1504) );
O2A1O1Ixp33_ASAP7_75t_L g1512 ( .A1(n_1488), .A2(n_1513), .B(n_1514), .C(n_1515), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_1488), .B(n_1505), .Y(n_1564) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1489), .Y(n_1563) );
AOI221xp5_ASAP7_75t_L g1596 ( .A1(n_1489), .A2(n_1583), .B1(n_1597), .B2(n_1598), .C(n_1602), .Y(n_1596) );
INVx3_ASAP7_75t_L g1555 ( .A(n_1490), .Y(n_1555) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1491), .B(n_1493), .Y(n_1490) );
AOI211xp5_ASAP7_75t_L g1495 ( .A1(n_1496), .A2(n_1497), .B(n_1500), .C(n_1505), .Y(n_1495) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_1504), .B(n_1522), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1511), .Y(n_1509) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1511), .Y(n_1566) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
NAND2xp5_ASAP7_75t_L g1518 ( .A(n_1519), .B(n_1529), .Y(n_1518) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1522), .Y(n_1558) );
AOI22xp5_ASAP7_75t_L g1572 ( .A1(n_1522), .A2(n_1573), .B1(n_1574), .B2(n_1576), .Y(n_1572) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
INVxp33_ASAP7_75t_SL g1604 ( .A(n_1525), .Y(n_1604) );
NOR2xp33_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1528), .Y(n_1525) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1535), .Y(n_1585) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
NAND3xp33_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1548), .C(n_1556), .Y(n_1541) );
INVxp67_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
AOI21xp33_ASAP7_75t_L g1543 ( .A1(n_1544), .A2(n_1546), .B(n_1547), .Y(n_1543) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
NOR2xp33_ASAP7_75t_L g1569 ( .A(n_1545), .B(n_1570), .Y(n_1569) );
AOI211xp5_ASAP7_75t_L g1548 ( .A1(n_1549), .A2(n_1551), .B(n_1554), .C(n_1555), .Y(n_1548) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
NOR2xp33_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1559), .Y(n_1557) );
OR2x2_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1561), .Y(n_1559) );
INVx2_ASAP7_75t_L g1570 ( .A(n_1561), .Y(n_1570) );
AOI211xp5_ASAP7_75t_L g1562 ( .A1(n_1563), .A2(n_1564), .B(n_1565), .C(n_1571), .Y(n_1562) );
AOI21xp33_ASAP7_75t_L g1565 ( .A1(n_1566), .A2(n_1567), .B(n_1569), .Y(n_1565) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
INVxp33_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
O2A1O1Ixp33_ASAP7_75t_L g1580 ( .A1(n_1581), .A2(n_1584), .B(n_1588), .C(n_1589), .Y(n_1580) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
AOI21xp5_ASAP7_75t_L g1589 ( .A1(n_1590), .A2(n_1591), .B(n_1594), .Y(n_1589) );
INVxp33_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
INVxp67_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
AOI21xp33_ASAP7_75t_L g1602 ( .A1(n_1603), .A2(n_1604), .B(n_1605), .Y(n_1602) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
CKINVDCx20_ASAP7_75t_R g1607 ( .A(n_1608), .Y(n_1607) );
CKINVDCx20_ASAP7_75t_R g1608 ( .A(n_1609), .Y(n_1608) );
HB1xp67_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
HB1xp67_ASAP7_75t_L g1679 ( .A(n_1612), .Y(n_1679) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
NAND3xp33_ASAP7_75t_L g1613 ( .A(n_1614), .B(n_1621), .C(n_1645), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1618), .Y(n_1616) );
OAI21xp33_ASAP7_75t_L g1621 ( .A1(n_1622), .A2(n_1634), .B(n_1644), .Y(n_1621) );
OAI211xp5_ASAP7_75t_L g1622 ( .A1(n_1623), .A2(n_1624), .B(n_1626), .C(n_1629), .Y(n_1622) );
OAI211xp5_ASAP7_75t_L g1629 ( .A1(n_1630), .A2(n_1631), .B(n_1632), .C(n_1633), .Y(n_1629) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
NOR3xp33_ASAP7_75t_L g1645 ( .A(n_1646), .B(n_1654), .C(n_1661), .Y(n_1645) );
INVxp67_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
INVx2_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
CKINVDCx20_ASAP7_75t_R g1666 ( .A(n_1667), .Y(n_1666) );
CKINVDCx20_ASAP7_75t_R g1667 ( .A(n_1668), .Y(n_1667) );
INVx3_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
HB1xp67_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
BUFx3_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
INVxp67_ASAP7_75t_SL g1677 ( .A(n_1678), .Y(n_1677) );
INVx2_ASAP7_75t_SL g1680 ( .A(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
OAI21xp5_ASAP7_75t_L g1682 ( .A1(n_1683), .A2(n_1684), .B(n_1685), .Y(n_1682) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
endmodule