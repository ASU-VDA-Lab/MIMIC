module fake_ibex_67_n_2271 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_403, n_423, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_426, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_427, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_414, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_428, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2271);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_428;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2271;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2163;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2189;
wire n_745;
wire n_2112;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_2256;
wire n_737;
wire n_606;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_1543;
wire n_823;
wire n_2233;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1793;
wire n_1237;
wire n_859;
wire n_1109;
wire n_965;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_585;
wire n_1982;
wire n_2252;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_2243;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_961;
wire n_634;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_1353;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1415;
wire n_1238;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_950;
wire n_512;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_2225;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_1788;
wire n_2093;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_753;
wire n_2126;
wire n_747;
wire n_1147;
wire n_645;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_470;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2079;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1397;
wire n_1211;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2092;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2262;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_1902;
wire n_1194;
wire n_683;
wire n_1150;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

BUFx3_ASAP7_75t_L g430 ( 
.A(n_70),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_37),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_290),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_419),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_351),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_266),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_45),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_41),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_40),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_380),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_28),
.Y(n_440)
);

BUFx10_ASAP7_75t_L g441 ( 
.A(n_260),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_52),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_273),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_258),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_360),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_373),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_269),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_425),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_87),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_294),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_167),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_302),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_150),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_92),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_283),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_404),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_258),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_163),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_386),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_274),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_285),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_276),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_407),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_150),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_391),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_308),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_43),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_320),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_397),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_307),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_229),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_28),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_335),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_151),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_345),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_0),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_51),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_231),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_179),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_85),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_309),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_108),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_36),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_70),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_147),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_187),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_138),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_116),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_207),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_322),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_259),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_297),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_126),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_180),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_96),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_111),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_184),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_146),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_261),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_253),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_298),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_61),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_18),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_92),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_123),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_187),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_158),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_245),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_195),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_55),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_207),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_48),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_189),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_175),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_41),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_186),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_62),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_182),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_376),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_111),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_381),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_180),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_112),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_206),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_305),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_193),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_336),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_62),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_5),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_186),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_228),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_0),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_282),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_275),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_68),
.Y(n_537)
);

BUFx10_ASAP7_75t_L g538 ( 
.A(n_357),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_257),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_139),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_347),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_325),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_256),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_162),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_131),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_340),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_301),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_371),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_318),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_191),
.Y(n_550)
);

BUFx8_ASAP7_75t_SL g551 ( 
.A(n_133),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_106),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_312),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_326),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_368),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_402),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_219),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_226),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_375),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_141),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_311),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_191),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_383),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_223),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_310),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_63),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_178),
.Y(n_567)
);

INVx4_ASAP7_75t_R g568 ( 
.A(n_323),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_136),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_68),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_66),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_159),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_427),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_93),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_316),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_356),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_230),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_330),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_422),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_100),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_167),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_416),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_366),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_141),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_129),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_2),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_235),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_60),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_300),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_132),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_213),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_327),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_395),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_254),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_296),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_55),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_315),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_409),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_385),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_225),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_16),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_429),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_134),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_163),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_204),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_83),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_169),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_251),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_154),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_244),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_174),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_135),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_123),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_72),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_367),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_195),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_11),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_378),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_4),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_280),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_231),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_97),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_162),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_80),
.Y(n_624)
);

CKINVDCx16_ASAP7_75t_R g625 ( 
.A(n_410),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_19),
.Y(n_626)
);

CKINVDCx16_ASAP7_75t_R g627 ( 
.A(n_176),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_71),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_243),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_218),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_329),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_426),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_165),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_130),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_408),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_67),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_52),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_74),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_2),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_412),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_135),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_133),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_203),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_321),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_350),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_152),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_263),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_281),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_56),
.Y(n_649)
);

CKINVDCx16_ASAP7_75t_R g650 ( 
.A(n_38),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_382),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_32),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_400),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_287),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_355),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_27),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_11),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_252),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_333),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_74),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_136),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_104),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_374),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_58),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_205),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_264),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_424),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_232),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_238),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_342),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_372),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_159),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_337),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_411),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_168),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_38),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_354),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_369),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_200),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_148),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_97),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_401),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_85),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_223),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_64),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_107),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_379),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_394),
.Y(n_688)
);

BUFx10_ASAP7_75t_L g689 ( 
.A(n_80),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_220),
.Y(n_690)
);

CKINVDCx14_ASAP7_75t_R g691 ( 
.A(n_324),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_39),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_396),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_227),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_12),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_256),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_217),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_109),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_389),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_169),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_271),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_178),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_15),
.Y(n_703)
);

INVxp67_ASAP7_75t_SL g704 ( 
.A(n_115),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_44),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_334),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_377),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_370),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_414),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_157),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_127),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_313),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_183),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_496),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_446),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_591),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_591),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_529),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_488),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_627),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_669),
.B(n_1),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_591),
.Y(n_722)
);

INVxp67_ASAP7_75t_SL g723 ( 
.A(n_430),
.Y(n_723)
);

NOR2xp67_ASAP7_75t_L g724 ( 
.A(n_474),
.B(n_1),
.Y(n_724)
);

INVxp33_ASAP7_75t_SL g725 ( 
.A(n_611),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_430),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_554),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_576),
.B(n_3),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_535),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_494),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_559),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_711),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_576),
.B(n_3),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_582),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_521),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_589),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_474),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_650),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_623),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_635),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_473),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_623),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_672),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_672),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_703),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_647),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_708),
.B(n_4),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_495),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_703),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_494),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_620),
.B(n_6),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_653),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_453),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_670),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_520),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_453),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_499),
.Y(n_757)
);

NOR2xp67_ASAP7_75t_L g758 ( 
.A(n_451),
.B(n_6),
.Y(n_758)
);

BUFx6f_ASAP7_75t_SL g759 ( 
.A(n_441),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_436),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_701),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_546),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_571),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_619),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_502),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_619),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_565),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_479),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_479),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_630),
.Y(n_770)
);

XOR2xp5_ASAP7_75t_L g771 ( 
.A(n_504),
.B(n_7),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_436),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_514),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_702),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_625),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_702),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_437),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_551),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_454),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_620),
.B(n_8),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_522),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_534),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_567),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_587),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_607),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_458),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_520),
.B(n_8),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_629),
.Y(n_788)
);

INVxp33_ASAP7_75t_SL g789 ( 
.A(n_438),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_649),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_466),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_660),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_696),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_478),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_432),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_482),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_484),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_432),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_487),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_438),
.Y(n_800)
);

INVxp33_ASAP7_75t_SL g801 ( 
.A(n_440),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_440),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_442),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_500),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_505),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_507),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_442),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_444),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_510),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_511),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_592),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_729),
.B(n_444),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_737),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_735),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_739),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_735),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_722),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_723),
.B(n_449),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_735),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_726),
.B(n_449),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_735),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_742),
.B(n_459),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_722),
.B(n_524),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_722),
.B(n_528),
.Y(n_824)
);

AND2x6_ASAP7_75t_L g825 ( 
.A(n_747),
.B(n_787),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_743),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_744),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_730),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_745),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_749),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_766),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_714),
.B(n_732),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_760),
.B(n_691),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_716),
.B(n_459),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_766),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_750),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_766),
.Y(n_837)
);

INVx5_ASAP7_75t_L g838 ( 
.A(n_811),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_717),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_811),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_753),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_756),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_768),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_769),
.Y(n_844)
);

INVx6_ASAP7_75t_L g845 ( 
.A(n_759),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_789),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_763),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_764),
.B(n_531),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_770),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_SL g850 ( 
.A(n_759),
.B(n_433),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_780),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_774),
.Y(n_852)
);

BUFx8_ASAP7_75t_L g853 ( 
.A(n_759),
.Y(n_853)
);

OAI21x1_ASAP7_75t_L g854 ( 
.A1(n_777),
.A2(n_599),
.B(n_592),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_776),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_779),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_786),
.Y(n_857)
);

BUFx8_ASAP7_75t_L g858 ( 
.A(n_801),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_791),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_794),
.B(n_532),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_808),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_725),
.A2(n_661),
.B1(n_668),
.B2(n_469),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_796),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_797),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_728),
.B(n_599),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_795),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_799),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_804),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_805),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_806),
.B(n_543),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_809),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_755),
.B(n_618),
.Y(n_872)
);

NOR2x1_ASAP7_75t_L g873 ( 
.A(n_810),
.B(n_443),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_733),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_751),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_724),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_798),
.B(n_520),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_721),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_758),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_762),
.Y(n_880)
);

INVx5_ASAP7_75t_L g881 ( 
.A(n_767),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_775),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_800),
.B(n_469),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_800),
.B(n_606),
.Y(n_884)
);

NAND2x1_ASAP7_75t_L g885 ( 
.A(n_778),
.B(n_568),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_802),
.A2(n_668),
.B1(n_679),
.B2(n_661),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_802),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_807),
.B(n_618),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_803),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_807),
.B(n_679),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_803),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_715),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_771),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_718),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_727),
.B(n_680),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_738),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_731),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_734),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_736),
.B(n_680),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_740),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_719),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_719),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_720),
.B(n_545),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_746),
.B(n_606),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_752),
.B(n_681),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_754),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_720),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_761),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_765),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_773),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_781),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_782),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_741),
.B(n_552),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_783),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_748),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_748),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_757),
.Y(n_917)
);

INVx6_ASAP7_75t_L g918 ( 
.A(n_757),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_784),
.B(n_609),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_784),
.Y(n_920)
);

OAI21x1_ASAP7_75t_L g921 ( 
.A1(n_785),
.A2(n_455),
.B(n_452),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_785),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_788),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_788),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_790),
.B(n_684),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_790),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_792),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_793),
.B(n_685),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_735),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_735),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_737),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_737),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_780),
.B(n_456),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_737),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_722),
.A2(n_460),
.B(n_457),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_780),
.B(n_463),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_735),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_735),
.Y(n_938)
);

BUFx8_ASAP7_75t_L g939 ( 
.A(n_759),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_722),
.A2(n_468),
.B(n_464),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_737),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_780),
.B(n_475),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_737),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_737),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_780),
.B(n_477),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_735),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_722),
.B(n_560),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_737),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_735),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_737),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_735),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_737),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_737),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_735),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_735),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_737),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_735),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_808),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_722),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_735),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_737),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_737),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_735),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_729),
.B(n_690),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_735),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_737),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_722),
.A2(n_492),
.B(n_483),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_722),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_729),
.B(n_690),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_737),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_729),
.B(n_493),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_737),
.Y(n_972)
);

AND3x1_ASAP7_75t_L g973 ( 
.A(n_787),
.B(n_566),
.C(n_564),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_772),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_808),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_722),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_735),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_737),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_722),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_735),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_851),
.B(n_441),
.Y(n_981)
);

BUFx10_ASAP7_75t_L g982 ( 
.A(n_845),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_817),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_817),
.Y(n_984)
);

INVx8_ASAP7_75t_L g985 ( 
.A(n_825),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_853),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_835),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_874),
.B(n_712),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_959),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_859),
.B(n_434),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_959),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_832),
.B(n_609),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_959),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_831),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_831),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_878),
.B(n_860),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_935),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_831),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_874),
.B(n_875),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_974),
.B(n_609),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_853),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_861),
.B(n_694),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_846),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_L g1004 ( 
.A(n_973),
.B(n_698),
.C(n_697),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_878),
.B(n_441),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_859),
.A2(n_569),
.B1(n_586),
.B2(n_580),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_968),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_845),
.Y(n_1008)
);

AND2x6_ASAP7_75t_L g1009 ( 
.A(n_860),
.B(n_501),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_878),
.B(n_435),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_875),
.B(n_435),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_828),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_968),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_863),
.A2(n_867),
.B1(n_868),
.B2(n_860),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_863),
.A2(n_601),
.B1(n_605),
.B2(n_604),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_867),
.B(n_868),
.Y(n_1016)
);

INVx6_ASAP7_75t_L g1017 ( 
.A(n_939),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_976),
.Y(n_1018)
);

AND2x6_ASAP7_75t_L g1019 ( 
.A(n_870),
.B(n_523),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_828),
.Y(n_1020)
);

AND2x6_ASAP7_75t_L g1021 ( 
.A(n_870),
.B(n_527),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_833),
.B(n_689),
.Y(n_1022)
);

AND2x6_ASAP7_75t_L g1023 ( 
.A(n_870),
.B(n_541),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_848),
.B(n_850),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_818),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_935),
.B(n_555),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_979),
.Y(n_1027)
);

AND2x6_ASAP7_75t_L g1028 ( 
.A(n_873),
.B(n_563),
.Y(n_1028)
);

AND2x6_ASAP7_75t_L g1029 ( 
.A(n_823),
.B(n_573),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_940),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_979),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_813),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_856),
.A2(n_857),
.B1(n_869),
.B2(n_864),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_836),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_L g1035 ( 
.A(n_825),
.B(n_439),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_933),
.B(n_538),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_836),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_815),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_826),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_825),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_940),
.B(n_579),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_858),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_827),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_877),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_858),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_829),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_825),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_862),
.B(n_689),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_933),
.B(n_538),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_830),
.Y(n_1050)
);

INVx4_ASAP7_75t_L g1051 ( 
.A(n_881),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_967),
.B(n_693),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_866),
.B(n_705),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_931),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_871),
.B(n_445),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_848),
.B(n_445),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_967),
.B(n_699),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_866),
.B(n_697),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_848),
.B(n_820),
.Y(n_1059)
);

AND2x6_ASAP7_75t_L g1060 ( 
.A(n_823),
.B(n_583),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_852),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_852),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_888),
.A2(n_705),
.B1(n_698),
.B2(n_713),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_888),
.B(n_480),
.C(n_476),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_936),
.B(n_538),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_823),
.B(n_824),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_932),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_881),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_824),
.B(n_447),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_876),
.B(n_704),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_824),
.B(n_447),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_947),
.B(n_450),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_934),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_884),
.B(n_485),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_852),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_840),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_852),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_841),
.B(n_598),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_941),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_947),
.B(n_450),
.Y(n_1080)
);

AND2x6_ASAP7_75t_L g1081 ( 
.A(n_947),
.B(n_631),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_855),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_958),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_975),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_943),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_840),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_944),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_936),
.B(n_578),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_948),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_906),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_855),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_950),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_839),
.A2(n_614),
.B1(n_621),
.B2(n_617),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_881),
.Y(n_1094)
);

BUFx4f_ASAP7_75t_L g1095 ( 
.A(n_898),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_812),
.A2(n_710),
.B1(n_624),
.B2(n_628),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_952),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_837),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_881),
.Y(n_1099)
);

OR2x6_ASAP7_75t_L g1100 ( 
.A(n_898),
.B(n_562),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_837),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_883),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_843),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_890),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_906),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_854),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_925),
.B(n_481),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_942),
.B(n_578),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_822),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_847),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_SL g1111 ( 
.A(n_903),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_854),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_953),
.Y(n_1113)
);

AND2x2_ASAP7_75t_SL g1114 ( 
.A(n_903),
.B(n_431),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_847),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_918),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_956),
.Y(n_1117)
);

AND2x6_ASAP7_75t_L g1118 ( 
.A(n_904),
.B(n_632),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_961),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_847),
.B(n_648),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_843),
.Y(n_1121)
);

INVx4_ASAP7_75t_L g1122 ( 
.A(n_838),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_886),
.B(n_486),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_844),
.Y(n_1124)
);

AND2x6_ASAP7_75t_L g1125 ( 
.A(n_880),
.B(n_654),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_928),
.B(n_508),
.Y(n_1126)
);

NAND2xp33_ASAP7_75t_L g1127 ( 
.A(n_850),
.B(n_978),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_962),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_838),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_964),
.B(n_489),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_919),
.Y(n_1131)
);

OR2x6_ASAP7_75t_L g1132 ( 
.A(n_898),
.B(n_657),
.Y(n_1132)
);

INVx4_ASAP7_75t_SL g1133 ( 
.A(n_966),
.Y(n_1133)
);

NAND3xp33_ASAP7_75t_L g1134 ( 
.A(n_969),
.B(n_491),
.C(n_490),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_901),
.B(n_509),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_945),
.B(n_615),
.Y(n_1136)
);

INVx4_ASAP7_75t_L g1137 ( 
.A(n_838),
.Y(n_1137)
);

BUFx4_ASAP7_75t_L g1138 ( 
.A(n_911),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_970),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_971),
.A2(n_638),
.B1(n_652),
.B2(n_646),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_885),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_972),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_921),
.Y(n_1143)
);

BUFx10_ASAP7_75t_L g1144 ( 
.A(n_903),
.Y(n_1144)
);

BUFx10_ASAP7_75t_L g1145 ( 
.A(n_882),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_879),
.B(n_664),
.Y(n_1146)
);

BUFx8_ASAP7_75t_SL g1147 ( 
.A(n_914),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_834),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_945),
.B(n_615),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_901),
.B(n_544),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_842),
.B(n_659),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_849),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_902),
.B(n_584),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_849),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_892),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_918),
.Y(n_1156)
);

OAI221xp5_ASAP7_75t_L g1157 ( 
.A1(n_971),
.A2(n_665),
.B1(n_675),
.B2(n_662),
.C(n_658),
.Y(n_1157)
);

OR2x6_ASAP7_75t_L g1158 ( 
.A(n_892),
.B(n_897),
.Y(n_1158)
);

BUFx10_ASAP7_75t_L g1159 ( 
.A(n_872),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_865),
.B(n_461),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_921),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_892),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_865),
.B(n_461),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_872),
.B(n_894),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_895),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_899),
.B(n_462),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_905),
.B(n_682),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_918),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_913),
.B(n_497),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_816),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_897),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_913),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_913),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_814),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_814),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_900),
.B(n_615),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_908),
.A2(n_676),
.B1(n_686),
.B2(n_683),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_902),
.B(n_613),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_897),
.B(n_462),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_907),
.B(n_465),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_819),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_819),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_907),
.B(n_692),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_821),
.B(n_465),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_954),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_929),
.B(n_467),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_896),
.B(n_498),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_954),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_930),
.B(n_467),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_887),
.A2(n_700),
.B1(n_506),
.B2(n_513),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_914),
.Y(n_1191)
);

NAND2xp33_ASAP7_75t_L g1192 ( 
.A(n_954),
.B(n_709),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_889),
.B(n_470),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_955),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_891),
.B(n_512),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_986),
.B(n_917),
.Y(n_1196)
);

AO22x2_ASAP7_75t_L g1197 ( 
.A1(n_1161),
.A2(n_917),
.B1(n_926),
.B2(n_924),
.Y(n_1197)
);

OAI221xp5_ASAP7_75t_L g1198 ( 
.A1(n_1131),
.A2(n_927),
.B1(n_909),
.B2(n_920),
.C(n_922),
.Y(n_1198)
);

AO22x2_ASAP7_75t_L g1199 ( 
.A1(n_1083),
.A2(n_917),
.B1(n_923),
.B2(n_916),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_1003),
.Y(n_1200)
);

AO22x2_ASAP7_75t_L g1201 ( 
.A1(n_1083),
.A2(n_1004),
.B1(n_1047),
.B2(n_1040),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1003),
.B(n_915),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1114),
.A2(n_431),
.B1(n_516),
.B2(n_515),
.Y(n_1203)
);

AO22x2_ASAP7_75t_L g1204 ( 
.A1(n_1040),
.A2(n_912),
.B1(n_910),
.B2(n_893),
.Y(n_1204)
);

NOR2xp67_ASAP7_75t_L g1205 ( 
.A(n_1001),
.B(n_914),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1152),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1025),
.B(n_517),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1105),
.B(n_915),
.Y(n_1208)
);

OAI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1102),
.A2(n_695),
.B1(n_642),
.B2(n_616),
.C(n_525),
.Y(n_1209)
);

AO22x2_ASAP7_75t_L g1210 ( 
.A1(n_1047),
.A2(n_915),
.B1(n_914),
.B2(n_687),
.Y(n_1210)
);

AO22x2_ASAP7_75t_L g1211 ( 
.A1(n_1190),
.A2(n_915),
.B1(n_503),
.B2(n_548),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_996),
.B(n_471),
.Y(n_1212)
);

NAND2xp33_ASAP7_75t_L g1213 ( 
.A(n_1009),
.B(n_471),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1066),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1066),
.Y(n_1215)
);

AO22x2_ASAP7_75t_L g1216 ( 
.A1(n_1190),
.A2(n_549),
.B1(n_667),
.B2(n_448),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1032),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1102),
.A2(n_519),
.B1(n_526),
.B2(n_518),
.Y(n_1218)
);

BUFx8_ASAP7_75t_L g1219 ( 
.A(n_1111),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1025),
.B(n_530),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1042),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1038),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1171),
.B(n_472),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1109),
.B(n_663),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1039),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1148),
.B(n_663),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1152),
.Y(n_1227)
);

AO22x2_ASAP7_75t_L g1228 ( 
.A1(n_1172),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1053),
.B(n_533),
.Y(n_1229)
);

AO22x2_ASAP7_75t_L g1230 ( 
.A1(n_1173),
.A2(n_13),
.B1(n_9),
.B2(n_10),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1059),
.B(n_537),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1043),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1046),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1050),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1144),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1054),
.A2(n_539),
.B(n_550),
.C(n_540),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1067),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1104),
.A2(n_558),
.B1(n_570),
.B2(n_557),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1045),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1158),
.B(n_666),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1017),
.A2(n_574),
.B1(n_577),
.B2(n_572),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1073),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1154),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1079),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1158),
.B(n_666),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1059),
.B(n_581),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1085),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1087),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1089),
.Y(n_1249)
);

AO22x2_ASAP7_75t_L g1250 ( 
.A1(n_1168),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_SL g1251 ( 
.A(n_1100),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1092),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1097),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1113),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1117),
.Y(n_1255)
);

OAI221xp5_ASAP7_75t_L g1256 ( 
.A1(n_1104),
.A2(n_590),
.B1(n_594),
.B2(n_588),
.C(n_585),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1014),
.B(n_596),
.Y(n_1257)
);

AO22x2_ASAP7_75t_L g1258 ( 
.A1(n_1168),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1119),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1128),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1014),
.B(n_600),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1114),
.A2(n_673),
.B1(n_674),
.B2(n_671),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1033),
.B(n_1011),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1090),
.A2(n_608),
.B1(n_610),
.B2(n_603),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1139),
.Y(n_1265)
);

AO22x2_ASAP7_75t_L g1266 ( 
.A1(n_1024),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1266)
);

OAI221xp5_ASAP7_75t_L g1267 ( 
.A1(n_1177),
.A2(n_626),
.B1(n_633),
.B2(n_622),
.C(n_612),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1142),
.Y(n_1268)
);

OAI221xp5_ASAP7_75t_L g1269 ( 
.A1(n_1177),
.A2(n_637),
.B1(n_639),
.B2(n_636),
.C(n_634),
.Y(n_1269)
);

AO22x2_ASAP7_75t_L g1270 ( 
.A1(n_1183),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1158),
.B(n_671),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1165),
.B(n_673),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1011),
.B(n_641),
.Y(n_1273)
);

AO22x2_ASAP7_75t_L g1274 ( 
.A1(n_1183),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1008),
.B(n_674),
.Y(n_1275)
);

AO22x2_ASAP7_75t_L g1276 ( 
.A1(n_1162),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1084),
.Y(n_1277)
);

AO22x2_ASAP7_75t_L g1278 ( 
.A1(n_1096),
.A2(n_1002),
.B1(n_1058),
.B2(n_1123),
.Y(n_1278)
);

BUFx8_ASAP7_75t_L g1279 ( 
.A(n_1111),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1055),
.B(n_643),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1016),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1016),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1130),
.B(n_656),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1017),
.Y(n_1284)
);

AO22x2_ASAP7_75t_L g1285 ( 
.A1(n_1096),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1082),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_992),
.B(n_677),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1082),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1044),
.B(n_678),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1091),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1091),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1008),
.B(n_688),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_999),
.Y(n_1293)
);

AO22x2_ASAP7_75t_L g1294 ( 
.A1(n_1056),
.A2(n_30),
.B1(n_26),
.B2(n_29),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1017),
.B(n_985),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_999),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_1100),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1155),
.B(n_521),
.Y(n_1298)
);

AO22x2_ASAP7_75t_L g1299 ( 
.A1(n_1048),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1009),
.A2(n_707),
.B1(n_709),
.B2(n_706),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1110),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1110),
.Y(n_1302)
);

BUFx8_ASAP7_75t_L g1303 ( 
.A(n_1074),
.Y(n_1303)
);

AO22x2_ASAP7_75t_L g1304 ( 
.A1(n_1135),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1141),
.B(n_33),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1144),
.Y(n_1306)
);

AO22x2_ASAP7_75t_L g1307 ( 
.A1(n_1150),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1100),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1169),
.B(n_34),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1115),
.Y(n_1310)
);

OAI221xp5_ASAP7_75t_L g1311 ( 
.A1(n_1157),
.A2(n_1063),
.B1(n_1140),
.B2(n_1093),
.C(n_1006),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_990),
.Y(n_1312)
);

AO22x2_ASAP7_75t_L g1313 ( 
.A1(n_1153),
.A2(n_39),
.B1(n_35),
.B2(n_37),
.Y(n_1313)
);

AO22x2_ASAP7_75t_L g1314 ( 
.A1(n_1178),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_1314)
);

AO22x2_ASAP7_75t_L g1315 ( 
.A1(n_1107),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1000),
.B(n_46),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1126),
.B(n_47),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1103),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1007),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1022),
.B(n_47),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1013),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1027),
.Y(n_1322)
);

AO22x2_ASAP7_75t_L g1323 ( 
.A1(n_1064),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1323)
);

AO22x2_ASAP7_75t_L g1324 ( 
.A1(n_1069),
.A2(n_53),
.B1(n_49),
.B2(n_51),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1147),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1031),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1116),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1132),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1098),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1164),
.B(n_53),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1098),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1121),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1101),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1101),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1187),
.B(n_54),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1124),
.Y(n_1336)
);

AO22x2_ASAP7_75t_L g1337 ( 
.A1(n_1069),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1132),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_L g1339 ( 
.A(n_1134),
.B(n_57),
.Y(n_1339)
);

BUFx8_ASAP7_75t_L g1340 ( 
.A(n_1191),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_985),
.B(n_575),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_983),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_984),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_994),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_995),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1164),
.B(n_58),
.Y(n_1346)
);

INVxp67_ASAP7_75t_L g1347 ( 
.A(n_1005),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_989),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_998),
.Y(n_1349)
);

OR2x6_ASAP7_75t_L g1350 ( 
.A(n_985),
.B(n_575),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1005),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_991),
.Y(n_1352)
);

INVxp67_ASAP7_75t_L g1353 ( 
.A(n_1071),
.Y(n_1353)
);

AO22x2_ASAP7_75t_L g1354 ( 
.A1(n_1071),
.A2(n_63),
.B1(n_59),
.B2(n_60),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_993),
.Y(n_1355)
);

CKINVDCx16_ASAP7_75t_R g1356 ( 
.A(n_982),
.Y(n_1356)
);

AO22x2_ASAP7_75t_L g1357 ( 
.A1(n_1072),
.A2(n_65),
.B1(n_59),
.B2(n_64),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1072),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1080),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1080),
.Y(n_1360)
);

AO22x2_ASAP7_75t_L g1361 ( 
.A1(n_1143),
.A2(n_69),
.B1(n_65),
.B2(n_67),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_981),
.B(n_536),
.Y(n_1362)
);

AO22x2_ASAP7_75t_L g1363 ( 
.A1(n_1143),
.A2(n_72),
.B1(n_69),
.B2(n_71),
.Y(n_1363)
);

AO22x2_ASAP7_75t_L g1364 ( 
.A1(n_1026),
.A2(n_76),
.B1(n_73),
.B2(n_75),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1018),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1193),
.B(n_547),
.C(n_542),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1179),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1018),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1151),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1156),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1151),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_997),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1075),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1009),
.A2(n_556),
.B1(n_561),
.B2(n_553),
.Y(n_1374)
);

AO22x2_ASAP7_75t_L g1375 ( 
.A1(n_1026),
.A2(n_1041),
.B1(n_1057),
.B2(n_1052),
.Y(n_1375)
);

AO22x2_ASAP7_75t_L g1376 ( 
.A1(n_1041),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1180),
.Y(n_1377)
);

AO22x2_ASAP7_75t_L g1378 ( 
.A1(n_1052),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1378)
);

NAND2x1p5_ASAP7_75t_L g1379 ( 
.A(n_1095),
.B(n_575),
.Y(n_1379)
);

NAND2x1p5_ASAP7_75t_L g1380 ( 
.A(n_1051),
.B(n_640),
.Y(n_1380)
);

BUFx8_ASAP7_75t_L g1381 ( 
.A(n_1019),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1180),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1051),
.B(n_640),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_988),
.Y(n_1384)
);

OAI221xp5_ASAP7_75t_L g1385 ( 
.A1(n_1140),
.A2(n_597),
.B1(n_602),
.B2(n_595),
.C(n_593),
.Y(n_1385)
);

AO22x2_ASAP7_75t_L g1386 ( 
.A1(n_1057),
.A2(n_81),
.B1(n_78),
.B2(n_79),
.Y(n_1386)
);

NAND2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1068),
.B(n_640),
.Y(n_1387)
);

NAND2x1p5_ASAP7_75t_L g1388 ( 
.A(n_1068),
.B(n_640),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1078),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1078),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1019),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1120),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1120),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1070),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_981),
.B(n_644),
.Y(n_1395)
);

AO22x2_ASAP7_75t_L g1396 ( 
.A1(n_1070),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1138),
.B(n_1195),
.Y(n_1397)
);

AO22x2_ASAP7_75t_L g1398 ( 
.A1(n_1133),
.A2(n_86),
.B1(n_82),
.B2(n_84),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1021),
.Y(n_1399)
);

AO22x2_ASAP7_75t_L g1400 ( 
.A1(n_1133),
.A2(n_88),
.B1(n_84),
.B2(n_86),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1179),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1160),
.Y(n_1402)
);

AO22x2_ASAP7_75t_L g1403 ( 
.A1(n_1133),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_982),
.B(n_645),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1160),
.Y(n_1405)
);

OAI221xp5_ASAP7_75t_L g1406 ( 
.A1(n_1093),
.A2(n_655),
.B1(n_651),
.B2(n_938),
.C(n_937),
.Y(n_1406)
);

AO22x2_ASAP7_75t_L g1407 ( 
.A1(n_1146),
.A2(n_93),
.B1(n_90),
.B2(n_91),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1010),
.B(n_91),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1163),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1163),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1122),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1021),
.A2(n_946),
.B1(n_949),
.B2(n_938),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1023),
.A2(n_1029),
.B1(n_1081),
.B2(n_1060),
.Y(n_1413)
);

OAI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_1006),
.A2(n_951),
.B1(n_957),
.B2(n_949),
.C(n_946),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1159),
.B(n_1193),
.Y(n_1415)
);

OA22x2_ASAP7_75t_L g1416 ( 
.A1(n_1146),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1118),
.B(n_94),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1023),
.Y(n_1418)
);

AO22x2_ASAP7_75t_L g1419 ( 
.A1(n_1167),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1023),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1029),
.A2(n_957),
.B1(n_960),
.B2(n_951),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1029),
.A2(n_960),
.B1(n_965),
.B2(n_963),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1166),
.B(n_98),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1166),
.B(n_99),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1184),
.Y(n_1425)
);

AO22x2_ASAP7_75t_L g1426 ( 
.A1(n_1167),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1426)
);

AO22x2_ASAP7_75t_L g1427 ( 
.A1(n_1127),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1118),
.B(n_105),
.Y(n_1428)
);

BUFx8_ASAP7_75t_L g1429 ( 
.A(n_1118),
.Y(n_1429)
);

AO22x2_ASAP7_75t_L g1430 ( 
.A1(n_1029),
.A2(n_108),
.B1(n_105),
.B2(n_107),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1106),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1200),
.B(n_1145),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1281),
.B(n_1282),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1272),
.B(n_1145),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1224),
.B(n_1129),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1226),
.B(n_1129),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1413),
.B(n_1030),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1358),
.B(n_1094),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1223),
.B(n_1099),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1360),
.B(n_1118),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1214),
.B(n_1118),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1223),
.B(n_1099),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1240),
.B(n_1122),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1215),
.B(n_1029),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1240),
.B(n_1137),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1245),
.B(n_1137),
.Y(n_1446)
);

NAND2xp33_ASAP7_75t_SL g1447 ( 
.A(n_1417),
.B(n_1106),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1353),
.B(n_1359),
.Y(n_1448)
);

NAND2xp33_ASAP7_75t_SL g1449 ( 
.A(n_1417),
.B(n_1106),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1271),
.B(n_1186),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1381),
.B(n_1189),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1429),
.B(n_1189),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1367),
.B(n_1060),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1300),
.B(n_1176),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1295),
.B(n_1060),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1212),
.B(n_1176),
.Y(n_1456)
);

AND2x2_ASAP7_75t_SL g1457 ( 
.A(n_1428),
.B(n_1035),
.Y(n_1457)
);

NAND2xp33_ASAP7_75t_SL g1458 ( 
.A(n_1428),
.B(n_1112),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1277),
.B(n_1356),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1401),
.B(n_1060),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1235),
.B(n_1036),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1198),
.B(n_1049),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1306),
.B(n_1049),
.Y(n_1463)
);

NAND2xp33_ASAP7_75t_SL g1464 ( 
.A(n_1330),
.B(n_1081),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1262),
.B(n_1065),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1346),
.B(n_1081),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1264),
.B(n_1088),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1374),
.B(n_1108),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1297),
.B(n_1136),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1308),
.B(n_1136),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1377),
.B(n_1081),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1338),
.B(n_1149),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1415),
.B(n_1347),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1351),
.B(n_1149),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1229),
.B(n_1015),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1382),
.B(n_1081),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1284),
.B(n_1015),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1207),
.B(n_987),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1220),
.B(n_1061),
.Y(n_1479)
);

NAND2xp33_ASAP7_75t_SL g1480 ( 
.A(n_1251),
.B(n_1125),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1402),
.B(n_1125),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1241),
.B(n_1061),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1218),
.B(n_1062),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1238),
.B(n_1062),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1328),
.B(n_1077),
.Y(n_1485)
);

NAND2xp33_ASAP7_75t_SL g1486 ( 
.A(n_1391),
.B(n_1125),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1405),
.B(n_1125),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1303),
.B(n_1012),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1287),
.B(n_1125),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1303),
.B(n_1020),
.Y(n_1490)
);

NAND2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1399),
.B(n_1028),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1278),
.B(n_1028),
.Y(n_1492)
);

NAND2xp33_ASAP7_75t_R g1493 ( 
.A(n_1239),
.B(n_109),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1278),
.B(n_1028),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1202),
.B(n_1028),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1370),
.B(n_1034),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1409),
.B(n_1028),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1317),
.B(n_110),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1289),
.B(n_1312),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1410),
.B(n_1037),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1295),
.B(n_1076),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1217),
.B(n_1086),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1222),
.B(n_1192),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1216),
.B(n_110),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1225),
.B(n_112),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1232),
.B(n_1174),
.Y(n_1506)
);

NAND2xp33_ASAP7_75t_SL g1507 ( 
.A(n_1372),
.B(n_1263),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1340),
.B(n_1194),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1340),
.B(n_1175),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1233),
.B(n_113),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1305),
.B(n_1175),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1234),
.B(n_113),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1237),
.B(n_114),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1397),
.B(n_114),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1242),
.B(n_115),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1408),
.B(n_1188),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1408),
.B(n_1181),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1244),
.B(n_116),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1216),
.B(n_117),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1247),
.B(n_117),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1208),
.B(n_118),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1231),
.B(n_118),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1246),
.B(n_1182),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1320),
.B(n_119),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1248),
.B(n_120),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1203),
.B(n_1185),
.Y(n_1526)
);

NAND2xp33_ASAP7_75t_SL g1527 ( 
.A(n_1425),
.B(n_1170),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1394),
.B(n_120),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1211),
.B(n_1283),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1219),
.B(n_1279),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1279),
.B(n_980),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1418),
.B(n_1420),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1211),
.B(n_121),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1221),
.B(n_977),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1316),
.B(n_1335),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1299),
.B(n_121),
.Y(n_1536)
);

NAND2xp33_ASAP7_75t_SL g1537 ( 
.A(n_1423),
.B(n_122),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1249),
.B(n_122),
.Y(n_1538)
);

AND2x2_ASAP7_75t_SL g1539 ( 
.A(n_1213),
.B(n_124),
.Y(n_1539)
);

NAND2xp33_ASAP7_75t_SL g1540 ( 
.A(n_1424),
.B(n_124),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1252),
.B(n_125),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1253),
.B(n_1254),
.Y(n_1542)
);

NAND2xp33_ASAP7_75t_SL g1543 ( 
.A(n_1318),
.B(n_125),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1255),
.B(n_126),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1259),
.B(n_127),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1260),
.B(n_128),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_SL g1547 ( 
.A(n_1318),
.B(n_128),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1257),
.B(n_1261),
.Y(n_1548)
);

NAND2xp33_ASAP7_75t_SL g1549 ( 
.A(n_1336),
.B(n_129),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1411),
.B(n_1280),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1265),
.B(n_130),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1299),
.B(n_131),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1268),
.B(n_132),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1309),
.B(n_134),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1397),
.B(n_137),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1273),
.B(n_137),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1362),
.B(n_139),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1395),
.B(n_140),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1365),
.B(n_142),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1368),
.B(n_142),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1327),
.B(n_143),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1196),
.B(n_1366),
.Y(n_1562)
);

NAND2xp33_ASAP7_75t_SL g1563 ( 
.A(n_1431),
.B(n_143),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1205),
.B(n_144),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1236),
.B(n_144),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1332),
.B(n_145),
.Y(n_1566)
);

NAND2xp33_ASAP7_75t_SL g1567 ( 
.A(n_1431),
.B(n_145),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_SL g1568 ( 
.A(n_1293),
.B(n_146),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1379),
.B(n_147),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1339),
.B(n_148),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1311),
.B(n_149),
.Y(n_1571)
);

NAND2xp33_ASAP7_75t_SL g1572 ( 
.A(n_1296),
.B(n_151),
.Y(n_1572)
);

NAND2xp33_ASAP7_75t_SL g1573 ( 
.A(n_1384),
.B(n_153),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1275),
.B(n_153),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1315),
.B(n_154),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1292),
.B(n_155),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1344),
.B(n_156),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_SL g1578 ( 
.A(n_1369),
.B(n_156),
.Y(n_1578)
);

NAND2xp33_ASAP7_75t_SL g1579 ( 
.A(n_1371),
.B(n_157),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1345),
.B(n_158),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1349),
.B(n_160),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1298),
.B(n_160),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1342),
.B(n_161),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1389),
.B(n_161),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1390),
.B(n_164),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1392),
.B(n_164),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1393),
.B(n_166),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1421),
.B(n_166),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1315),
.B(n_170),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1343),
.B(n_170),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1380),
.B(n_171),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1383),
.B(n_172),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1387),
.B(n_173),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1388),
.B(n_174),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1348),
.B(n_175),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1199),
.B(n_176),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1352),
.B(n_177),
.Y(n_1597)
);

NAND2xp33_ASAP7_75t_SL g1598 ( 
.A(n_1319),
.B(n_179),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1286),
.B(n_181),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1206),
.B(n_181),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1355),
.B(n_182),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1227),
.B(n_183),
.Y(n_1602)
);

NAND2xp33_ASAP7_75t_SL g1603 ( 
.A(n_1321),
.B(n_184),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1197),
.B(n_1199),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1197),
.B(n_185),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1243),
.B(n_188),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1422),
.B(n_190),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1404),
.B(n_192),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1412),
.B(n_192),
.Y(n_1609)
);

NAND2xp33_ASAP7_75t_SL g1610 ( 
.A(n_1322),
.B(n_193),
.Y(n_1610)
);

NAND2xp33_ASAP7_75t_SL g1611 ( 
.A(n_1326),
.B(n_1301),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1201),
.B(n_194),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1288),
.B(n_196),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1270),
.B(n_196),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1290),
.B(n_197),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1291),
.B(n_197),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1302),
.B(n_198),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1270),
.B(n_198),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1310),
.B(n_1341),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1329),
.B(n_199),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1331),
.B(n_199),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1333),
.B(n_200),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1334),
.B(n_201),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1274),
.B(n_201),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_SL g1625 ( 
.A(n_1373),
.B(n_202),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1416),
.B(n_203),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1325),
.B(n_206),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1210),
.B(n_208),
.Y(n_1628)
);

NAND2xp33_ASAP7_75t_SL g1629 ( 
.A(n_1341),
.B(n_208),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1350),
.B(n_209),
.Y(n_1630)
);

NAND2xp33_ASAP7_75t_SL g1631 ( 
.A(n_1350),
.B(n_209),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1256),
.B(n_210),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1204),
.B(n_210),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1204),
.B(n_211),
.Y(n_1634)
);

NAND2xp33_ASAP7_75t_SL g1635 ( 
.A(n_1430),
.B(n_211),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1209),
.B(n_212),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1274),
.B(n_212),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1385),
.B(n_213),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1406),
.B(n_214),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1267),
.B(n_1269),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1430),
.B(n_214),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1398),
.B(n_1400),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1398),
.B(n_215),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1400),
.B(n_215),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1403),
.B(n_216),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1403),
.B(n_216),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1250),
.B(n_217),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1250),
.B(n_219),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1258),
.B(n_220),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1258),
.B(n_221),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1294),
.B(n_222),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1294),
.B(n_224),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1324),
.B(n_224),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1407),
.B(n_227),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1337),
.B(n_228),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1354),
.B(n_229),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1407),
.B(n_230),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1354),
.B(n_232),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1357),
.B(n_233),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1357),
.B(n_233),
.Y(n_1660)
);

NAND2xp33_ASAP7_75t_SL g1661 ( 
.A(n_1361),
.B(n_234),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1276),
.B(n_234),
.Y(n_1662)
);

NAND2xp33_ASAP7_75t_SL g1663 ( 
.A(n_1361),
.B(n_235),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1396),
.B(n_1285),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1276),
.B(n_1363),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1363),
.B(n_1285),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1396),
.B(n_236),
.Y(n_1667)
);

NAND2xp33_ASAP7_75t_SL g1668 ( 
.A(n_1304),
.B(n_236),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_SL g1669 ( 
.A(n_1304),
.B(n_237),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1307),
.B(n_238),
.Y(n_1670)
);

NAND2xp33_ASAP7_75t_SL g1671 ( 
.A(n_1313),
.B(n_239),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1313),
.B(n_239),
.Y(n_1672)
);

NAND2xp33_ASAP7_75t_SL g1673 ( 
.A(n_1314),
.B(n_240),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1314),
.B(n_240),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1228),
.B(n_241),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1228),
.B(n_241),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1230),
.B(n_242),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1419),
.B(n_243),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1419),
.B(n_244),
.Y(n_1679)
);

NAND2xp33_ASAP7_75t_SL g1680 ( 
.A(n_1427),
.B(n_246),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1426),
.B(n_246),
.Y(n_1681)
);

NAND2xp33_ASAP7_75t_SL g1682 ( 
.A(n_1427),
.B(n_247),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1323),
.B(n_247),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1266),
.B(n_248),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1266),
.B(n_248),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1414),
.B(n_249),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1386),
.B(n_250),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_SL g1688 ( 
.A(n_1364),
.B(n_1376),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1386),
.B(n_250),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1455),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1527),
.A2(n_1375),
.B(n_1376),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1437),
.A2(n_1375),
.B(n_1378),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1448),
.B(n_252),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1475),
.B(n_1378),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1455),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1657),
.B(n_253),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1571),
.A2(n_254),
.B(n_255),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1433),
.B(n_255),
.Y(n_1698)
);

BUFx12f_ASAP7_75t_L g1699 ( 
.A(n_1514),
.Y(n_1699)
);

NAND3x1_ASAP7_75t_L g1700 ( 
.A(n_1536),
.B(n_257),
.C(n_262),
.Y(n_1700)
);

AO31x2_ASAP7_75t_L g1701 ( 
.A1(n_1612),
.A2(n_265),
.A3(n_267),
.B(n_268),
.Y(n_1701)
);

NAND3x1_ASAP7_75t_L g1702 ( 
.A(n_1552),
.B(n_270),
.C(n_272),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1548),
.A2(n_277),
.B(n_278),
.Y(n_1703)
);

AO21x2_ASAP7_75t_L g1704 ( 
.A1(n_1642),
.A2(n_279),
.B(n_284),
.Y(n_1704)
);

NAND3xp33_ASAP7_75t_L g1705 ( 
.A(n_1688),
.B(n_286),
.C(n_288),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1464),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1641),
.A2(n_293),
.B(n_295),
.Y(n_1707)
);

INVx3_ASAP7_75t_SL g1708 ( 
.A(n_1530),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1538),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1641),
.A2(n_1637),
.B1(n_1657),
.B2(n_1457),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1542),
.B(n_299),
.Y(n_1711)
);

INVx6_ASAP7_75t_L g1712 ( 
.A(n_1637),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1462),
.B(n_1529),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1481),
.A2(n_1487),
.B(n_1497),
.Y(n_1714)
);

INVxp67_ASAP7_75t_SL g1715 ( 
.A(n_1538),
.Y(n_1715)
);

A2O1A1Ixp33_ASAP7_75t_L g1716 ( 
.A1(n_1688),
.A2(n_303),
.B(n_304),
.C(n_306),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1493),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1661),
.A2(n_314),
.B(n_317),
.C(n_319),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1447),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1555),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1664),
.B(n_428),
.Y(n_1721)
);

CKINVDCx14_ASAP7_75t_R g1722 ( 
.A(n_1657),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1538),
.Y(n_1723)
);

NOR4xp25_ASAP7_75t_L g1724 ( 
.A(n_1666),
.B(n_328),
.C(n_331),
.D(n_332),
.Y(n_1724)
);

BUFx3_ASAP7_75t_L g1725 ( 
.A(n_1541),
.Y(n_1725)
);

INVx4_ASAP7_75t_L g1726 ( 
.A(n_1455),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1641),
.A2(n_338),
.B1(n_339),
.B2(n_341),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_L g1728 ( 
.A(n_1680),
.B(n_343),
.C(n_344),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1541),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1637),
.A2(n_346),
.B1(n_348),
.B2(n_349),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1539),
.B(n_352),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1457),
.A2(n_353),
.B1(n_359),
.B2(n_361),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1539),
.B(n_1629),
.Y(n_1733)
);

AO32x2_ASAP7_75t_L g1734 ( 
.A1(n_1680),
.A2(n_362),
.A3(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_1734)
);

AOI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1668),
.A2(n_1669),
.B1(n_1673),
.B2(n_1671),
.C(n_1456),
.Y(n_1735)
);

BUFx4_ASAP7_75t_SL g1736 ( 
.A(n_1686),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1473),
.B(n_384),
.Y(n_1737)
);

AO32x2_ASAP7_75t_L g1738 ( 
.A1(n_1682),
.A2(n_387),
.A3(n_388),
.B1(n_390),
.B2(n_392),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1665),
.A2(n_393),
.B1(n_398),
.B2(n_399),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1541),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1522),
.B(n_403),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1459),
.B(n_405),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1654),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1467),
.B(n_423),
.Y(n_1744)
);

NAND2x1p5_ASAP7_75t_L g1745 ( 
.A(n_1508),
.B(n_413),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1438),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1544),
.Y(n_1747)
);

BUFx12f_ASAP7_75t_L g1748 ( 
.A(n_1544),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1544),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1434),
.B(n_415),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1438),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1466),
.A2(n_417),
.B1(n_418),
.B2(n_420),
.Y(n_1752)
);

BUFx2_ASAP7_75t_R g1753 ( 
.A(n_1662),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1575),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1617),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1499),
.B(n_421),
.Y(n_1756)
);

AO21x1_ASAP7_75t_L g1757 ( 
.A1(n_1682),
.A2(n_1635),
.B(n_1663),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1599),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1477),
.B(n_1474),
.Y(n_1759)
);

OAI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1640),
.A2(n_1440),
.B(n_1471),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1617),
.Y(n_1761)
);

AO31x2_ASAP7_75t_L g1762 ( 
.A1(n_1687),
.A2(n_1689),
.A3(n_1681),
.B(n_1660),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1589),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1684),
.A2(n_1535),
.B1(n_1617),
.B2(n_1599),
.Y(n_1764)
);

NAND2xp33_ASAP7_75t_L g1765 ( 
.A(n_1447),
.B(n_1449),
.Y(n_1765)
);

OAI21x1_ASAP7_75t_SL g1766 ( 
.A1(n_1677),
.A2(n_1667),
.B(n_1476),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1498),
.B(n_1524),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_SL g1768 ( 
.A(n_1684),
.B(n_1599),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1769)
);

BUFx2_ASAP7_75t_SL g1770 ( 
.A(n_1684),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1494),
.B(n_1554),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1449),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1521),
.B(n_1528),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1639),
.A2(n_1500),
.B(n_1638),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1626),
.A2(n_1672),
.B(n_1674),
.C(n_1670),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1517),
.B(n_1450),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1480),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1469),
.B(n_1470),
.Y(n_1778)
);

INVx3_ASAP7_75t_L g1779 ( 
.A(n_1438),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1505),
.Y(n_1780)
);

OAI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1453),
.A2(n_1460),
.B1(n_1441),
.B2(n_1511),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1502),
.Y(n_1782)
);

AOI211x1_ASAP7_75t_L g1783 ( 
.A1(n_1675),
.A2(n_1676),
.B(n_1679),
.C(n_1678),
.Y(n_1783)
);

A2O1A1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1668),
.A2(n_1671),
.B(n_1673),
.C(n_1669),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1452),
.B(n_1451),
.Y(n_1785)
);

AOI221x1_ASAP7_75t_L g1786 ( 
.A1(n_1635),
.A2(n_1549),
.B1(n_1543),
.B2(n_1547),
.C(n_1572),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1472),
.B(n_1495),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1435),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1510),
.A2(n_1513),
.B(n_1512),
.Y(n_1789)
);

O2A1O1Ixp5_ASAP7_75t_L g1790 ( 
.A1(n_1507),
.A2(n_1607),
.B(n_1609),
.C(n_1629),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1461),
.B(n_1463),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1443),
.B(n_1445),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1614),
.B(n_1618),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1624),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1436),
.B(n_1515),
.Y(n_1795)
);

BUFx10_ASAP7_75t_L g1796 ( 
.A(n_1619),
.Y(n_1796)
);

AO22x2_ASAP7_75t_L g1797 ( 
.A1(n_1647),
.A2(n_1648),
.B1(n_1649),
.B2(n_1650),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1458),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1444),
.A2(n_1516),
.B1(n_1533),
.B2(n_1636),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1506),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1506),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1518),
.B(n_1520),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1525),
.B(n_1545),
.Y(n_1803)
);

INVx3_ASAP7_75t_L g1804 ( 
.A(n_1501),
.Y(n_1804)
);

AOI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1651),
.A2(n_1653),
.B(n_1652),
.Y(n_1805)
);

CKINVDCx16_ASAP7_75t_R g1806 ( 
.A(n_1504),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1546),
.Y(n_1807)
);

INVx4_ASAP7_75t_L g1808 ( 
.A(n_1501),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1551),
.B(n_1553),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1432),
.B(n_1488),
.Y(n_1810)
);

NAND3x1_ASAP7_75t_L g1811 ( 
.A(n_1519),
.B(n_1596),
.C(n_1683),
.Y(n_1811)
);

OAI22x1_ASAP7_75t_L g1812 ( 
.A1(n_1633),
.A2(n_1634),
.B1(n_1645),
.B2(n_1646),
.Y(n_1812)
);

OR2x6_ASAP7_75t_L g1813 ( 
.A(n_1490),
.B(n_1509),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1458),
.A2(n_1507),
.B(n_1468),
.Y(n_1814)
);

NOR2xp67_ASAP7_75t_L g1815 ( 
.A(n_1628),
.B(n_1643),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1561),
.B(n_1446),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1631),
.B(n_1619),
.Y(n_1817)
);

INVx5_ASAP7_75t_L g1818 ( 
.A(n_1619),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1506),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1627),
.B(n_1655),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1656),
.A2(n_1659),
.B1(n_1658),
.B2(n_1685),
.C(n_1644),
.Y(n_1821)
);

OAI21x1_ASAP7_75t_L g1822 ( 
.A1(n_1600),
.A2(n_1602),
.B(n_1606),
.Y(n_1822)
);

NOR2xp67_ASAP7_75t_L g1823 ( 
.A(n_1630),
.B(n_1582),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1583),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1590),
.Y(n_1825)
);

AO31x2_ASAP7_75t_L g1826 ( 
.A1(n_1595),
.A2(n_1597),
.A3(n_1601),
.B(n_1503),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1465),
.A2(n_1454),
.B(n_1565),
.Y(n_1827)
);

OAI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1632),
.A2(n_1523),
.B(n_1550),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1439),
.B(n_1442),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1556),
.B(n_1478),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1557),
.A2(n_1558),
.B1(n_1482),
.B2(n_1559),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1588),
.A2(n_1526),
.B(n_1479),
.Y(n_1832)
);

A2O1A1Ixp33_ASAP7_75t_L g1833 ( 
.A1(n_1598),
.A2(n_1603),
.B(n_1610),
.C(n_1540),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1562),
.B(n_1608),
.Y(n_1834)
);

INVx5_ASAP7_75t_L g1835 ( 
.A(n_1603),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1560),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1563),
.Y(n_1837)
);

A2O1A1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1537),
.A2(n_1540),
.B(n_1579),
.C(n_1578),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1574),
.B(n_1576),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1537),
.B(n_1613),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1615),
.B(n_1616),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1577),
.A2(n_1580),
.B(n_1581),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1483),
.A2(n_1484),
.B(n_1586),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1566),
.Y(n_1844)
);

NAND2xp33_ASAP7_75t_R g1845 ( 
.A(n_1578),
.B(n_1579),
.Y(n_1845)
);

OAI22x1_ASAP7_75t_L g1846 ( 
.A1(n_1570),
.A2(n_1531),
.B1(n_1564),
.B2(n_1569),
.Y(n_1846)
);

AO32x2_ASAP7_75t_L g1847 ( 
.A1(n_1568),
.A2(n_1573),
.A3(n_1563),
.B1(n_1567),
.B2(n_1625),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1620),
.Y(n_1848)
);

O2A1O1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1584),
.A2(n_1585),
.B(n_1587),
.C(n_1623),
.Y(n_1849)
);

AOI211x1_ASAP7_75t_L g1850 ( 
.A1(n_1621),
.A2(n_1622),
.B(n_1591),
.C(n_1592),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1573),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1611),
.A2(n_1486),
.B(n_1491),
.C(n_1532),
.Y(n_1852)
);

BUFx12f_ASAP7_75t_L g1853 ( 
.A(n_1496),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1534),
.Y(n_1854)
);

OAI21x1_ASAP7_75t_L g1855 ( 
.A1(n_1594),
.A2(n_1593),
.B(n_1485),
.Y(n_1855)
);

NOR2xp67_ASAP7_75t_SL g1856 ( 
.A(n_1530),
.B(n_1017),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1475),
.B(n_1448),
.Y(n_1857)
);

AO31x2_ASAP7_75t_L g1858 ( 
.A1(n_1604),
.A2(n_1161),
.A3(n_1612),
.B(n_1605),
.Y(n_1858)
);

OAI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1571),
.A2(n_1263),
.B(n_1377),
.Y(n_1859)
);

AO22x2_ASAP7_75t_L g1860 ( 
.A1(n_1666),
.A2(n_1642),
.B1(n_1665),
.B2(n_1637),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1475),
.B(n_1448),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1448),
.B(n_1003),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1475),
.B(n_1448),
.Y(n_1863)
);

O2A1O1Ixp5_ASAP7_75t_L g1864 ( 
.A1(n_1639),
.A2(n_1507),
.B(n_1688),
.C(n_1642),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1448),
.B(n_1003),
.Y(n_1865)
);

INVx4_ASAP7_75t_SL g1866 ( 
.A(n_1637),
.Y(n_1866)
);

OAI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1462),
.A2(n_1401),
.B(n_1367),
.Y(n_1867)
);

AO31x2_ASAP7_75t_L g1868 ( 
.A1(n_1604),
.A2(n_1161),
.A3(n_1612),
.B(n_1605),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1538),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1539),
.B(n_1083),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1475),
.B(n_1448),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1455),
.B(n_1433),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1475),
.B(n_1448),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1455),
.Y(n_1874)
);

BUFx3_ASAP7_75t_L g1875 ( 
.A(n_1555),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1455),
.B(n_1433),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1782),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1757),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1857),
.B(n_1861),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_L g1880 ( 
.A(n_1806),
.B(n_1754),
.Y(n_1880)
);

OAI21x1_ASAP7_75t_SL g1881 ( 
.A1(n_1710),
.A2(n_1764),
.B(n_1735),
.Y(n_1881)
);

AO21x2_ASAP7_75t_L g1882 ( 
.A1(n_1691),
.A2(n_1766),
.B(n_1814),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1770),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1851),
.Y(n_1884)
);

NOR2x1_ASAP7_75t_L g1885 ( 
.A(n_1813),
.B(n_1707),
.Y(n_1885)
);

INVx6_ASAP7_75t_L g1886 ( 
.A(n_1796),
.Y(n_1886)
);

AO21x2_ASAP7_75t_L g1887 ( 
.A1(n_1833),
.A2(n_1838),
.B(n_1827),
.Y(n_1887)
);

BUFx4f_ASAP7_75t_L g1888 ( 
.A(n_1708),
.Y(n_1888)
);

AOI222xp33_ASAP7_75t_L g1889 ( 
.A1(n_1866),
.A2(n_1871),
.B1(n_1863),
.B2(n_1873),
.C1(n_1867),
.C2(n_1793),
.Y(n_1889)
);

BUFx10_ASAP7_75t_L g1890 ( 
.A(n_1785),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1862),
.B(n_1865),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1763),
.B(n_1743),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1722),
.A2(n_1712),
.B1(n_1715),
.B2(n_1748),
.Y(n_1893)
);

A2O1A1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1768),
.A2(n_1784),
.B(n_1775),
.C(n_1733),
.Y(n_1894)
);

AO21x2_ASAP7_75t_L g1895 ( 
.A1(n_1827),
.A2(n_1692),
.B(n_1843),
.Y(n_1895)
);

NAND2x1p5_ASAP7_75t_L g1896 ( 
.A(n_1856),
.B(n_1818),
.Y(n_1896)
);

AO32x2_ASAP7_75t_L g1897 ( 
.A1(n_1799),
.A2(n_1831),
.A3(n_1730),
.B1(n_1727),
.B2(n_1860),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1794),
.B(n_1693),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_SL g1899 ( 
.A1(n_1768),
.A2(n_1712),
.B1(n_1860),
.B2(n_1696),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1725),
.A2(n_1729),
.B1(n_1749),
.B2(n_1758),
.Y(n_1900)
);

AOI221xp5_ASAP7_75t_SL g1901 ( 
.A1(n_1870),
.A2(n_1812),
.B1(n_1713),
.B2(n_1820),
.C(n_1767),
.Y(n_1901)
);

AO32x2_ASAP7_75t_L g1902 ( 
.A1(n_1781),
.A2(n_1732),
.A3(n_1762),
.B1(n_1808),
.B2(n_1858),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1759),
.B(n_1872),
.Y(n_1903)
);

AO32x2_ASAP7_75t_L g1904 ( 
.A1(n_1762),
.A2(n_1808),
.A3(n_1858),
.B1(n_1868),
.B2(n_1783),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1720),
.B(n_1875),
.Y(n_1905)
);

CKINVDCx16_ASAP7_75t_R g1906 ( 
.A(n_1699),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1876),
.B(n_1726),
.Y(n_1907)
);

BUFx2_ASAP7_75t_L g1908 ( 
.A(n_1853),
.Y(n_1908)
);

AO21x2_ASAP7_75t_L g1909 ( 
.A1(n_1805),
.A2(n_1705),
.B(n_1815),
.Y(n_1909)
);

OA21x2_ASAP7_75t_L g1910 ( 
.A1(n_1786),
.A2(n_1864),
.B(n_1821),
.Y(n_1910)
);

OAI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1859),
.A2(n_1774),
.B(n_1789),
.Y(n_1911)
);

OAI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1717),
.A2(n_1835),
.B1(n_1845),
.B2(n_1837),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1751),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1709),
.Y(n_1914)
);

INVx4_ASAP7_75t_L g1915 ( 
.A(n_1818),
.Y(n_1915)
);

BUFx12f_ASAP7_75t_L g1916 ( 
.A(n_1785),
.Y(n_1916)
);

A2O1A1Ixp33_ASAP7_75t_L g1917 ( 
.A1(n_1815),
.A2(n_1837),
.B(n_1731),
.C(n_1821),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1876),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1723),
.Y(n_1919)
);

BUFx8_ASAP7_75t_L g1920 ( 
.A(n_1777),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1797),
.A2(n_1780),
.B1(n_1807),
.B2(n_1824),
.Y(n_1921)
);

NAND3xp33_ASAP7_75t_L g1922 ( 
.A(n_1783),
.B(n_1850),
.C(n_1697),
.Y(n_1922)
);

AO31x2_ASAP7_75t_L g1923 ( 
.A1(n_1852),
.A2(n_1694),
.A3(n_1716),
.B(n_1718),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1726),
.B(n_1746),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1774),
.A2(n_1789),
.B(n_1802),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1695),
.B(n_1874),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1771),
.B(n_1769),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_SL g1928 ( 
.A(n_1753),
.B(n_1835),
.Y(n_1928)
);

OAI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1803),
.A2(n_1809),
.B(n_1790),
.Y(n_1929)
);

AOI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1825),
.A2(n_1797),
.B1(n_1697),
.B2(n_1773),
.C(n_1791),
.Y(n_1930)
);

O2A1O1Ixp33_ASAP7_75t_L g1931 ( 
.A1(n_1840),
.A2(n_1778),
.B(n_1834),
.C(n_1839),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1835),
.A2(n_1811),
.B1(n_1869),
.B2(n_1740),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1747),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1698),
.Y(n_1934)
);

AOI222xp33_ASAP7_75t_L g1935 ( 
.A1(n_1817),
.A2(n_1816),
.B1(n_1787),
.B2(n_1810),
.C1(n_1736),
.C2(n_1776),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1746),
.B(n_1779),
.Y(n_1936)
);

AOI21xp33_ASAP7_75t_L g1937 ( 
.A1(n_1849),
.A2(n_1846),
.B(n_1841),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1779),
.B(n_1818),
.Y(n_1938)
);

INVxp33_ASAP7_75t_L g1939 ( 
.A(n_1751),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1844),
.A2(n_1836),
.B1(n_1761),
.B2(n_1755),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1690),
.B(n_1751),
.Y(n_1941)
);

NAND2x1p5_ASAP7_75t_L g1942 ( 
.A(n_1810),
.B(n_1690),
.Y(n_1942)
);

INVxp33_ASAP7_75t_L g1943 ( 
.A(n_1695),
.Y(n_1943)
);

A2O1A1Ixp33_ASAP7_75t_L g1944 ( 
.A1(n_1728),
.A2(n_1739),
.B(n_1823),
.C(n_1706),
.Y(n_1944)
);

OA21x2_ASAP7_75t_L g1945 ( 
.A1(n_1760),
.A2(n_1832),
.B(n_1714),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1760),
.A2(n_1828),
.B(n_1823),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1695),
.B(n_1874),
.Y(n_1947)
);

BUFx12f_ASAP7_75t_L g1948 ( 
.A(n_1813),
.Y(n_1948)
);

BUFx2_ASAP7_75t_R g1949 ( 
.A(n_1721),
.Y(n_1949)
);

CKINVDCx20_ASAP7_75t_R g1950 ( 
.A(n_1796),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1742),
.B(n_1874),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1788),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1792),
.B(n_1829),
.Y(n_1953)
);

OAI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1828),
.A2(n_1795),
.B(n_1830),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1700),
.A2(n_1739),
.B1(n_1702),
.B2(n_1772),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1762),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1800),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_SL g1958 ( 
.A1(n_1765),
.A2(n_1798),
.B1(n_1772),
.B2(n_1719),
.Y(n_1958)
);

OA21x2_ASAP7_75t_L g1959 ( 
.A1(n_1714),
.A2(n_1703),
.B(n_1842),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_1804),
.Y(n_1960)
);

OAI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1822),
.A2(n_1855),
.B(n_1848),
.Y(n_1961)
);

INVx2_ASAP7_75t_SL g1962 ( 
.A(n_1801),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1819),
.B(n_1711),
.Y(n_1963)
);

OAI21x1_ASAP7_75t_L g1964 ( 
.A1(n_1756),
.A2(n_1744),
.B(n_1745),
.Y(n_1964)
);

BUFx3_ASAP7_75t_L g1965 ( 
.A(n_1854),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1750),
.B(n_1737),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1826),
.B(n_1850),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1826),
.B(n_1868),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1719),
.B(n_1798),
.Y(n_1969)
);

OA21x2_ASAP7_75t_L g1970 ( 
.A1(n_1741),
.A2(n_1752),
.B(n_1847),
.Y(n_1970)
);

CKINVDCx20_ASAP7_75t_R g1971 ( 
.A(n_1704),
.Y(n_1971)
);

OA21x2_ASAP7_75t_L g1972 ( 
.A1(n_1724),
.A2(n_1701),
.B(n_1734),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1826),
.B(n_1701),
.Y(n_1973)
);

AOI22xp33_ASAP7_75t_L g1974 ( 
.A1(n_1738),
.A2(n_1666),
.B1(n_1710),
.B2(n_1637),
.Y(n_1974)
);

INVx2_ASAP7_75t_SL g1975 ( 
.A(n_1738),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1857),
.B(n_1861),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1806),
.B(n_893),
.Y(n_1977)
);

NOR2x1p5_ASAP7_75t_L g1978 ( 
.A(n_1748),
.B(n_1042),
.Y(n_1978)
);

NOR2xp67_ASAP7_75t_L g1979 ( 
.A(n_1710),
.B(n_1530),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1866),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1866),
.B(n_1872),
.Y(n_1981)
);

NAND3xp33_ASAP7_75t_L g1982 ( 
.A(n_1735),
.B(n_1669),
.C(n_1668),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1857),
.B(n_1861),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1782),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1866),
.B(n_1768),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1857),
.B(n_1861),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1884),
.Y(n_1987)
);

NAND2x1p5_ASAP7_75t_L g1988 ( 
.A(n_1985),
.B(n_1885),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1967),
.B(n_1891),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1884),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1914),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1878),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1878),
.B(n_1887),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1879),
.B(n_1976),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1887),
.B(n_1956),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1980),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1913),
.Y(n_1997)
);

BUFx2_ASAP7_75t_L g1998 ( 
.A(n_1969),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1956),
.B(n_1919),
.Y(n_1999)
);

NAND2x1p5_ASAP7_75t_L g2000 ( 
.A(n_1981),
.B(n_1915),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1950),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1933),
.B(n_1911),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1975),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1968),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1904),
.Y(n_2005)
);

OAI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1929),
.A2(n_1925),
.B(n_1982),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_SL g2007 ( 
.A1(n_1928),
.A2(n_1881),
.B1(n_1955),
.B2(n_1948),
.Y(n_2007)
);

INVx3_ASAP7_75t_L g2008 ( 
.A(n_1981),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1913),
.Y(n_2009)
);

INVx3_ASAP7_75t_SL g2010 ( 
.A(n_1886),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_1886),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1927),
.B(n_1921),
.Y(n_2012)
);

BUFx3_ASAP7_75t_L g2013 ( 
.A(n_1888),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1952),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_1908),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1877),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1915),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1904),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1889),
.A2(n_1935),
.B1(n_1979),
.B2(n_1930),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1974),
.B(n_1945),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1984),
.B(n_1899),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1977),
.B(n_1898),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1973),
.Y(n_2023)
);

CKINVDCx16_ASAP7_75t_R g2024 ( 
.A(n_1906),
.Y(n_2024)
);

AND2x4_ASAP7_75t_L g2025 ( 
.A(n_1894),
.B(n_1961),
.Y(n_2025)
);

BUFx10_ASAP7_75t_L g2026 ( 
.A(n_1978),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_SL g2027 ( 
.A1(n_1893),
.A2(n_1920),
.B1(n_1916),
.B2(n_1890),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1983),
.B(n_1986),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1957),
.B(n_1897),
.Y(n_2029)
);

CKINVDCx6p67_ASAP7_75t_R g2030 ( 
.A(n_1890),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1892),
.B(n_1905),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1897),
.B(n_1895),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1897),
.B(n_1918),
.Y(n_2033)
);

NOR2x1p5_ASAP7_75t_L g2034 ( 
.A(n_1922),
.B(n_1883),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1882),
.Y(n_2035)
);

INVxp67_ASAP7_75t_L g2036 ( 
.A(n_1880),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1910),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1910),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1953),
.B(n_1934),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1972),
.Y(n_2040)
);

BUFx3_ASAP7_75t_L g2041 ( 
.A(n_1888),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1883),
.Y(n_2042)
);

OAI221xp5_ASAP7_75t_L g2043 ( 
.A1(n_1901),
.A2(n_1937),
.B1(n_1946),
.B2(n_1944),
.C(n_1966),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_SL g2044 ( 
.A1(n_1920),
.A2(n_1907),
.B1(n_1971),
.B2(n_1972),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1903),
.B(n_1931),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_1907),
.A2(n_1951),
.B1(n_1936),
.B2(n_1965),
.Y(n_2046)
);

BUFx24_ASAP7_75t_SL g2047 ( 
.A(n_2027),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2014),
.B(n_1926),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_SL g2049 ( 
.A(n_2010),
.B(n_1932),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1989),
.B(n_1940),
.Y(n_2050)
);

INVx1_ASAP7_75t_SL g2051 ( 
.A(n_2015),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2042),
.B(n_1939),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_1998),
.B(n_1947),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_2024),
.Y(n_2054)
);

NAND2xp33_ASAP7_75t_R g2055 ( 
.A(n_2017),
.B(n_1938),
.Y(n_2055)
);

XNOR2xp5_ASAP7_75t_L g2056 ( 
.A(n_2001),
.B(n_1912),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_2001),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_1996),
.Y(n_2058)
);

NAND2xp33_ASAP7_75t_R g2059 ( 
.A(n_2017),
.B(n_1924),
.Y(n_2059)
);

NAND2xp33_ASAP7_75t_R g2060 ( 
.A(n_2017),
.B(n_2008),
.Y(n_2060)
);

CKINVDCx11_ASAP7_75t_R g2061 ( 
.A(n_2026),
.Y(n_2061)
);

NAND2xp33_ASAP7_75t_R g2062 ( 
.A(n_2008),
.B(n_1924),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2031),
.B(n_1941),
.Y(n_2063)
);

NAND2xp33_ASAP7_75t_R g2064 ( 
.A(n_2008),
.B(n_1994),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_2023),
.B(n_1917),
.Y(n_2065)
);

BUFx10_ASAP7_75t_L g2066 ( 
.A(n_2011),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_2026),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1989),
.B(n_2002),
.Y(n_2068)
);

NAND2xp33_ASAP7_75t_R g2069 ( 
.A(n_2028),
.B(n_1970),
.Y(n_2069)
);

INVxp67_ASAP7_75t_L g2070 ( 
.A(n_2039),
.Y(n_2070)
);

NAND2xp33_ASAP7_75t_SL g2071 ( 
.A(n_2010),
.B(n_1960),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_2036),
.B(n_1949),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2002),
.B(n_1954),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2012),
.B(n_1962),
.Y(n_2074)
);

OR2x6_ASAP7_75t_L g2075 ( 
.A(n_2013),
.B(n_1896),
.Y(n_2075)
);

NAND2xp33_ASAP7_75t_R g2076 ( 
.A(n_2033),
.B(n_1970),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_2013),
.Y(n_2077)
);

OR2x6_ASAP7_75t_L g2078 ( 
.A(n_2041),
.B(n_1942),
.Y(n_2078)
);

NAND2xp33_ASAP7_75t_R g2079 ( 
.A(n_2033),
.B(n_1959),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1991),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_R g2081 ( 
.A(n_2041),
.B(n_1960),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_L g2082 ( 
.A(n_2022),
.B(n_1943),
.Y(n_2082)
);

BUFx3_ASAP7_75t_L g2083 ( 
.A(n_2010),
.Y(n_2083)
);

BUFx6f_ASAP7_75t_L g2084 ( 
.A(n_2030),
.Y(n_2084)
);

NAND2xp33_ASAP7_75t_R g2085 ( 
.A(n_2021),
.B(n_1959),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_1999),
.B(n_1909),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2034),
.B(n_1958),
.Y(n_2087)
);

INVxp67_ASAP7_75t_L g2088 ( 
.A(n_2011),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_R g2089 ( 
.A(n_2030),
.B(n_1963),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_2000),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2012),
.B(n_1900),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2045),
.B(n_1923),
.Y(n_2092)
);

INVxp67_ASAP7_75t_L g2093 ( 
.A(n_1997),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_1999),
.B(n_1923),
.Y(n_2094)
);

XNOR2xp5_ASAP7_75t_L g2095 ( 
.A(n_2007),
.B(n_1964),
.Y(n_2095)
);

OR2x6_ASAP7_75t_L g2096 ( 
.A(n_2000),
.B(n_1902),
.Y(n_2096)
);

NAND2xp33_ASAP7_75t_R g2097 ( 
.A(n_2029),
.B(n_2025),
.Y(n_2097)
);

CKINVDCx16_ASAP7_75t_R g2098 ( 
.A(n_2009),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2016),
.B(n_1923),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2068),
.B(n_1987),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_2086),
.B(n_1995),
.Y(n_2101)
);

AND2x4_ASAP7_75t_L g2102 ( 
.A(n_2086),
.B(n_1995),
.Y(n_2102)
);

INVxp67_ASAP7_75t_L g2103 ( 
.A(n_2059),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2094),
.B(n_2020),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_SL g2105 ( 
.A1(n_2089),
.A2(n_1988),
.B1(n_2043),
.B2(n_2032),
.Y(n_2105)
);

NAND2x1p5_ASAP7_75t_L g2106 ( 
.A(n_2090),
.B(n_2025),
.Y(n_2106)
);

OR2x2_ASAP7_75t_L g2107 ( 
.A(n_2092),
.B(n_1992),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2073),
.B(n_1987),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2096),
.B(n_1993),
.Y(n_2109)
);

OAI21xp33_ASAP7_75t_SL g2110 ( 
.A1(n_2064),
.A2(n_2019),
.B(n_2029),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_2096),
.B(n_2035),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2080),
.B(n_2003),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_2051),
.B(n_2072),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2099),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2065),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2070),
.B(n_1990),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2098),
.B(n_1990),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2050),
.B(n_1992),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2065),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2048),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2058),
.B(n_2052),
.Y(n_2121)
);

AND2x4_ASAP7_75t_L g2122 ( 
.A(n_2053),
.B(n_2035),
.Y(n_2122)
);

OR2x2_ASAP7_75t_L g2123 ( 
.A(n_2074),
.B(n_2004),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2093),
.B(n_2006),
.Y(n_2124)
);

OAI21xp33_ASAP7_75t_L g2125 ( 
.A1(n_2087),
.A2(n_2044),
.B(n_2025),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2125),
.A2(n_2047),
.B1(n_2082),
.B2(n_2063),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2104),
.B(n_2005),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2104),
.B(n_2005),
.Y(n_2128)
);

AO21x2_ASAP7_75t_L g2129 ( 
.A1(n_2124),
.A2(n_2038),
.B(n_2037),
.Y(n_2129)
);

INVx2_ASAP7_75t_SL g2130 ( 
.A(n_2122),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2114),
.Y(n_2131)
);

BUFx3_ASAP7_75t_L g2132 ( 
.A(n_2106),
.Y(n_2132)
);

NOR2x1_ASAP7_75t_SL g2133 ( 
.A(n_2109),
.B(n_2084),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_2114),
.Y(n_2134)
);

NOR2x1_ASAP7_75t_L g2135 ( 
.A(n_2111),
.B(n_2083),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2107),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_2113),
.B(n_2054),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2101),
.B(n_2018),
.Y(n_2138)
);

OR2x2_ASAP7_75t_L g2139 ( 
.A(n_2123),
.B(n_2040),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2101),
.B(n_2018),
.Y(n_2140)
);

AOI322xp5_ASAP7_75t_L g2141 ( 
.A1(n_2110),
.A2(n_2103),
.A3(n_2105),
.B1(n_2120),
.B2(n_2109),
.C1(n_2049),
.C2(n_2116),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2107),
.Y(n_2142)
);

OAI21xp33_ASAP7_75t_L g2143 ( 
.A1(n_2110),
.A2(n_2095),
.B(n_2056),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2123),
.B(n_2118),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_2112),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2136),
.B(n_2120),
.Y(n_2146)
);

HB1xp67_ASAP7_75t_L g2147 ( 
.A(n_2134),
.Y(n_2147)
);

OR2x6_ASAP7_75t_L g2148 ( 
.A(n_2135),
.B(n_2106),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2138),
.B(n_2101),
.Y(n_2149)
);

INVx4_ASAP7_75t_L g2150 ( 
.A(n_2132),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2144),
.B(n_2121),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_2144),
.B(n_2100),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2138),
.B(n_2140),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2140),
.B(n_2101),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2135),
.B(n_2111),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2134),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2131),
.Y(n_2157)
);

HB1xp67_ASAP7_75t_L g2158 ( 
.A(n_2145),
.Y(n_2158)
);

INVx3_ASAP7_75t_L g2159 ( 
.A(n_2132),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2127),
.B(n_2102),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2127),
.B(n_2102),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2129),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2131),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2129),
.Y(n_2164)
);

OR2x2_ASAP7_75t_L g2165 ( 
.A(n_2145),
.B(n_2108),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2128),
.B(n_2102),
.Y(n_2166)
);

AOI22xp33_ASAP7_75t_L g2167 ( 
.A1(n_2143),
.A2(n_2102),
.B1(n_2115),
.B2(n_2119),
.Y(n_2167)
);

NAND2xp33_ASAP7_75t_SL g2168 ( 
.A(n_2150),
.B(n_2055),
.Y(n_2168)
);

OR2x2_ASAP7_75t_L g2169 ( 
.A(n_2165),
.B(n_2139),
.Y(n_2169)
);

NOR4xp25_ASAP7_75t_SL g2170 ( 
.A(n_2156),
.B(n_2143),
.C(n_2060),
.D(n_2062),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2167),
.B(n_2136),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_L g2172 ( 
.A(n_2151),
.B(n_2137),
.Y(n_2172)
);

NOR2xp67_ASAP7_75t_L g2173 ( 
.A(n_2150),
.B(n_2130),
.Y(n_2173)
);

BUFx3_ASAP7_75t_L g2174 ( 
.A(n_2150),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2158),
.B(n_2142),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2157),
.B(n_2142),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2158),
.B(n_2141),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_2150),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_2151),
.B(n_2057),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2153),
.B(n_2141),
.Y(n_2180)
);

AOI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2149),
.A2(n_2126),
.B1(n_2097),
.B2(n_2085),
.Y(n_2181)
);

NOR2xp67_ASAP7_75t_L g2182 ( 
.A(n_2159),
.B(n_2130),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_2146),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2171),
.B(n_2149),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2169),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2176),
.Y(n_2186)
);

INVx1_ASAP7_75t_SL g2187 ( 
.A(n_2174),
.Y(n_2187)
);

INVx1_ASAP7_75t_SL g2188 ( 
.A(n_2178),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2176),
.Y(n_2189)
);

OAI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_2180),
.A2(n_2159),
.B1(n_2148),
.B2(n_2155),
.Y(n_2190)
);

INVxp33_ASAP7_75t_L g2191 ( 
.A(n_2173),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_2168),
.A2(n_2148),
.B(n_2159),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2175),
.B(n_2165),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2177),
.B(n_2156),
.Y(n_2194)
);

INVxp67_ASAP7_75t_L g2195 ( 
.A(n_2172),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_2178),
.B(n_2152),
.Y(n_2196)
);

AOI22xp33_ASAP7_75t_L g2197 ( 
.A1(n_2181),
.A2(n_2126),
.B1(n_2155),
.B2(n_2119),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2183),
.B(n_2153),
.Y(n_2198)
);

HB1xp67_ASAP7_75t_L g2199 ( 
.A(n_2182),
.Y(n_2199)
);

HB1xp67_ASAP7_75t_L g2200 ( 
.A(n_2179),
.Y(n_2200)
);

AND2x4_ASAP7_75t_L g2201 ( 
.A(n_2170),
.B(n_2155),
.Y(n_2201)
);

HB1xp67_ASAP7_75t_L g2202 ( 
.A(n_2174),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_2183),
.B(n_2061),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_2194),
.B(n_2152),
.Y(n_2204)
);

BUFx2_ASAP7_75t_L g2205 ( 
.A(n_2202),
.Y(n_2205)
);

NAND2xp33_ASAP7_75t_L g2206 ( 
.A(n_2187),
.B(n_2200),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_2195),
.A2(n_2159),
.B1(n_2155),
.B2(n_2130),
.Y(n_2207)
);

OAI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_2197),
.A2(n_2148),
.B1(n_2147),
.B2(n_2132),
.Y(n_2208)
);

AOI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_2192),
.A2(n_2148),
.B(n_2147),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2185),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2193),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2201),
.B(n_2149),
.Y(n_2212)
);

NAND4xp25_ASAP7_75t_SL g2213 ( 
.A(n_2194),
.B(n_2117),
.C(n_2166),
.D(n_2161),
.Y(n_2213)
);

OAI32xp33_ASAP7_75t_L g2214 ( 
.A1(n_2191),
.A2(n_2146),
.A3(n_2077),
.B1(n_2106),
.B2(n_2161),
.Y(n_2214)
);

OAI22xp33_ASAP7_75t_L g2215 ( 
.A1(n_2191),
.A2(n_2148),
.B1(n_2084),
.B2(n_2139),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_SL g2216 ( 
.A(n_2201),
.B(n_2084),
.Y(n_2216)
);

BUFx2_ASAP7_75t_L g2217 ( 
.A(n_2201),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_2196),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2211),
.B(n_2186),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2205),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2218),
.B(n_2184),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2217),
.B(n_2210),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2206),
.B(n_2184),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2204),
.B(n_2189),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2212),
.Y(n_2225)
);

OAI221xp5_ASAP7_75t_L g2226 ( 
.A1(n_2216),
.A2(n_2190),
.B1(n_2199),
.B2(n_2188),
.C(n_2196),
.Y(n_2226)
);

OR2x2_ASAP7_75t_L g2227 ( 
.A(n_2208),
.B(n_2193),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2207),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2208),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_2213),
.B(n_2203),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2209),
.B(n_2198),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2220),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2222),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2229),
.Y(n_2234)
);

INVx4_ASAP7_75t_L g2235 ( 
.A(n_2231),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2221),
.Y(n_2236)
);

BUFx2_ASAP7_75t_L g2237 ( 
.A(n_2228),
.Y(n_2237)
);

CKINVDCx6p67_ASAP7_75t_R g2238 ( 
.A(n_2223),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2225),
.Y(n_2239)
);

INVx8_ASAP7_75t_L g2240 ( 
.A(n_2230),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2224),
.Y(n_2241)
);

NOR3xp33_ASAP7_75t_L g2242 ( 
.A(n_2235),
.B(n_2226),
.C(n_2219),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2233),
.Y(n_2243)
);

NOR2x1p5_ASAP7_75t_L g2244 ( 
.A(n_2238),
.B(n_2219),
.Y(n_2244)
);

NAND3xp33_ASAP7_75t_L g2245 ( 
.A(n_2235),
.B(n_2227),
.C(n_2215),
.Y(n_2245)
);

NAND3xp33_ASAP7_75t_L g2246 ( 
.A(n_2234),
.B(n_2164),
.C(n_2162),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2237),
.B(n_2157),
.Y(n_2247)
);

OA211x2_ASAP7_75t_L g2248 ( 
.A1(n_2240),
.A2(n_2213),
.B(n_2214),
.C(n_2088),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_2234),
.B(n_2067),
.Y(n_2249)
);

AND4x1_ASAP7_75t_L g2250 ( 
.A(n_2242),
.B(n_2245),
.C(n_2243),
.D(n_2236),
.Y(n_2250)
);

NAND3xp33_ASAP7_75t_SL g2251 ( 
.A(n_2249),
.B(n_2232),
.C(n_2233),
.Y(n_2251)
);

OAI322xp33_ASAP7_75t_SL g2252 ( 
.A1(n_2247),
.A2(n_2241),
.A3(n_2239),
.B1(n_2240),
.B2(n_2164),
.C1(n_2162),
.C2(n_2091),
.Y(n_2252)
);

NOR4xp25_ASAP7_75t_L g2253 ( 
.A(n_2244),
.B(n_2239),
.C(n_2240),
.D(n_2164),
.Y(n_2253)
);

AOI22xp5_ASAP7_75t_L g2254 ( 
.A1(n_2248),
.A2(n_2075),
.B1(n_2148),
.B2(n_2066),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2250),
.B(n_2246),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2251),
.Y(n_2256)
);

OAI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2254),
.A2(n_2162),
.B1(n_2075),
.B2(n_2078),
.Y(n_2257)
);

NOR2x1_ASAP7_75t_L g2258 ( 
.A(n_2253),
.B(n_2078),
.Y(n_2258)
);

NAND3xp33_ASAP7_75t_L g2259 ( 
.A(n_2256),
.B(n_2252),
.C(n_2071),
.Y(n_2259)
);

NAND2xp33_ASAP7_75t_L g2260 ( 
.A(n_2255),
.B(n_2081),
.Y(n_2260)
);

OAI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_2259),
.A2(n_2258),
.B1(n_2257),
.B2(n_2046),
.Y(n_2261)
);

OAI221xp5_ASAP7_75t_R g2262 ( 
.A1(n_2260),
.A2(n_2079),
.B1(n_2069),
.B2(n_2076),
.C(n_2066),
.Y(n_2262)
);

NOR2x1_ASAP7_75t_L g2263 ( 
.A(n_2261),
.B(n_2163),
.Y(n_2263)
);

OR2x2_ASAP7_75t_L g2264 ( 
.A(n_2262),
.B(n_2153),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2264),
.Y(n_2265)
);

AOI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_2265),
.A2(n_2263),
.B1(n_2154),
.B2(n_2160),
.Y(n_2266)
);

INVx1_ASAP7_75t_SL g2267 ( 
.A(n_2266),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2267),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2268),
.Y(n_2269)
);

OAI221xp5_ASAP7_75t_R g2270 ( 
.A1(n_2269),
.A2(n_2133),
.B1(n_2154),
.B2(n_2161),
.C(n_2160),
.Y(n_2270)
);

AOI211xp5_ASAP7_75t_L g2271 ( 
.A1(n_2270),
.A2(n_2154),
.B(n_2160),
.C(n_2166),
.Y(n_2271)
);


endmodule