module fake_jpeg_29223_n_382 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_382);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_46),
.B(n_24),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_21),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_52),
.Y(n_70)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_19),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_22),
.A2(n_10),
.B(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_66),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_24),
.B1(n_41),
.B2(n_37),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_11),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_20),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_76),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_82),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_46),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_103),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_47),
.B(n_26),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_90),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_42),
.B1(n_40),
.B2(n_43),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_100),
.B1(n_25),
.B2(n_41),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_28),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_33),
.B1(n_40),
.B2(n_42),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_64),
.B1(n_33),
.B2(n_66),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_29),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_46),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_120),
.Y(n_141)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_116),
.B1(n_126),
.B2(n_27),
.Y(n_143)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_69),
.B1(n_61),
.B2(n_62),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_111),
.B1(n_133),
.B2(n_64),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_42),
.B1(n_30),
.B2(n_28),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_103),
.B1(n_89),
.B2(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_49),
.B1(n_67),
.B2(n_59),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_31),
.B(n_66),
.Y(n_154)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_132),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_34),
.B(n_27),
.C(n_30),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_137),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_53),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_31),
.Y(n_148)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_71),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_70),
.A2(n_55),
.B1(n_97),
.B2(n_74),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_76),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_138),
.B(n_95),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

BUFx4f_ASAP7_75t_SL g161 ( 
.A(n_139),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_152),
.B1(n_154),
.B2(n_122),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_136),
.B1(n_133),
.B2(n_112),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_33),
.A3(n_66),
.B1(n_79),
.B2(n_28),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_155),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_153),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_98),
.B(n_82),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_150),
.B(n_134),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_87),
.B(n_86),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_107),
.B1(n_123),
.B2(n_108),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_130),
.B(n_60),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_112),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_72),
.B1(n_138),
.B2(n_91),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_156),
.A2(n_91),
.B1(n_95),
.B2(n_48),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_81),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_136),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_123),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_164),
.C(n_128),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_63),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_63),
.Y(n_165)
);

NAND2x1p5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_72),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_118),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_184),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_136),
.B1(n_81),
.B2(n_74),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_192),
.B1(n_196),
.B2(n_198),
.Y(n_207)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

BUFx24_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_178),
.Y(n_210)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_163),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_180),
.A2(n_187),
.B1(n_190),
.B2(n_166),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_189),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_125),
.B(n_137),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_193),
.B(n_150),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_194),
.B(n_145),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_118),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_188),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_73),
.B1(n_124),
.B2(n_127),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_125),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_104),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_73),
.B1(n_129),
.B2(n_113),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_169),
.B(n_147),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_129),
.B1(n_109),
.B2(n_119),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_117),
.B(n_31),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_114),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_131),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_141),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_106),
.B1(n_40),
.B2(n_120),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_170),
.B1(n_161),
.B2(n_168),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_40),
.B1(n_87),
.B2(n_86),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

AOI21x1_ASAP7_75t_L g248 ( 
.A1(n_200),
.A2(n_209),
.B(n_175),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_222),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_142),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_202),
.B(n_206),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_164),
.C(n_153),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_204),
.C(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_182),
.C(n_181),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_165),
.B1(n_154),
.B2(n_157),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_219),
.B1(n_225),
.B2(n_198),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_189),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_211),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_193),
.A2(n_184),
.B(n_173),
.C(n_191),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_212),
.A2(n_218),
.B(n_227),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_148),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_144),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_153),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_151),
.C(n_167),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_194),
.A2(n_154),
.B1(n_166),
.B2(n_168),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_183),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_232),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_172),
.B1(n_196),
.B2(n_195),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_188),
.B1(n_176),
.B2(n_187),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_220),
.B(n_184),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_184),
.B1(n_190),
.B2(n_154),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_207),
.A2(n_162),
.B1(n_159),
.B2(n_146),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_253),
.B1(n_32),
.B2(n_35),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_199),
.B1(n_162),
.B2(n_159),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_235),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_220),
.B(n_214),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_241),
.C(n_203),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_199),
.B1(n_146),
.B2(n_29),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_225),
.B1(n_224),
.B2(n_206),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_151),
.B1(n_170),
.B2(n_167),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_170),
.B1(n_175),
.B2(n_177),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_246),
.B1(n_212),
.B2(n_216),
.Y(n_270)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_175),
.B1(n_177),
.B2(n_27),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_95),
.B(n_50),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_161),
.Y(n_250)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_252),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_212),
.A2(n_175),
.B1(n_30),
.B2(n_35),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_250),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_271),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_260),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_282),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_210),
.C(n_200),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_266),
.C(n_238),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_212),
.C(n_221),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_212),
.B1(n_221),
.B2(n_216),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_270),
.B1(n_278),
.B2(n_281),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_16),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_279),
.B1(n_246),
.B2(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_32),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_273),
.Y(n_294)
);

AOI21x1_ASAP7_75t_L g300 ( 
.A1(n_274),
.A2(n_277),
.B(n_280),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_244),
.Y(n_276)
);

NOR3xp33_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_139),
.C(n_9),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_0),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_230),
.A2(n_25),
.B1(n_37),
.B2(n_9),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_237),
.A2(n_14),
.B1(n_19),
.B2(n_17),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_242),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_139),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_2),
.B(n_3),
.Y(n_302)
);

A2O1A1O1Ixp25_ASAP7_75t_L g282 ( 
.A1(n_232),
.A2(n_95),
.B(n_63),
.C(n_139),
.D(n_33),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_256),
.B(n_248),
.C(n_243),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_283),
.A2(n_264),
.B(n_262),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_287),
.C(n_8),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_241),
.C(n_229),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_291),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_289),
.B(n_279),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_290),
.A2(n_302),
.B1(n_276),
.B2(n_277),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_265),
.B(n_236),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_256),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_298),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_259),
.B(n_236),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_295),
.B(n_303),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_260),
.A2(n_247),
.B1(n_245),
.B2(n_251),
.Y(n_296)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_297)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_297),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_263),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_301),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_281),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_8),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_293),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_280),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_313),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_308),
.B(n_315),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_268),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_302),
.Y(n_334)
);

XNOR2x1_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_282),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_283),
.A2(n_275),
.B1(n_258),
.B2(n_262),
.Y(n_314)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_275),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_318),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_258),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_285),
.B(n_264),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_319),
.B(n_322),
.Y(n_333)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_305),
.A2(n_283),
.B1(n_300),
.B2(n_294),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_324),
.A2(n_313),
.B1(n_310),
.B2(n_13),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_306),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_331),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_284),
.C(n_303),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_335),
.C(n_7),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_304),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_284),
.Y(n_332)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_332),
.Y(n_339)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_283),
.C(n_12),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_312),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_336),
.B(n_337),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_322),
.B(n_12),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_309),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_320),
.B(n_314),
.Y(n_340)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_349),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_326),
.A2(n_317),
.B(n_307),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_342),
.A2(n_346),
.B(n_343),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_343),
.B(n_329),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_345),
.B(n_348),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_335),
.A2(n_17),
.B(n_13),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_334),
.B(n_15),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_351),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_2),
.Y(n_351)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_358),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_345),
.A2(n_324),
.B(n_325),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_356),
.A2(n_3),
.B(n_5),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_329),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_357),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_323),
.C(n_330),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_361),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_327),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_325),
.C(n_4),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_362),
.B(n_353),
.Y(n_365)
);

NAND2x1_ASAP7_75t_SL g363 ( 
.A(n_360),
.B(n_347),
.Y(n_363)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_363),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_359),
.A2(n_344),
.B1(n_4),
.B2(n_5),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_364),
.B(n_365),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_366),
.A2(n_362),
.B(n_352),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_371),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_368),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_374),
.Y(n_378)
);

O2A1O1Ixp33_ASAP7_75t_SL g375 ( 
.A1(n_369),
.A2(n_357),
.B(n_361),
.C(n_3),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_375),
.A2(n_376),
.B(n_365),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_370),
.A2(n_3),
.B(n_5),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_377),
.A2(n_372),
.B(n_373),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_378),
.C(n_379),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_381),
.B(n_367),
.Y(n_382)
);


endmodule