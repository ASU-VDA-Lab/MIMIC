module fake_jpeg_6174_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_10),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.C(n_1),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_24),
.B1(n_30),
.B2(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_21),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_23),
.B(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_31),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_47),
.Y(n_85)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_61),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_17),
.B1(n_23),
.B2(n_30),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_63),
.B1(n_71),
.B2(n_22),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_17),
.B1(n_32),
.B2(n_25),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_57),
.B1(n_62),
.B2(n_67),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_17),
.B1(n_32),
.B2(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_25),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_26),
.B1(n_27),
.B2(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_19),
.B1(n_18),
.B2(n_22),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_41),
.B1(n_40),
.B2(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_24),
.B1(n_22),
.B2(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_38),
.B(n_44),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_87),
.C(n_91),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_84),
.B1(n_93),
.B2(n_67),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_57),
.B(n_19),
.C(n_27),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_53),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_39),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_46),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_41),
.B1(n_40),
.B2(n_35),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_38),
.C(n_44),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_96),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_29),
.B(n_28),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_41),
.B1(n_33),
.B2(n_32),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_58),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_98),
.A2(n_104),
.B1(n_109),
.B2(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_65),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_99),
.Y(n_144)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_103),
.Y(n_132)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_62),
.B1(n_56),
.B2(n_52),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_50),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_72),
.B1(n_59),
.B2(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_94),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_77),
.A2(n_59),
.B1(n_48),
.B2(n_68),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_87),
.B1(n_95),
.B2(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_49),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_122),
.Y(n_140)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

OAI32xp33_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_69),
.A3(n_66),
.B1(n_36),
.B2(n_59),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_86),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_60),
.Y(n_122)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_68),
.B(n_36),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_123),
.A2(n_68),
.B1(n_93),
.B2(n_120),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_75),
.B1(n_79),
.B2(n_81),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_105),
.B1(n_112),
.B2(n_115),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_88),
.B1(n_91),
.B2(n_87),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_139),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_123),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_146),
.B1(n_147),
.B2(n_39),
.Y(n_170)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_97),
.C(n_92),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_73),
.C(n_80),
.Y(n_175)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_151),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_98),
.A2(n_97),
.B1(n_92),
.B2(n_74),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_109),
.B1(n_121),
.B2(n_102),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_102),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_94),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_152),
.A2(n_113),
.B(n_123),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_153),
.A2(n_170),
.B1(n_39),
.B2(n_129),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_123),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_111),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_166),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_171),
.B(n_178),
.Y(n_200)
);

AO22x1_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_107),
.B1(n_113),
.B2(n_94),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_159),
.A2(n_144),
.B1(n_134),
.B2(n_152),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_118),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_74),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_73),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_144),
.B(n_16),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_174),
.Y(n_193)
);

CKINVDCx10_ASAP7_75t_R g164 ( 
.A(n_145),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_168),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_49),
.B(n_103),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_16),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_143),
.C(n_147),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_80),
.B(n_2),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_151),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_132),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_188),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_191),
.C(n_194),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_165),
.B(n_126),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_190),
.B(n_195),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_136),
.C(n_134),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_197),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_170),
.C(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_159),
.A2(n_136),
.B1(n_129),
.B2(n_127),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_178),
.B(n_172),
.Y(n_218)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_169),
.A2(n_45),
.B1(n_100),
.B2(n_119),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_36),
.C(n_45),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_171),
.C(n_180),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_29),
.Y(n_207)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_194),
.A2(n_198),
.B1(n_189),
.B2(n_153),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_211),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_177),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_213),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_189),
.B(n_158),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_166),
.B(n_2),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_220),
.C(n_223),
.Y(n_235)
);

NOR3xp33_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_159),
.C(n_173),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_219),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_168),
.Y(n_241)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_191),
.C(n_206),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_172),
.C(n_155),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_177),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_203),
.C(n_196),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_197),
.C(n_187),
.Y(n_236)
);

AOI22x1_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_45),
.B1(n_36),
.B2(n_174),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_228),
.A2(n_201),
.B1(n_181),
.B2(n_182),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_161),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_230),
.Y(n_243)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_186),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_33),
.B(n_2),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_179),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_207),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_236),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_237),
.A2(n_248),
.B1(n_228),
.B2(n_232),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_193),
.C(n_163),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_240),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_193),
.C(n_186),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_246),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_251),
.B(n_229),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_224),
.B(n_8),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_31),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_33),
.C(n_31),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_247),
.B(n_252),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_227),
.A2(n_33),
.B1(n_7),
.B2(n_8),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_225),
.B(n_222),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_250),
.A2(n_224),
.B(n_215),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_0),
.C(n_2),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_7),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_252),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_211),
.Y(n_254)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_256),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_257),
.A2(n_265),
.B(n_266),
.Y(n_282)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

AO221x1_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_241),
.B1(n_253),
.B2(n_234),
.C(n_235),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_255),
.A2(n_216),
.B1(n_208),
.B2(n_249),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_262),
.B(n_263),
.Y(n_278)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_265),
.B(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_208),
.B(n_230),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_254),
.A2(n_216),
.B1(n_226),
.B2(n_212),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_269),
.B1(n_239),
.B2(n_240),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_268),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_228),
.B1(n_231),
.B2(n_210),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_274),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_283),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_235),
.C(n_247),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_285),
.C(n_289),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

XOR2x2_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_8),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_9),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_258),
.B1(n_273),
.B2(n_274),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_0),
.C(n_3),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_257),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_262),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_4),
.C(n_5),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_4),
.C(n_5),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_6),
.C(n_9),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_6),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_259),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_297),
.B(n_300),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_261),
.B(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_259),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_275),
.C(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_286),
.C(n_280),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_6),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_303),
.A2(n_290),
.B(n_283),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_304),
.A2(n_282),
.B(n_288),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_293),
.Y(n_318)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_280),
.B1(n_281),
.B2(n_289),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_308),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_311),
.B(n_314),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_6),
.Y(n_311)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_292),
.B(n_291),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_317),
.B(n_318),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_304),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_302),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_322),
.C(n_311),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_295),
.Y(n_322)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_324),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_312),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_326),
.B(n_327),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_307),
.B(n_14),
.C(n_15),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_12),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_12),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_323),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_330),
.B(n_328),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_15),
.Y(n_333)
);


endmodule