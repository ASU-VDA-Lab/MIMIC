module fake_jpeg_3841_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

OR2x2_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_40),
.B(n_25),
.C(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_18),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_38),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_27),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_14),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_15),
.B1(n_19),
.B2(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_25),
.B1(n_17),
.B2(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_52),
.B1(n_54),
.B2(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_42),
.CI(n_32),
.CON(n_76),
.SN(n_76)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_25),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_15),
.B1(n_17),
.B2(n_19),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_23),
.B1(n_29),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_60),
.B1(n_43),
.B2(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_58),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_20),
.B1(n_29),
.B2(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_16),
.B1(n_27),
.B2(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_32),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_53),
.Y(n_88)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_SL g85 ( 
.A(n_68),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_83),
.B1(n_50),
.B2(n_43),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_77),
.Y(n_103)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_80),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_46),
.B1(n_63),
.B2(n_44),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_49),
.B1(n_44),
.B2(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_39),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_39),
.B1(n_35),
.B2(n_38),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_88),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_78),
.B1(n_66),
.B2(n_73),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_94),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_59),
.B1(n_50),
.B2(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

OR2x2_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_13),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_101),
.B(n_102),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_16),
.B(n_24),
.C(n_31),
.Y(n_128)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_49),
.B(n_64),
.C(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_58),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_69),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_38),
.B1(n_31),
.B2(n_21),
.Y(n_100)
);

XNOR2x1_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_44),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_47),
.C(n_28),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_28),
.B(n_22),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_74),
.B(n_67),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_111),
.B(n_112),
.Y(n_142)
);

AO21x1_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_76),
.B(n_67),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_99),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_119),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_84),
.B(n_22),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_126),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_87),
.B(n_94),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_128),
.B(n_72),
.Y(n_143)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

AO21x2_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_84),
.B(n_24),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_90),
.B1(n_72),
.B2(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_106),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_92),
.B(n_86),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_137),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_89),
.C(n_102),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_138),
.C(n_117),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_93),
.B1(n_104),
.B2(n_88),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_146),
.B1(n_128),
.B2(n_125),
.Y(n_152)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_122),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_95),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_96),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_143),
.B(n_147),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_150),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_106),
.B1(n_24),
.B2(n_31),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_106),
.B(n_28),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_28),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_22),
.B(n_28),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_128),
.B1(n_125),
.B2(n_113),
.Y(n_167)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_28),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_109),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_160),
.B1(n_165),
.B2(n_167),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_150),
.B(n_116),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_166),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_107),
.C(n_111),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_109),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_121),
.B1(n_108),
.B2(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_22),
.B(n_24),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_117),
.C(n_119),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_163),
.B(n_148),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_172),
.C(n_138),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_128),
.B1(n_125),
.B2(n_119),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_115),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_133),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_125),
.C(n_128),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_142),
.B1(n_140),
.B2(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_180),
.C(n_181),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_145),
.B1(n_139),
.B2(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_144),
.C(n_147),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_146),
.C(n_136),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_184),
.C(n_177),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_47),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_170),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_134),
.C(n_133),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_162),
.A2(n_21),
.B1(n_16),
.B2(n_2),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_21),
.B1(n_1),
.B2(n_0),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_165),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_204),
.B1(n_191),
.B2(n_190),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_169),
.C(n_170),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_5),
.Y(n_216)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_197),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_181),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_187),
.A2(n_171),
.B1(n_168),
.B2(n_153),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_200),
.B(n_188),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_161),
.C(n_156),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_184),
.C(n_173),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_159),
.B1(n_21),
.B2(n_5),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_206),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_212),
.C(n_216),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_217),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_218),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_193),
.A2(n_175),
.B1(n_185),
.B2(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_189),
.B1(n_175),
.B2(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_6),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_6),
.C(n_7),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_6),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_219),
.B(n_206),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_205),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_223),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_203),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_211),
.B(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_213),
.B1(n_218),
.B2(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_225),
.Y(n_233)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_235),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_237),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_9),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_197),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_236),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_225),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_222),
.A2(n_196),
.B(n_8),
.Y(n_236)
);

OAI321xp33_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_196),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_7),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_230),
.A2(n_229),
.B1(n_224),
.B2(n_227),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_243),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_231),
.B(n_8),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_11),
.C(n_13),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_232),
.B(n_12),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_246),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_11),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_13),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

AOI221xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_240),
.B1(n_247),
.B2(n_249),
.C(n_235),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_240),
.Y(n_252)
);


endmodule