module fake_jpeg_30266_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_0),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_51),
.Y(n_78)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_70),
.Y(n_81)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_70),
.A2(n_61),
.B1(n_44),
.B2(n_46),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_83),
.B1(n_6),
.B2(n_7),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_49),
.B(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_2),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_3),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_59),
.B1(n_57),
.B2(n_56),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_55),
.B1(n_50),
.B2(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_5),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_86),
.B(n_25),
.Y(n_118)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_87),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_92),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_52),
.B1(n_47),
.B2(n_23),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_102),
.B1(n_77),
.B2(n_10),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_95),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_94),
.Y(n_115)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_14),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_5),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_22),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_100),
.A2(n_8),
.B(n_9),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_7),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_101),
.B(n_9),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_26),
.B1(n_42),
.B2(n_41),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_111),
.B(n_113),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_107),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_11),
.B(n_12),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_17),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_21),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_24),
.Y(n_117)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_27),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_43),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_108),
.C(n_103),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_100),
.B1(n_31),
.B2(n_34),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

NOR4xp25_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_104),
.C(n_126),
.D(n_123),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_29),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_132),
.B(n_107),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_135),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_112),
.C(n_115),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_122),
.C(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_137),
.B(n_127),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_138),
.B1(n_131),
.B2(n_130),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_133),
.B(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_114),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);


endmodule