module fake_jpeg_17440_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_1),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_13),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_26),
.Y(n_30)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_24),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_13),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_16),
.B1(n_10),
.B2(n_27),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_27),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_14),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_16),
.B1(n_19),
.B2(n_10),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_24),
.B1(n_21),
.B2(n_3),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_22),
.A2(n_19),
.B1(n_12),
.B2(n_18),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_46),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_35),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_41),
.B(n_29),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_4),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_5),
.C(n_6),
.Y(n_58)
);

OAI22x1_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_41),
.B1(n_48),
.B2(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_48),
.B1(n_29),
.B2(n_43),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_32),
.C(n_33),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_3),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_55),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_2),
.B1(n_3),
.B2(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_55),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_63),
.B(n_59),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_61),
.C(n_63),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_71),
.C(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_65),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.C(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_53),
.Y(n_76)
);


endmodule