module real_aes_7522_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_1106;
wire n_800;
wire n_778;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_792;
wire n_673;
wire n_386;
wire n_635;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_1064;
wire n_540;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_852;
wire n_766;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_955;
wire n_696;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_951;
wire n_467;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_931;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_960;
wire n_725;
wire n_1081;
wire n_671;
wire n_973;
wire n_1084;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1017;
wire n_737;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1103;
wire n_1037;
wire n_1031;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_898;
wire n_734;
wire n_604;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_727;
wire n_1014;
wire n_397;
wire n_649;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_1002;
wire n_934;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_972;
wire n_1127;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_717;
wire n_456;
wire n_982;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_1114;
wire n_871;
wire n_1045;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_1055;
wire n_988;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_646;
wire n_650;
wire n_743;
wire n_710;
wire n_393;
wire n_652;
wire n_703;
wire n_823;
wire n_500;
wire n_601;
wire n_1097;
wire n_1076;
wire n_463;
wire n_661;
wire n_804;
wire n_396;
wire n_1101;
wire n_447;
wire n_1102;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1039;
wire n_802;
wire n_868;
wire n_877;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_1104;
wire n_842;
wire n_1061;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_0), .A2(n_173), .B1(n_626), .B2(n_627), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_1), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_2), .B(n_489), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_3), .B(n_484), .Y(n_858) );
OA22x2_ASAP7_75t_L g396 ( .A1(n_4), .A2(n_397), .B1(n_398), .B2(n_490), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_4), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_5), .A2(n_162), .B1(n_619), .B2(n_649), .C(n_820), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_6), .A2(n_293), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_7), .A2(n_940), .B1(n_967), .B2(n_968), .Y(n_939) );
INVx1_ASAP7_75t_L g968 ( .A(n_7), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_8), .A2(n_349), .B1(n_839), .B2(n_840), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_9), .Y(n_512) );
AO22x2_ASAP7_75t_L g415 ( .A1(n_10), .A2(n_227), .B1(n_407), .B2(n_412), .Y(n_415) );
INVx1_ASAP7_75t_L g1072 ( .A(n_10), .Y(n_1072) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_11), .A2(n_212), .B1(n_716), .B2(n_717), .Y(n_715) );
AOI22xp5_ASAP7_75t_SL g1003 ( .A1(n_12), .A2(n_380), .B1(n_530), .B2(n_627), .Y(n_1003) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_13), .A2(n_305), .B1(n_480), .B2(n_508), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_14), .A2(n_63), .B1(n_745), .B2(n_746), .Y(n_744) );
AOI22xp5_ASAP7_75t_SL g999 ( .A1(n_15), .A2(n_254), .B1(n_523), .B2(n_868), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_16), .A2(n_105), .B1(n_521), .B2(n_711), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_17), .A2(n_23), .B1(n_550), .B2(n_589), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_18), .Y(n_963) );
CKINVDCx20_ASAP7_75t_R g1118 ( .A(n_19), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_20), .A2(n_381), .B1(n_531), .B2(n_644), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_21), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_22), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_24), .A2(n_273), .B1(n_441), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_25), .A2(n_338), .B1(n_651), .B2(n_751), .Y(n_859) );
AOI22xp33_ASAP7_75t_SL g997 ( .A1(n_26), .A2(n_174), .B1(n_591), .B2(n_652), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_27), .A2(n_341), .B1(n_445), .B2(n_543), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_28), .A2(n_107), .B1(n_629), .B2(n_789), .Y(n_951) );
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_29), .A2(n_51), .B1(n_642), .B2(n_758), .Y(n_757) );
AO22x2_ASAP7_75t_L g417 ( .A1(n_30), .A2(n_111), .B1(n_407), .B2(n_408), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_31), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_32), .A2(n_268), .B1(n_567), .B2(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_33), .A2(n_52), .B1(n_656), .B2(n_840), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_34), .A2(n_204), .B1(n_440), .B2(n_443), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g1081 ( .A1(n_35), .A2(n_99), .B1(n_745), .B2(n_1020), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_36), .A2(n_284), .B1(n_655), .B2(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_37), .Y(n_1028) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_38), .A2(n_326), .B1(n_629), .B2(n_631), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_39), .A2(n_231), .B1(n_656), .B2(n_975), .Y(n_974) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_40), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_41), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g541 ( .A1(n_42), .A2(n_280), .B1(n_436), .B2(n_451), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_43), .B(n_617), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_44), .B(n_614), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_45), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_46), .Y(n_924) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_47), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_48), .A2(n_198), .B1(n_612), .B2(n_614), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_49), .A2(n_146), .B1(n_523), .B2(n_526), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_50), .A2(n_360), .B1(n_566), .B2(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_53), .B(n_510), .Y(n_509) );
AOI222xp33_ASAP7_75t_L g824 ( .A1(n_54), .A2(n_221), .B1(n_318), .B2(n_612), .C1(n_825), .C2(n_826), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g866 ( .A1(n_55), .A2(n_322), .B1(n_530), .B2(n_711), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g882 ( .A(n_56), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_57), .A2(n_223), .B1(n_531), .B2(n_918), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_58), .A2(n_190), .B1(n_440), .B2(n_915), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_59), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g1021 ( .A(n_60), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g1043 ( .A(n_61), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_62), .B(n_583), .Y(n_1115) );
CKINVDCx20_ASAP7_75t_R g927 ( .A(n_64), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_65), .A2(n_364), .B1(n_426), .B2(n_441), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_66), .A2(n_302), .B1(n_559), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_67), .A2(n_213), .B1(n_784), .B2(n_792), .Y(n_902) );
INVx1_ASAP7_75t_L g1005 ( .A(n_68), .Y(n_1005) );
AOI222xp33_ASAP7_75t_L g985 ( .A1(n_69), .A2(n_210), .B1(n_245), .B2(n_460), .C1(n_659), .C2(n_986), .Y(n_985) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_70), .Y(n_1023) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_71), .Y(n_965) );
AOI22xp33_ASAP7_75t_SL g1046 ( .A1(n_72), .A2(n_214), .B1(n_481), .B2(n_589), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_73), .A2(n_134), .B1(n_644), .B2(n_1125), .Y(n_1124) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_74), .A2(n_277), .B1(n_434), .B2(n_533), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_75), .A2(n_286), .B1(n_758), .B2(n_784), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_76), .A2(n_98), .B1(n_424), .B2(n_434), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_77), .A2(n_262), .B1(n_466), .B2(n_478), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_78), .A2(n_155), .B1(n_627), .B2(n_868), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g944 ( .A(n_79), .Y(n_944) );
AOI22xp5_ASAP7_75t_SL g1000 ( .A1(n_80), .A2(n_259), .B1(n_526), .B2(n_1001), .Y(n_1000) );
AOI22xp33_ASAP7_75t_SL g750 ( .A1(n_81), .A2(n_232), .B1(n_673), .B2(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_82), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_83), .A2(n_94), .B1(n_634), .B2(n_794), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_84), .A2(n_308), .B1(n_531), .B2(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_85), .A2(n_116), .B1(n_523), .B2(n_758), .Y(n_983) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_86), .Y(n_546) );
AO22x2_ASAP7_75t_L g411 ( .A1(n_87), .A2(n_267), .B1(n_407), .B2(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g1069 ( .A(n_87), .Y(n_1069) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_88), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_89), .A2(n_264), .B1(n_449), .B2(n_527), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_90), .A2(n_369), .B1(n_789), .B2(n_1128), .Y(n_1127) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_91), .Y(n_768) );
AOI22xp33_ASAP7_75t_SL g1087 ( .A1(n_92), .A2(n_319), .B1(n_418), .B2(n_1088), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_93), .A2(n_379), .B1(n_535), .B2(n_642), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_95), .Y(n_946) );
AOI22xp5_ASAP7_75t_SL g1004 ( .A1(n_96), .A2(n_217), .B1(n_434), .B2(n_784), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_97), .A2(n_303), .B1(n_642), .B2(n_645), .Y(n_984) );
AOI211xp5_ASAP7_75t_L g1089 ( .A1(n_100), .A2(n_868), .B(n_1090), .C(n_1093), .Y(n_1089) );
AOI22xp33_ASAP7_75t_SL g1083 ( .A1(n_101), .A2(n_290), .B1(n_477), .B2(n_480), .Y(n_1083) );
AOI222xp33_ASAP7_75t_L g658 ( .A1(n_102), .A2(n_237), .B1(n_248), .B2(n_460), .C1(n_480), .C2(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g592 ( .A(n_103), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_104), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_106), .A2(n_199), .B1(n_508), .B2(n_550), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_108), .A2(n_205), .B1(n_484), .B2(n_487), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g909 ( .A1(n_109), .A2(n_910), .B1(n_933), .B2(n_934), .Y(n_909) );
INVx1_ASAP7_75t_L g933 ( .A(n_109), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_110), .A2(n_178), .B1(n_465), .B2(n_478), .Y(n_731) );
INVx1_ASAP7_75t_L g1073 ( .A(n_111), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_112), .A2(n_258), .B1(n_644), .B2(n_645), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_113), .B(n_929), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g1017 ( .A(n_114), .Y(n_1017) );
XOR2xp5_ASAP7_75t_L g639 ( .A(n_115), .B(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g981 ( .A1(n_117), .A2(n_335), .B1(n_478), .B2(n_550), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g633 ( .A1(n_118), .A2(n_202), .B1(n_402), .B2(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_119), .B(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_120), .A2(n_332), .B1(n_567), .B2(n_677), .Y(n_1050) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_121), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_122), .A2(n_191), .B1(n_898), .B2(n_915), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_123), .A2(n_315), .B1(n_648), .B2(n_649), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_124), .A2(n_216), .B1(n_621), .B2(n_622), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_125), .A2(n_359), .B1(n_792), .B2(n_898), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_126), .A2(n_247), .B1(n_784), .B2(n_785), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_127), .A2(n_142), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g1075 ( .A1(n_128), .A2(n_1076), .B1(n_1077), .B2(n_1095), .Y(n_1075) );
CKINVDCx20_ASAP7_75t_R g1095 ( .A(n_128), .Y(n_1095) );
AOI22xp33_ASAP7_75t_SL g754 ( .A1(n_129), .A2(n_187), .B1(n_567), .B2(n_655), .Y(n_754) );
AOI22xp33_ASAP7_75t_SL g872 ( .A1(n_130), .A2(n_328), .B1(n_526), .B2(n_566), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_131), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_132), .A2(n_336), .B1(n_642), .B2(n_789), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_133), .A2(n_249), .B1(n_478), .B2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_135), .A2(n_255), .B1(n_477), .B2(n_480), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_136), .A2(n_366), .B1(n_794), .B2(n_797), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_137), .A2(n_346), .B1(n_508), .B2(n_612), .Y(n_993) );
AOI22xp33_ASAP7_75t_SL g448 ( .A1(n_138), .A2(n_211), .B1(n_449), .B2(n_454), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_139), .A2(n_194), .B1(n_487), .B2(n_553), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_140), .A2(n_361), .B1(n_792), .B2(n_840), .Y(n_1036) );
XNOR2x2_ASAP7_75t_L g832 ( .A(n_141), .B(n_833), .Y(n_832) );
OA22x2_ASAP7_75t_L g851 ( .A1(n_143), .A2(n_852), .B1(n_853), .B2(n_873), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_143), .Y(n_852) );
INVx1_ASAP7_75t_L g683 ( .A(n_144), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_145), .B(n_489), .Y(n_554) );
AND2x6_ASAP7_75t_L g385 ( .A(n_147), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1066 ( .A(n_147), .Y(n_1066) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_148), .A2(n_368), .B1(n_530), .B2(n_531), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_149), .A2(n_189), .B1(n_402), .B2(n_681), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_150), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_151), .B(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_152), .A2(n_350), .B1(n_533), .B2(n_535), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_153), .B(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g1044 ( .A1(n_154), .A2(n_276), .B1(n_704), .B2(n_826), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_156), .Y(n_978) );
AO22x1_ASAP7_75t_L g800 ( .A1(n_157), .A2(n_801), .B1(n_827), .B2(n_828), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_157), .Y(n_827) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_158), .A2(n_179), .B1(n_681), .B2(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_159), .B(n_670), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_160), .Y(n_705) );
AOI222xp33_ASAP7_75t_L g846 ( .A1(n_161), .A2(n_215), .B1(n_342), .B2(n_510), .C1(n_583), .C2(n_704), .Y(n_846) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_163), .A2(n_240), .B1(n_553), .B2(n_617), .Y(n_1084) );
CKINVDCx20_ASAP7_75t_R g1117 ( .A(n_164), .Y(n_1117) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_165), .A2(n_256), .B1(n_407), .B2(n_408), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g1070 ( .A(n_165), .B(n_1071), .Y(n_1070) );
CKINVDCx20_ASAP7_75t_R g1011 ( .A(n_166), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_167), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g1094 ( .A(n_168), .Y(n_1094) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_169), .A2(n_295), .B1(n_403), .B2(n_428), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_170), .Y(n_956) );
AOI22xp33_ASAP7_75t_SL g1031 ( .A1(n_171), .A2(n_182), .B1(n_796), .B2(n_839), .Y(n_1031) );
AOI22xp33_ASAP7_75t_SL g1086 ( .A1(n_172), .A2(n_275), .B1(n_535), .B2(n_797), .Y(n_1086) );
CKINVDCx20_ASAP7_75t_R g926 ( .A(n_175), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_176), .A2(n_209), .B1(n_533), .B2(n_681), .Y(n_1051) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_177), .A2(n_183), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_180), .A2(n_269), .B1(n_441), .B2(n_642), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_181), .A2(n_192), .B1(n_484), .B2(n_487), .Y(n_1047) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_184), .A2(n_325), .B1(n_449), .B2(n_631), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_185), .A2(n_317), .B1(n_440), .B2(n_792), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g802 ( .A1(n_186), .A2(n_208), .B1(n_443), .B2(n_803), .C(n_804), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_188), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g1109 ( .A(n_193), .Y(n_1109) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_195), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_196), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_197), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g1080 ( .A(n_200), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_201), .A2(n_307), .B1(n_566), .B2(n_645), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_203), .B(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_206), .A2(n_257), .B1(n_426), .B2(n_441), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_207), .A2(n_304), .B1(n_788), .B2(n_789), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g1112 ( .A(n_218), .Y(n_1112) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_219), .A2(n_383), .B(n_391), .C(n_1074), .Y(n_382) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_220), .A2(n_246), .B1(n_521), .B2(n_523), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_222), .A2(n_239), .B1(n_525), .B2(n_526), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g810 ( .A1(n_224), .A2(n_243), .B1(n_531), .B2(n_811), .C(n_812), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_225), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_226), .A2(n_344), .B1(n_788), .B2(n_818), .Y(n_920) );
NAND2xp5_ASAP7_75t_SL g996 ( .A(n_228), .B(n_619), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_229), .A2(n_327), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_230), .A2(n_272), .B1(n_445), .B2(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_233), .A2(n_310), .B1(n_789), .B2(n_900), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_234), .B(n_631), .Y(n_1092) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_235), .Y(n_888) );
OA22x2_ASAP7_75t_L g492 ( .A1(n_236), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_236), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_238), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_241), .A2(n_260), .B1(n_677), .B2(n_713), .Y(n_976) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_242), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_244), .A2(n_329), .B1(n_443), .B2(n_656), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g1027 ( .A(n_250), .Y(n_1027) );
CKINVDCx20_ASAP7_75t_R g992 ( .A(n_251), .Y(n_992) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_252), .A2(n_301), .B1(n_543), .B2(n_677), .Y(n_722) );
AND2x2_ASAP7_75t_L g389 ( .A(n_253), .B(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_261), .A2(n_289), .B1(n_589), .B2(n_591), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_263), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_265), .Y(n_773) );
XNOR2x1_ASAP7_75t_L g739 ( .A(n_266), .B(n_740), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_270), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_271), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_274), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g1114 ( .A(n_278), .Y(n_1114) );
OA22x2_ASAP7_75t_L g1037 ( .A1(n_279), .A2(n_1038), .B1(n_1039), .B2(n_1055), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g1038 ( .A(n_279), .Y(n_1038) );
AOI22xp33_ASAP7_75t_SL g1034 ( .A1(n_281), .A2(n_300), .B1(n_426), .B2(n_1035), .Y(n_1034) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_282), .Y(n_954) );
AOI22x1_ASAP7_75t_L g764 ( .A1(n_283), .A2(n_765), .B1(n_798), .B2(n_799), .Y(n_764) );
INVx1_ASAP7_75t_L g798 ( .A(n_283), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_285), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_287), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_288), .B(n_619), .Y(n_980) );
INVx1_ASAP7_75t_L g407 ( .A(n_291), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_291), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_292), .Y(n_1025) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_294), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g1110 ( .A(n_296), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_297), .B(n_484), .Y(n_587) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_298), .A2(n_330), .B1(n_525), .B2(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_299), .A2(n_367), .B1(n_402), .B2(n_418), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_306), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_309), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_311), .A2(n_605), .B1(n_606), .B2(n_636), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_311), .Y(n_605) );
XNOR2x1_ASAP7_75t_L g689 ( .A(n_312), .B(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_313), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_314), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_316), .Y(n_736) );
INVx1_ASAP7_75t_L g390 ( .A(n_320), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_321), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_323), .Y(n_886) );
INVx1_ASAP7_75t_L g386 ( .A(n_324), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_331), .A2(n_375), .B1(n_472), .B2(n_480), .Y(n_700) );
XOR2x2_ASAP7_75t_L g875 ( .A(n_333), .B(n_876), .Y(n_875) );
AOI22xp33_ASAP7_75t_SL g870 ( .A1(n_334), .A2(n_340), .B1(n_434), .B2(n_871), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_337), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_339), .B(n_648), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_343), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_345), .A2(n_374), .B1(n_549), .B2(n_550), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_347), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_348), .B(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g582 ( .A1(n_351), .A2(n_356), .B1(n_507), .B2(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_352), .A2(n_362), .B1(n_434), .B2(n_711), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g961 ( .A(n_353), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g1091 ( .A(n_354), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_355), .A2(n_377), .B1(n_631), .B2(n_642), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_357), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_358), .B(n_489), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g949 ( .A(n_363), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_365), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_370), .B(n_507), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_371), .Y(n_610) );
INVx1_ASAP7_75t_L g1104 ( .A(n_372), .Y(n_1104) );
OA22x2_ASAP7_75t_L g1105 ( .A1(n_372), .A2(n_1104), .B1(n_1106), .B2(n_1129), .Y(n_1105) );
CKINVDCx20_ASAP7_75t_R g1016 ( .A(n_373), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g987 ( .A(n_376), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_378), .B(n_857), .Y(n_995) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
HB1xp67_ASAP7_75t_L g1065 ( .A(n_386), .Y(n_1065) );
OAI21xp5_ASAP7_75t_L g1102 ( .A1(n_387), .A2(n_1064), .B(n_1103), .Y(n_1102) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_907), .B1(n_908), .B2(n_1060), .C(n_1061), .Y(n_391) );
INVxp67_ASAP7_75t_L g1060 ( .A(n_392), .Y(n_1060) );
XOR2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_762), .Y(n_392) );
XNOR2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_597), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_491), .B2(n_596), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g490 ( .A(n_398), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_457), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_438), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_423), .Y(n_400) );
BUFx4f_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g841 ( .A(n_403), .Y(n_841) );
BUFx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g530 ( .A(n_404), .Y(n_530) );
BUFx3_ASAP7_75t_L g655 ( .A(n_404), .Y(n_655) );
BUFx3_ASAP7_75t_L g677 ( .A(n_404), .Y(n_677) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_413), .Y(n_404) );
AND2x2_ASAP7_75t_L g453 ( .A(n_405), .B(n_437), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_405), .B(n_413), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g815 ( .A(n_405), .B(n_437), .Y(n_815) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_410), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_406), .B(n_411), .Y(n_422) );
INVx2_ASAP7_75t_L g432 ( .A(n_406), .Y(n_432) );
AND2x2_ASAP7_75t_L g469 ( .A(n_406), .B(n_415), .Y(n_469) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_409), .Y(n_412) );
INVx1_ASAP7_75t_L g482 ( .A(n_410), .Y(n_482) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g433 ( .A(n_411), .Y(n_433) );
AND2x2_ASAP7_75t_L g447 ( .A(n_411), .B(n_432), .Y(n_447) );
INVx1_ASAP7_75t_L g468 ( .A(n_411), .Y(n_468) );
AND2x4_ASAP7_75t_L g420 ( .A(n_413), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g442 ( .A(n_413), .B(n_431), .Y(n_442) );
AND2x4_ASAP7_75t_L g446 ( .A(n_413), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
OR2x2_ASAP7_75t_L g430 ( .A(n_414), .B(n_417), .Y(n_430) );
AND2x2_ASAP7_75t_L g437 ( .A(n_414), .B(n_417), .Y(n_437) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g462 ( .A(n_415), .B(n_417), .Y(n_462) );
AND2x2_ASAP7_75t_L g467 ( .A(n_416), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g514 ( .A(n_416), .Y(n_514) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g456 ( .A(n_417), .Y(n_456) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI221xp5_ASAP7_75t_SL g948 ( .A1(n_419), .A2(n_919), .B1(n_949), .B2(n_950), .C(n_951), .Y(n_948) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g531 ( .A(n_420), .Y(n_531) );
BUFx3_ASAP7_75t_L g559 ( .A(n_420), .Y(n_559) );
BUFx2_ASAP7_75t_SL g567 ( .A(n_420), .Y(n_567) );
BUFx2_ASAP7_75t_L g627 ( .A(n_420), .Y(n_627) );
BUFx3_ASAP7_75t_L g656 ( .A(n_420), .Y(n_656) );
BUFx2_ASAP7_75t_SL g1035 ( .A(n_420), .Y(n_1035) );
AND2x2_ASAP7_75t_L g543 ( .A(n_421), .B(n_514), .Y(n_543) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x6_ASAP7_75t_L g455 ( .A(n_422), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx5_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_427), .A2(n_435), .B1(n_570), .B2(n_571), .Y(n_569) );
INVx4_ASAP7_75t_L g711 ( .A(n_427), .Y(n_711) );
INVx2_ASAP7_75t_SL g734 ( .A(n_427), .Y(n_734) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_427), .Y(n_943) );
INVx2_ASAP7_75t_L g975 ( .A(n_427), .Y(n_975) );
INVx11_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx11_ASAP7_75t_L g534 ( .A(n_428), .Y(n_534) );
AND2x6_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
AND2x4_ASAP7_75t_L g486 ( .A(n_429), .B(n_447), .Y(n_486) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g500 ( .A(n_430), .B(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g436 ( .A(n_431), .B(n_437), .Y(n_436) );
AND2x6_ASAP7_75t_L g461 ( .A(n_431), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g716 ( .A(n_435), .Y(n_716) );
INVx3_ASAP7_75t_L g758 ( .A(n_435), .Y(n_758) );
INVx2_ASAP7_75t_L g807 ( .A(n_435), .Y(n_807) );
INVx6_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx3_ASAP7_75t_L g535 ( .A(n_436), .Y(n_535) );
BUFx3_ASAP7_75t_L g681 ( .A(n_436), .Y(n_681) );
BUFx3_ASAP7_75t_L g796 ( .A(n_436), .Y(n_796) );
AND2x6_ASAP7_75t_L g489 ( .A(n_437), .B(n_447), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g504 ( .A(n_437), .B(n_447), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_448), .Y(n_438) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx3_ASAP7_75t_L g574 ( .A(n_441), .Y(n_574) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_441), .Y(n_634) );
BUFx3_ASAP7_75t_L g839 ( .A(n_441), .Y(n_839) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g522 ( .A(n_442), .Y(n_522) );
BUFx2_ASAP7_75t_SL g803 ( .A(n_442), .Y(n_803) );
BUFx2_ASAP7_75t_SL g868 ( .A(n_442), .Y(n_868) );
INVx4_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx3_ASAP7_75t_L g626 ( .A(n_444), .Y(n_626) );
INVx4_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g523 ( .A(n_446), .Y(n_523) );
BUFx3_ASAP7_75t_L g566 ( .A(n_446), .Y(n_566) );
BUFx3_ASAP7_75t_L g644 ( .A(n_446), .Y(n_644) );
INVx2_ASAP7_75t_L g919 ( .A(n_446), .Y(n_919) );
INVx1_ASAP7_75t_L g501 ( .A(n_447), .Y(n_501) );
INVx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_L g900 ( .A(n_451), .Y(n_900) );
BUFx2_ASAP7_75t_L g1001 ( .A(n_451), .Y(n_1001) );
INVx4_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx5_ASAP7_75t_L g525 ( .A(n_452), .Y(n_525) );
BUFx3_ASAP7_75t_L g630 ( .A(n_452), .Y(n_630) );
INVx3_ASAP7_75t_L g642 ( .A(n_452), .Y(n_642) );
INVx2_ASAP7_75t_L g717 ( .A(n_452), .Y(n_717) );
INVx1_ASAP7_75t_L g871 ( .A(n_452), .Y(n_871) );
INVx8_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx6_ASAP7_75t_SL g527 ( .A(n_455), .Y(n_527) );
INVx1_ASAP7_75t_SL g631 ( .A(n_455), .Y(n_631) );
INVx1_ASAP7_75t_L g789 ( .A(n_455), .Y(n_789) );
INVx1_ASAP7_75t_L g479 ( .A(n_456), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_475), .Y(n_457) );
OAI222xp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_463), .B1(n_464), .B2(n_470), .C1(n_471), .C2(n_474), .Y(n_458) );
INVx2_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g609 ( .A(n_460), .Y(n_609) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx3_ASAP7_75t_L g510 ( .A(n_461), .Y(n_510) );
INVx4_ASAP7_75t_L g547 ( .A(n_461), .Y(n_547) );
INVx2_ASAP7_75t_L g666 ( .A(n_461), .Y(n_666) );
INVx2_ASAP7_75t_SL g1022 ( .A(n_461), .Y(n_1022) );
INVx2_ASAP7_75t_L g1042 ( .A(n_461), .Y(n_1042) );
AND2x4_ASAP7_75t_L g481 ( .A(n_462), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g517 ( .A(n_462), .Y(n_517) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g958 ( .A(n_465), .Y(n_958) );
BUFx4f_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_466), .Y(n_507) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_466), .Y(n_651) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_466), .Y(n_673) );
BUFx2_ASAP7_75t_L g704 ( .A(n_466), .Y(n_704) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g473 ( .A(n_468), .Y(n_473) );
AND2x4_ASAP7_75t_L g472 ( .A(n_469), .B(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g478 ( .A(n_469), .B(n_479), .Y(n_478) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_469), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx12f_ASAP7_75t_L g508 ( .A(n_472), .Y(n_508) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_472), .Y(n_549) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_472), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_483), .Y(n_475) );
BUFx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g590 ( .A(n_478), .Y(n_590) );
BUFx3_ASAP7_75t_L g652 ( .A(n_478), .Y(n_652) );
BUFx2_ASAP7_75t_L g751 ( .A(n_478), .Y(n_751) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_481), .Y(n_550) );
BUFx2_ASAP7_75t_SL g591 ( .A(n_481), .Y(n_591) );
BUFx2_ASAP7_75t_SL g746 ( .A(n_481), .Y(n_746) );
INVx1_ASAP7_75t_L g518 ( .A(n_482), .Y(n_518) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx5_ASAP7_75t_L g553 ( .A(n_485), .Y(n_553) );
INVx2_ASAP7_75t_L g648 ( .A(n_485), .Y(n_648) );
INVx2_ASAP7_75t_L g670 ( .A(n_485), .Y(n_670) );
INVx4_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_SL g857 ( .A(n_488), .Y(n_857) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g586 ( .A(n_489), .Y(n_586) );
BUFx2_ASAP7_75t_L g617 ( .A(n_489), .Y(n_617) );
BUFx4f_ASAP7_75t_L g649 ( .A(n_489), .Y(n_649) );
INVx1_ASAP7_75t_L g596 ( .A(n_491), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_536), .B1(n_594), .B2(n_595), .Y(n_491) );
INVx2_ASAP7_75t_SL g594 ( .A(n_492), .Y(n_594) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND3x1_ASAP7_75t_L g495 ( .A(n_496), .B(n_519), .C(n_528), .Y(n_495) );
NOR3xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_505), .C(n_511), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B1(n_502), .B2(n_503), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_499), .A2(n_695), .B1(n_773), .B2(n_774), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_499), .A2(n_695), .B1(n_923), .B2(n_924), .Y(n_922) );
BUFx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_500), .A2(n_693), .B1(n_694), .B2(n_695), .Y(n_692) );
INVx2_ASAP7_75t_L g881 ( .A(n_500), .Y(n_881) );
BUFx6f_ASAP7_75t_L g1015 ( .A(n_500), .Y(n_1015) );
INVx2_ASAP7_75t_L g884 ( .A(n_503), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_503), .A2(n_954), .B1(n_955), .B2(n_956), .Y(n_953) );
OAI22xp5_ASAP7_75t_SL g1014 ( .A1(n_503), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g696 ( .A(n_504), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_509), .Y(n_505) );
INVx4_ASAP7_75t_L g613 ( .A(n_507), .Y(n_613) );
BUFx2_ASAP7_75t_L g986 ( .A(n_507), .Y(n_986) );
BUFx4f_ASAP7_75t_SL g583 ( .A(n_508), .Y(n_583) );
INVx2_ASAP7_75t_L g660 ( .A(n_508), .Y(n_660) );
INVx3_ASAP7_75t_L g699 ( .A(n_510), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B1(n_515), .B2(n_516), .Y(n_511) );
INVx4_ASAP7_75t_L g707 ( .A(n_513), .Y(n_707) );
BUFx3_ASAP7_75t_L g822 ( .A(n_513), .Y(n_822) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_513), .Y(n_892) );
CKINVDCx16_ASAP7_75t_R g780 ( .A(n_516), .Y(n_780) );
BUFx2_ASAP7_75t_L g966 ( .A(n_516), .Y(n_966) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_524), .Y(n_519) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx3_ASAP7_75t_L g713 ( .A(n_522), .Y(n_713) );
BUFx6f_ASAP7_75t_L g788 ( .A(n_525), .Y(n_788) );
BUFx2_ASAP7_75t_L g1128 ( .A(n_525), .Y(n_1128) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g645 ( .A(n_527), .Y(n_645) );
BUFx4f_ASAP7_75t_SL g818 ( .A(n_527), .Y(n_818) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_532), .Y(n_528) );
BUFx2_ASAP7_75t_L g797 ( .A(n_530), .Y(n_797) );
INVx4_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_SL g784 ( .A(n_534), .Y(n_784) );
INVx3_ASAP7_75t_L g811 ( .A(n_534), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g1093 ( .A(n_534), .B(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g595 ( .A(n_536), .Y(n_595) );
OA22x2_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B1(n_561), .B2(n_593), .Y(n_536) );
OAI22x1_ASAP7_75t_L g738 ( .A1(n_537), .A2(n_538), .B1(n_739), .B2(n_760), .Y(n_738) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
XOR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_560), .Y(n_538) );
NAND3x1_ASAP7_75t_SL g539 ( .A(n_540), .B(n_544), .C(n_556), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_545), .B(n_551), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_548), .Y(n_545) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_547), .A2(n_581), .B(n_582), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_547), .A2(n_726), .B(n_727), .Y(n_725) );
OAI21xp5_ASAP7_75t_SL g742 ( .A1(n_547), .A2(n_743), .B(n_744), .Y(n_742) );
INVx4_ASAP7_75t_L g825 ( .A(n_547), .Y(n_825) );
BUFx2_ASAP7_75t_L g861 ( .A(n_547), .Y(n_861) );
OAI21xp5_ASAP7_75t_SL g991 ( .A1(n_547), .A2(n_992), .B(n_993), .Y(n_991) );
BUFx4f_ASAP7_75t_L g614 ( .A(n_549), .Y(n_614) );
INVx1_ASAP7_75t_SL g623 ( .A(n_550), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .C(n_555), .Y(n_551) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_553), .Y(n_619) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx2_ASAP7_75t_L g786 ( .A(n_559), .Y(n_786) );
INVx1_ASAP7_75t_L g593 ( .A(n_561), .Y(n_593) );
XOR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_592), .Y(n_561) );
AND2x2_ASAP7_75t_SL g562 ( .A(n_563), .B(n_579), .Y(n_562) );
NOR3xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_569), .C(n_572), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_568), .Y(n_564) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_566), .Y(n_1088) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_575), .B2(n_576), .Y(n_572) );
INVx2_ASAP7_75t_L g898 ( .A(n_574), .Y(n_898) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g809 ( .A(n_577), .Y(n_809) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_584), .Y(n_579) );
INVx1_ASAP7_75t_L g964 ( .A(n_583), .Y(n_964) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .C(n_588), .Y(n_584) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g621 ( .A(n_590), .Y(n_621) );
OAI22xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_599), .B1(n_686), .B2(n_687), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_637), .B2(n_638), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g636 ( .A(n_606), .Y(n_636) );
NAND3x1_ASAP7_75t_L g606 ( .A(n_607), .B(n_624), .C(n_632), .Y(n_606) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_608), .B(n_615), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_610), .B(n_611), .Y(n_608) );
OAI21xp5_ASAP7_75t_SL g1079 ( .A1(n_609), .A2(n_1080), .B(n_1081), .Y(n_1079) );
INVx1_ASAP7_75t_L g1113 ( .A(n_612), .Y(n_1113) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g1024 ( .A(n_614), .Y(n_1024) );
NAND3xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .C(n_620), .Y(n_615) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_628), .Y(n_624) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
AO22x2_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_661), .B1(n_684), .B2(n_685), .Y(n_638) );
INVx1_ASAP7_75t_L g684 ( .A(n_639), .Y(n_684) );
NAND5xp2_ASAP7_75t_SL g640 ( .A(n_641), .B(n_643), .C(n_646), .D(n_653), .E(n_658), .Y(n_640) );
BUFx2_ASAP7_75t_L g792 ( .A(n_644), .Y(n_792) );
AND2x2_ASAP7_75t_SL g646 ( .A(n_647), .B(n_650), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_651), .Y(n_769) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_657), .Y(n_653) );
BUFx3_ASAP7_75t_L g915 ( .A(n_655), .Y(n_915) );
INVx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g685 ( .A(n_661), .Y(n_685) );
XOR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_683), .Y(n_661) );
NAND2x1p5_ASAP7_75t_L g662 ( .A(n_663), .B(n_674), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_668), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B(n_667), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g767 ( .A1(n_666), .A2(n_768), .B1(n_769), .B2(n_770), .C(n_771), .Y(n_767) );
OAI221xp5_ASAP7_75t_L g885 ( .A1(n_666), .A2(n_886), .B1(n_887), .B2(n_888), .C(n_889), .Y(n_885) );
OAI222xp33_ASAP7_75t_L g957 ( .A1(n_666), .A2(n_706), .B1(n_958), .B2(n_959), .C1(n_960), .C2(n_961), .Y(n_957) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .C(n_672), .Y(n_668) );
BUFx6f_ASAP7_75t_L g1020 ( .A(n_673), .Y(n_1020) );
NOR2x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_679), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
INVx3_ASAP7_75t_L g945 ( .A(n_681), .Y(n_945) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_737), .B1(n_738), .B2(n_761), .Y(n_687) );
INVx2_ASAP7_75t_L g761 ( .A(n_688), .Y(n_761) );
XOR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_719), .Y(n_688) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_708), .Y(n_690) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_697), .C(n_701), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g979 ( .A(n_696), .Y(n_979) );
OAI21xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B(n_700), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_705), .B2(n_706), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx3_ASAP7_75t_SL g777 ( .A(n_707), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_714), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_718), .Y(n_714) );
OAI22xp5_ASAP7_75t_SL g849 ( .A1(n_719), .A2(n_850), .B1(n_851), .B2(n_874), .Y(n_849) );
INVx2_ASAP7_75t_L g874 ( .A(n_719), .Y(n_874) );
XOR2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_736), .Y(n_719) );
NAND3x1_ASAP7_75t_L g720 ( .A(n_721), .B(n_724), .C(n_732), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NOR2x1_ASAP7_75t_L g724 ( .A(n_725), .B(n_728), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .C(n_731), .Y(n_728) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g1126 ( .A(n_734), .Y(n_1126) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g760 ( .A(n_739), .Y(n_760) );
AND2x4_ASAP7_75t_L g740 ( .A(n_741), .B(n_752), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_747), .Y(n_741) );
BUFx3_ASAP7_75t_L g826 ( .A(n_745), .Y(n_826) );
BUFx2_ASAP7_75t_L g929 ( .A(n_745), .Y(n_929) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .C(n_750), .Y(n_747) );
NOR2x1_ASAP7_75t_L g752 ( .A(n_753), .B(n_756), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_759), .Y(n_756) );
XNOR2x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_831), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_800), .B1(n_829), .B2(n_830), .Y(n_763) );
INVx1_ASAP7_75t_L g829 ( .A(n_764), .Y(n_829) );
INVx2_ASAP7_75t_SL g799 ( .A(n_765), .Y(n_799) );
AND2x4_ASAP7_75t_L g765 ( .A(n_766), .B(n_781), .Y(n_765) );
NOR3xp33_ASAP7_75t_SL g766 ( .A(n_767), .B(n_772), .C(n_775), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g925 ( .A1(n_769), .A2(n_861), .B1(n_926), .B2(n_927), .C(n_928), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_777), .A2(n_894), .B1(n_931), .B2(n_932), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_779), .A2(n_821), .B1(n_822), .B2(n_823), .Y(n_820) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g894 ( .A(n_780), .Y(n_894) );
NOR2x1_ASAP7_75t_L g781 ( .A(n_782), .B(n_790), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_787), .Y(n_782) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g830 ( .A(n_800), .Y(n_830) );
INVx1_ASAP7_75t_L g828 ( .A(n_801), .Y(n_828) );
AND4x1_ASAP7_75t_L g801 ( .A(n_802), .B(n_810), .C(n_819), .D(n_824), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_808), .B2(n_809), .Y(n_804) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_814), .B1(n_816), .B2(n_817), .Y(n_812) );
OAI21xp33_ASAP7_75t_L g1090 ( .A1(n_814), .A2(n_1091), .B(n_1092), .Y(n_1090) );
BUFx2_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
OAI22xp5_ASAP7_75t_SL g1026 ( .A1(n_822), .A2(n_894), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_822), .A2(n_966), .B1(n_1117), .B2(n_1118), .Y(n_1116) );
INVx2_ASAP7_75t_L g887 ( .A(n_826), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_847), .B1(n_905), .B2(n_906), .Y(n_831) );
INVx2_ASAP7_75t_L g905 ( .A(n_832), .Y(n_905) );
NAND4xp75_ASAP7_75t_L g833 ( .A(n_834), .B(n_837), .C(n_843), .D(n_846), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
AND2x2_ASAP7_75t_L g837 ( .A(n_838), .B(n_842), .Y(n_837) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
AND2x2_ASAP7_75t_SL g843 ( .A(n_844), .B(n_845), .Y(n_843) );
INVx1_ASAP7_75t_L g906 ( .A(n_847), .Y(n_906) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B1(n_875), .B2(n_904), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx2_ASAP7_75t_SL g873 ( .A(n_853), .Y(n_873) );
NAND2x1p5_ASAP7_75t_L g853 ( .A(n_854), .B(n_864), .Y(n_853) );
NOR2xp67_ASAP7_75t_SL g854 ( .A(n_855), .B(n_860), .Y(n_854) );
NAND3xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_858), .C(n_859), .Y(n_855) );
OAI21xp5_ASAP7_75t_SL g860 ( .A1(n_861), .A2(n_862), .B(n_863), .Y(n_860) );
OAI221xp5_ASAP7_75t_L g1111 ( .A1(n_861), .A2(n_1112), .B1(n_1113), .B2(n_1114), .C(n_1115), .Y(n_1111) );
NOR2x1_ASAP7_75t_L g864 ( .A(n_865), .B(n_869), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_872), .Y(n_869) );
INVx2_ASAP7_75t_L g904 ( .A(n_875), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_877), .B(n_895), .Y(n_876) );
NOR3xp33_ASAP7_75t_L g877 ( .A(n_878), .B(n_885), .C(n_890), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_880), .B1(n_882), .B2(n_883), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_880), .A2(n_883), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_SL g955 ( .A(n_881), .Y(n_955) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_892), .B1(n_893), .B2(n_894), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_901), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_897), .B(n_899), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_935), .B1(n_1058), .B2(n_1059), .Y(n_908) );
INVx1_ASAP7_75t_L g1059 ( .A(n_909), .Y(n_1059) );
INVx1_ASAP7_75t_SL g934 ( .A(n_910), .Y(n_934) );
AND2x2_ASAP7_75t_SL g910 ( .A(n_911), .B(n_921), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_916), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_917), .B(n_920), .Y(n_916) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NOR3xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_925), .C(n_930), .Y(n_921) );
INVx1_ASAP7_75t_L g1058 ( .A(n_935), .Y(n_1058) );
BUFx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
OAI22xp5_ASAP7_75t_SL g936 ( .A1(n_937), .A2(n_938), .B1(n_1007), .B2(n_1008), .Y(n_936) );
INVx2_ASAP7_75t_SL g937 ( .A(n_938), .Y(n_937) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_939), .A2(n_969), .B1(n_970), .B2(n_1006), .Y(n_938) );
INVx2_ASAP7_75t_L g1006 ( .A(n_939), .Y(n_1006) );
INVx1_ASAP7_75t_L g967 ( .A(n_940), .Y(n_967) );
AND2x2_ASAP7_75t_SL g940 ( .A(n_941), .B(n_952), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_942), .B(n_948), .Y(n_941) );
OAI221xp5_ASAP7_75t_SL g942 ( .A1(n_943), .A2(n_944), .B1(n_945), .B2(n_946), .C(n_947), .Y(n_942) );
NOR3xp33_ASAP7_75t_L g952 ( .A(n_953), .B(n_957), .C(n_962), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_963), .A2(n_964), .B1(n_965), .B2(n_966), .Y(n_962) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
XNOR2x2_ASAP7_75t_L g970 ( .A(n_971), .B(n_988), .Y(n_970) );
XOR2x2_ASAP7_75t_L g971 ( .A(n_972), .B(n_987), .Y(n_971) );
NAND4xp75_ASAP7_75t_L g972 ( .A(n_973), .B(n_977), .C(n_982), .D(n_985), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_974), .B(n_976), .Y(n_973) );
OA211x2_ASAP7_75t_L g977 ( .A1(n_978), .A2(n_979), .B(n_980), .C(n_981), .Y(n_977) );
AND2x2_ASAP7_75t_L g982 ( .A(n_983), .B(n_984), .Y(n_982) );
XOR2x2_ASAP7_75t_L g988 ( .A(n_989), .B(n_1005), .Y(n_988) );
NAND3x1_ASAP7_75t_L g989 ( .A(n_990), .B(n_998), .C(n_1002), .Y(n_989) );
NOR2x1_ASAP7_75t_L g990 ( .A(n_991), .B(n_994), .Y(n_990) );
NAND3xp33_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .C(n_997), .Y(n_994) );
AND2x2_ASAP7_75t_L g998 ( .A(n_999), .B(n_1000), .Y(n_998) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1004), .Y(n_1002) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
AOI22xp5_ASAP7_75t_L g1009 ( .A1(n_1010), .A2(n_1037), .B1(n_1056), .B2(n_1057), .Y(n_1009) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1010), .Y(n_1056) );
XNOR2x2_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1029), .Y(n_1012) );
NOR3xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1018), .C(n_1026), .Y(n_1013) );
OAI222xp33_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1021), .B1(n_1022), .B2(n_1023), .C1(n_1024), .C2(n_1025), .Y(n_1018) );
INVx2_ASAP7_75t_SL g1019 ( .A(n_1020), .Y(n_1019) );
NOR2xp33_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1033), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1032), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1036), .Y(n_1033) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1037), .Y(n_1057) );
INVx2_ASAP7_75t_L g1055 ( .A(n_1039), .Y(n_1055) );
NAND2x1_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1048), .Y(n_1039) );
NOR2xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1045), .Y(n_1040) );
OAI21xp5_ASAP7_75t_SL g1041 ( .A1(n_1042), .A2(n_1043), .B(n_1044), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1047), .Y(n_1045) );
NOR2x1_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1052), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1051), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1054), .Y(n_1052) );
INVx1_ASAP7_75t_SL g1061 ( .A(n_1062), .Y(n_1061) );
NOR2x1_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1067), .Y(n_1062) );
OR2x2_ASAP7_75t_SL g1132 ( .A(n_1063), .B(n_1068), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1066), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g1096 ( .A(n_1065), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_1065), .B(n_1100), .Y(n_1103) );
CKINVDCx16_ASAP7_75t_R g1100 ( .A(n_1066), .Y(n_1100) );
CKINVDCx20_ASAP7_75t_R g1067 ( .A(n_1068), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1070), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1073), .Y(n_1071) );
OAI322xp33_ASAP7_75t_L g1074 ( .A1(n_1075), .A2(n_1096), .A3(n_1097), .B1(n_1101), .B2(n_1104), .C1(n_1105), .C2(n_1130), .Y(n_1074) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
NAND3x1_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1085), .C(n_1089), .Y(n_1077) );
NOR2xp33_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1082), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1084), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1087), .Y(n_1085) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1106), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1119), .Y(n_1106) );
NOR3xp33_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1111), .C(n_1116), .Y(n_1107) );
NOR2xp67_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1123), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1122), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1127), .Y(n_1123) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
CKINVDCx20_ASAP7_75t_R g1130 ( .A(n_1131), .Y(n_1130) );
CKINVDCx20_ASAP7_75t_R g1131 ( .A(n_1132), .Y(n_1131) );
endmodule