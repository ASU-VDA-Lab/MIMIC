module fake_jpeg_15783_n_236 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_19),
.Y(n_29)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_28),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_44),
.B(n_49),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_31),
.Y(n_45)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_34),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_30),
.Y(n_73)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_21),
.B1(n_18),
.B2(n_25),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_35),
.B1(n_37),
.B2(n_29),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_32),
.B1(n_21),
.B2(n_20),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_70),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_37),
.B1(n_29),
.B2(n_30),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_32),
.C(n_29),
.Y(n_72)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_28),
.CI(n_41),
.CON(n_86),
.SN(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_30),
.B1(n_36),
.B2(n_38),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_77),
.A2(n_92),
.B1(n_41),
.B2(n_39),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_72),
.B(n_59),
.C(n_16),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_69),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_28),
.B1(n_42),
.B2(n_36),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_60),
.B(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_93),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_56),
.B1(n_43),
.B2(n_49),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_105),
.B1(n_113),
.B2(n_41),
.Y(n_126)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

AND2x4_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_66),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_43),
.B1(n_54),
.B2(n_45),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_114),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g107 ( 
.A(n_94),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_57),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_116),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_40),
.B1(n_66),
.B2(n_70),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_78),
.B1(n_83),
.B2(n_93),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_36),
.B(n_66),
.C(n_60),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_40),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_15),
.B(n_23),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_15),
.B(n_24),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_17),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_118),
.B1(n_111),
.B2(n_92),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_87),
.B1(n_86),
.B2(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_127),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_111),
.B1(n_97),
.B2(n_112),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_101),
.C(n_79),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_26),
.C(n_22),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_82),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_134),
.B(n_136),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_14),
.B1(n_24),
.B2(n_27),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_27),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_151),
.B(n_135),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_145),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_105),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_153),
.C(n_154),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_113),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_155),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_130),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_148),
.B1(n_156),
.B2(n_34),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_111),
.B1(n_107),
.B2(n_100),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_90),
.B1(n_85),
.B2(n_76),
.Y(n_149)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_33),
.B(n_17),
.C(n_39),
.D(n_26),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_33),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_17),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_34),
.B1(n_96),
.B2(n_68),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_120),
.CI(n_122),
.CON(n_161),
.SN(n_161)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_131),
.B(n_120),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_165),
.B1(n_166),
.B2(n_170),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_169),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_152),
.A2(n_127),
.B1(n_131),
.B2(n_119),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_119),
.B(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_153),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_180),
.C(n_184),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_162),
.A2(n_144),
.B1(n_154),
.B2(n_155),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_159),
.B1(n_14),
.B2(n_2),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_96),
.C(n_55),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_26),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_26),
.C(n_22),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_170),
.B1(n_168),
.B2(n_157),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_161),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_175),
.B(n_187),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_177),
.B(n_172),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_196),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_173),
.C(n_163),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_198),
.C(n_200),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_183),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_0),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_1),
.C(n_2),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_179),
.B(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_207),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_174),
.A3(n_184),
.B1(n_13),
.B2(n_12),
.C1(n_6),
.C2(n_7),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_4),
.B(n_6),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_210),
.C(n_201),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_12),
.C(n_5),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_193),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_212),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_8),
.B(n_9),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_219),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_204),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_217),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_211),
.A2(n_189),
.B(n_192),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_7),
.B(n_8),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_195),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_208),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_223),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_9),
.B(n_10),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_212),
.B(n_213),
.C(n_11),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g230 ( 
.A(n_227),
.Y(n_230)
);

NOR3x1_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_9),
.C(n_10),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_228),
.A2(n_229),
.B1(n_10),
.B2(n_11),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_230),
.A2(n_225),
.B(n_226),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_38),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_233),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_38),
.Y(n_236)
);


endmodule