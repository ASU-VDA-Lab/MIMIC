module fake_ariane_98_n_9276 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_106, n_12, n_53, n_111, n_21, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_112, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_108, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_9276);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_112;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_108;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_9276;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_7329;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_8165;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_8139;
wire n_416;
wire n_4962;
wire n_1430;
wire n_7832;
wire n_8438;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_8321;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_7922;
wire n_7805;
wire n_2790;
wire n_7542;
wire n_2207;
wire n_7053;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_462;
wire n_8699;
wire n_9263;
wire n_1131;
wire n_8037;
wire n_5479;
wire n_2646;
wire n_8257;
wire n_737;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_232;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_9096;
wire n_6358;
wire n_8546;
wire n_6293;
wire n_8997;
wire n_2482;
wire n_1682;
wire n_7001;
wire n_958;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_146;
wire n_9241;
wire n_4853;
wire n_8744;
wire n_338;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_7464;
wire n_8449;
wire n_4260;
wire n_903;
wire n_7626;
wire n_3348;
wire n_239;
wire n_3261;
wire n_1761;
wire n_8953;
wire n_7965;
wire n_7368;
wire n_1690;
wire n_8399;
wire n_2807;
wire n_6664;
wire n_8598;
wire n_7562;
wire n_7534;
wire n_1018;
wire n_7428;
wire n_4512;
wire n_6190;
wire n_8460;
wire n_4132;
wire n_1364;
wire n_7373;
wire n_2390;
wire n_8068;
wire n_6891;
wire n_4500;
wire n_625;
wire n_2322;
wire n_8734;
wire n_1107;
wire n_8720;
wire n_331;
wire n_559;
wire n_2663;
wire n_8097;
wire n_5481;
wire n_6539;
wire n_495;
wire n_8114;
wire n_8422;
wire n_4824;
wire n_7467;
wire n_350;
wire n_8126;
wire n_381;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_7526;
wire n_8664;
wire n_561;
wire n_4143;
wire n_4273;
wire n_507;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_786;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_9119;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_9058;
wire n_6197;
wire n_7200;
wire n_8326;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_8504;
wire n_3015;
wire n_5744;
wire n_8920;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_277;
wire n_5691;
wire n_7937;
wire n_8985;
wire n_3482;
wire n_7490;
wire n_6295;
wire n_5403;
wire n_823;
wire n_1900;
wire n_620;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_587;
wire n_863;
wire n_6992;
wire n_303;
wire n_3960;
wire n_2433;
wire n_352;
wire n_899;
wire n_3975;
wire n_8035;
wire n_5830;
wire n_365;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_8660;
wire n_334;
wire n_192;
wire n_3325;
wire n_6681;
wire n_661;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_8939;
wire n_533;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_6542;
wire n_9202;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_273;
wire n_4505;
wire n_6452;
wire n_1840;
wire n_5247;
wire n_8469;
wire n_8715;
wire n_5464;
wire n_7306;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_579;
wire n_7507;
wire n_844;
wire n_1267;
wire n_8176;
wire n_2956;
wire n_5210;
wire n_7441;
wire n_149;
wire n_1213;
wire n_2382;
wire n_7379;
wire n_7215;
wire n_237;
wire n_780;
wire n_5292;
wire n_1918;
wire n_8327;
wire n_8991;
wire n_7438;
wire n_8855;
wire n_4443;
wire n_4119;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_3458;
wire n_570;
wire n_5843;
wire n_7874;
wire n_8539;
wire n_8630;
wire n_8533;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_490;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_575;
wire n_8435;
wire n_7695;
wire n_6156;
wire n_1216;
wire n_4908;
wire n_8098;
wire n_3754;
wire n_8204;
wire n_5060;
wire n_9199;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_7331;
wire n_5913;
wire n_8958;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_7944;
wire n_3841;
wire n_5249;
wire n_249;
wire n_851;
wire n_123;
wire n_444;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_9265;
wire n_6872;
wire n_6644;
wire n_9143;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_8542;
wire n_8572;
wire n_5046;
wire n_7607;
wire n_7642;
wire n_8373;
wire n_8424;
wire n_8442;
wire n_1386;
wire n_6236;
wire n_7104;
wire n_8147;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_1842;
wire n_4993;
wire n_7397;
wire n_3678;
wire n_7205;
wire n_366;
wire n_2791;
wire n_1661;
wire n_555;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_7461;
wire n_8519;
wire n_1692;
wire n_2611;
wire n_8075;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_7638;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_8642;
wire n_8648;
wire n_7224;
wire n_6966;
wire n_5056;
wire n_9149;
wire n_1178;
wire n_2015;
wire n_7259;
wire n_7838;
wire n_8556;
wire n_5984;
wire n_5204;
wire n_6724;
wire n_6705;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_203;
wire n_4951;
wire n_8585;
wire n_3000;
wire n_150;
wire n_2930;
wire n_7840;
wire n_4959;
wire n_2745;
wire n_8455;
wire n_2087;
wire n_8444;
wire n_619;
wire n_9128;
wire n_2161;
wire n_746;
wire n_6624;
wire n_1357;
wire n_7888;
wire n_8560;
wire n_292;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_8108;
wire n_1389;
wire n_8158;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_6553;
wire n_4905;
wire n_9016;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_6261;
wire n_3651;
wire n_1812;
wire n_6659;
wire n_4894;
wire n_428;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_8814;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_7583;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_542;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_1087;
wire n_632;
wire n_9094;
wire n_2388;
wire n_2273;
wire n_8130;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_7488;
wire n_3700;
wire n_7690;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_6206;
wire n_7893;
wire n_2954;
wire n_382;
wire n_489;
wire n_4438;
wire n_6538;
wire n_7966;
wire n_251;
wire n_974;
wire n_506;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_7599;
wire n_7231;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_1447;
wire n_8675;
wire n_1220;
wire n_9095;
wire n_7900;
wire n_2019;
wire n_5708;
wire n_8123;
wire n_698;
wire n_9003;
wire n_9048;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_124;
wire n_5454;
wire n_307;
wire n_1209;
wire n_4254;
wire n_646;
wire n_8913;
wire n_3438;
wire n_8220;
wire n_404;
wire n_2625;
wire n_8355;
wire n_5373;
wire n_7403;
wire n_1578;
wire n_6665;
wire n_8883;
wire n_3147;
wire n_299;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_133;
wire n_1029;
wire n_2649;
wire n_6461;
wire n_6033;
wire n_1247;
wire n_6860;
wire n_9063;
wire n_522;
wire n_1568;
wire n_2919;
wire n_7322;
wire n_6060;
wire n_3108;
wire n_5983;
wire n_5788;
wire n_367;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_8816;
wire n_4314;
wire n_8418;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_3239;
wire n_2631;
wire n_9110;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_424;
wire n_4857;
wire n_8739;
wire n_8927;
wire n_1651;
wire n_3087;
wire n_7221;
wire n_6009;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_8243;
wire n_3704;
wire n_8798;
wire n_7963;
wire n_6382;
wire n_8423;
wire n_9028;
wire n_670;
wire n_2677;
wire n_4296;
wire n_379;
wire n_138;
wire n_162;
wire n_2483;
wire n_7938;
wire n_5088;
wire n_6615;
wire n_441;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_9270;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_8548;
wire n_8996;
wire n_207;
wire n_720;
wire n_6263;
wire n_1943;
wire n_8156;
wire n_6731;
wire n_5138;
wire n_8845;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_194;
wire n_5149;
wire n_9256;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_6234;
wire n_4153;
wire n_8992;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_8510;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_8961;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_8402;
wire n_8978;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_9105;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_8685;
wire n_1828;
wire n_9240;
wire n_1304;
wire n_7202;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_9212;
wire n_5985;
wire n_8595;
wire n_604;
wire n_478;
wire n_9040;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_7868;
wire n_3370;
wire n_874;
wire n_7654;
wire n_3949;
wire n_2286;
wire n_8779;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_129;
wire n_126;
wire n_3036;
wire n_2783;
wire n_8520;
wire n_4583;
wire n_8555;
wire n_6366;
wire n_1015;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_9146;
wire n_688;
wire n_7176;
wire n_636;
wire n_8565;
wire n_8334;
wire n_1490;
wire n_6074;
wire n_7547;
wire n_5552;
wire n_442;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_8030;
wire n_8513;
wire n_887;
wire n_9219;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_2861;
wire n_8245;
wire n_7942;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_8753;
wire n_1498;
wire n_1188;
wire n_7527;
wire n_4856;
wire n_2618;
wire n_7948;
wire n_7096;
wire n_4216;
wire n_957;
wire n_1242;
wire n_9206;
wire n_2707;
wire n_8485;
wire n_5596;
wire n_6482;
wire n_8106;
wire n_2849;
wire n_1489;
wire n_8325;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_616;
wire n_7293;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_9082;
wire n_7144;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_7316;
wire n_7508;
wire n_3070;
wire n_1005;
wire n_8677;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_4182;
wire n_2452;
wire n_8626;
wire n_2827;
wire n_7869;
wire n_3214;
wire n_8166;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_6631;
wire n_5889;
wire n_8602;
wire n_7151;
wire n_3944;
wire n_7762;
wire n_5632;
wire n_4729;
wire n_8002;
wire n_6728;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_7472;
wire n_4800;
wire n_1373;
wire n_7075;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_7611;
wire n_7796;
wire n_6508;
wire n_832;
wire n_7989;
wire n_8047;
wire n_744;
wire n_2821;
wire n_3696;
wire n_9233;
wire n_7936;
wire n_215;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_655;
wire n_4237;
wire n_8751;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_8800;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_2211;
wire n_8955;
wire n_951;
wire n_8039;
wire n_8193;
wire n_9073;
wire n_7546;
wire n_8432;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_8684;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_722;
wire n_7407;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_8628;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_7481;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_5435;
wire n_6484;
wire n_3340;
wire n_7182;
wire n_5053;
wire n_5476;
wire n_5483;
wire n_8617;
wire n_7605;
wire n_8591;
wire n_8090;
wire n_1243;
wire n_9268;
wire n_5511;
wire n_8661;
wire n_3486;
wire n_6639;
wire n_358;
wire n_608;
wire n_9187;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_317;
wire n_3197;
wire n_7423;
wire n_3256;
wire n_1878;
wire n_7375;
wire n_7076;
wire n_7689;
wire n_6344;
wire n_8189;
wire n_8811;
wire n_266;
wire n_7736;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_7419;
wire n_811;
wire n_6600;
wire n_7010;
wire n_791;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_8192;
wire n_9251;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_8573;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_480;
wire n_7918;
wire n_642;
wire n_1406;
wire n_6555;
wire n_5073;
wire n_4306;
wire n_6360;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_9181;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_474;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_8339;
wire n_386;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_197;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_7346;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_8775;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_1657;
wire n_8804;
wire n_6650;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_7385;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_9250;
wire n_1330;
wire n_906;
wire n_6204;
wire n_2295;
wire n_5225;
wire n_283;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_7148;
wire n_3142;
wire n_9171;
wire n_7169;
wire n_3129;
wire n_374;
wire n_3495;
wire n_3843;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_7600;
wire n_9124;
wire n_2386;
wire n_5826;
wire n_8697;
wire n_4822;
wire n_6946;
wire n_7947;
wire n_8645;
wire n_5931;
wire n_8820;
wire n_8146;
wire n_1829;
wire n_4635;
wire n_7847;
wire n_8154;
wire n_1450;
wire n_5532;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_8027;
wire n_7807;
wire n_1493;
wire n_2911;
wire n_515;
wire n_8063;
wire n_3313;
wire n_8406;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_8480;
wire n_4419;
wire n_8849;
wire n_5405;
wire n_7660;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_6442;
wire n_8241;
wire n_140;
wire n_6188;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_230;
wire n_3548;
wire n_4906;
wire n_6846;
wire n_4630;
wire n_8261;
wire n_6840;
wire n_142;
wire n_6645;
wire n_8535;
wire n_8348;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_7831;
wire n_8138;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_8702;
wire n_1995;
wire n_7455;
wire n_8273;
wire n_1397;
wire n_5921;
wire n_6247;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_8235;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_8294;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_9036;
wire n_9165;
wire n_7509;
wire n_6205;
wire n_2506;
wire n_8349;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_7497;
wire n_7315;
wire n_8429;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_7887;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_8486;
wire n_9052;
wire n_2070;
wire n_426;
wire n_6706;
wire n_7431;
wire n_8140;
wire n_398;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_166;
wire n_8117;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_7521;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_8129;
wire n_1291;
wire n_7253;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_7569;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_6551;
wire n_3386;
wire n_400;
wire n_7972;
wire n_8672;
wire n_7505;
wire n_3921;
wire n_282;
wire n_467;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_7524;
wire n_4196;
wire n_1197;
wire n_8934;
wire n_7318;
wire n_2613;
wire n_7411;
wire n_7326;
wire n_5667;
wire n_168;
wire n_1517;
wire n_2647;
wire n_8847;
wire n_8005;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_9030;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_8221;
wire n_7573;
wire n_6630;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_8191;
wire n_6798;
wire n_5999;
wire n_1504;
wire n_2110;
wire n_7498;
wire n_7895;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_8225;
wire n_3822;
wire n_889;
wire n_4355;
wire n_7453;
wire n_3818;
wire n_7932;
wire n_7890;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6403;
wire n_3497;
wire n_6395;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_565;
wire n_3927;
wire n_6141;
wire n_8559;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_8689;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_452;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_8330;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_6944;
wire n_4452;
wire n_284;
wire n_3887;
wire n_3195;
wire n_8304;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_8163;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_7240;
wire n_8907;
wire n_409;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_1056;
wire n_526;
wire n_5584;
wire n_674;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_6559;
wire n_4088;
wire n_9038;
wire n_8777;
wire n_2669;
wire n_8698;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_6248;
wire n_6541;
wire n_9034;
wire n_848;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_629;
wire n_4733;
wire n_7927;
wire n_161;
wire n_8928;
wire n_1814;
wire n_7219;
wire n_2441;
wire n_8081;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_216;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_7402;
wire n_6351;
wire n_4509;
wire n_4935;
wire n_2073;
wire n_7382;
wire n_8384;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_8650;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_7767;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_3433;
wire n_2931;
wire n_8284;
wire n_8374;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_7510;
wire n_9041;
wire n_3786;
wire n_875;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_7434;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_9035;
wire n_9011;
wire n_1715;
wire n_4204;
wire n_7691;
wire n_296;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_9135;
wire n_6744;
wire n_3645;
wire n_793;
wire n_5705;
wire n_6927;
wire n_7335;
wire n_132;
wire n_4996;
wire n_9107;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_7735;
wire n_8531;
wire n_6116;
wire n_8074;
wire n_494;
wire n_3550;
wire n_8780;
wire n_7956;
wire n_5510;
wire n_7495;
wire n_7651;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_8580;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_185;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_8358;
wire n_972;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_164;
wire n_2843;
wire n_3714;
wire n_9093;
wire n_184;
wire n_7671;
wire n_4832;
wire n_8033;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_118;
wire n_1679;
wire n_5834;
wire n_7926;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_8643;
wire n_2356;
wire n_5618;
wire n_6495;
wire n_7528;
wire n_6209;
wire n_4672;
wire n_8094;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_7413;
wire n_7993;
wire n_7821;
wire n_160;
wire n_7620;
wire n_119;
wire n_1008;
wire n_3963;
wire n_581;
wire n_3091;
wire n_6274;
wire n_1024;
wire n_176;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_6237;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_7343;
wire n_5982;
wire n_8477;
wire n_1775;
wire n_908;
wire n_1036;
wire n_7109;
wire n_8028;
wire n_341;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_549;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_6809;
wire n_6099;
wire n_3225;
wire n_8530;
wire n_3621;
wire n_5529;
wire n_244;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_8500;
wire n_6716;
wire n_8713;
wire n_3565;
wire n_7885;
wire n_8297;
wire n_6905;
wire n_8926;
wire n_8456;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_5824;
wire n_8025;
wire n_5354;
wire n_2453;
wire n_7898;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_3040;
wire n_4230;
wire n_6899;
wire n_7980;
wire n_7817;
wire n_6413;
wire n_445;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_9025;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_8293;
wire n_3211;
wire n_7299;
wire n_917;
wire n_5196;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_8029;
wire n_2215;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_8880;
wire n_1261;
wire n_7249;
wire n_5763;
wire n_3633;
wire n_857;
wire n_363;
wire n_6061;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_8471;
wire n_1462;
wire n_5701;
wire n_7002;
wire n_1064;
wire n_633;
wire n_1446;
wire n_1701;
wire n_6273;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_8726;
wire n_731;
wire n_8977;
wire n_1813;
wire n_315;
wire n_2997;
wire n_7018;
wire n_1573;
wire n_6746;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_8316;
wire n_6174;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_5907;
wire n_784;
wire n_4339;
wire n_7297;
wire n_7730;
wire n_8134;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4169;
wire n_4024;
wire n_3316;
wire n_8610;
wire n_4023;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_3632;
wire n_309;
wire n_1344;
wire n_115;
wire n_485;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_435;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_840;
wire n_2324;
wire n_6575;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_2139;
wire n_7613;
wire n_9061;
wire n_7995;
wire n_8113;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_8724;
wire n_7140;
wire n_614;
wire n_4066;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_8253;
wire n_9258;
wire n_9228;
wire n_3303;
wire n_7910;
wire n_6592;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_248;
wire n_7741;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_228;
wire n_6668;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_8232;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_8803;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_8818;
wire n_7698;
wire n_1875;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_1150;
wire n_7800;
wire n_4266;
wire n_6336;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_7835;
wire n_1136;
wire n_458;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_7415;
wire n_8823;
wire n_5399;
wire n_8536;
wire n_658;
wire n_362;
wire n_8795;
wire n_2846;
wire n_3371;
wire n_8674;
wire n_9186;
wire n_4918;
wire n_5856;
wire n_8016;
wire n_3872;
wire n_5760;
wire n_7747;
wire n_4415;
wire n_5110;
wire n_8966;
wire n_1964;
wire n_3659;
wire n_7552;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_5844;
wire n_6298;
wire n_8132;
wire n_7650;
wire n_3441;
wire n_199;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_708;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_7635;
wire n_4408;
wire n_2115;
wire n_8567;
wire n_8259;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_6525;
wire n_3555;
wire n_5938;
wire n_7274;
wire n_3534;
wire n_450;
wire n_8578;
wire n_4548;
wire n_7819;
wire n_8495;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_896;
wire n_4574;
wire n_8160;
wire n_8980;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_8336;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_7788;
wire n_6974;
wire n_1168;
wire n_4663;
wire n_219;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_8600;
wire n_8229;
wire n_415;
wire n_4686;
wire n_9236;
wire n_2384;
wire n_7794;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_8761;
wire n_1846;
wire n_7630;
wire n_4161;
wire n_304;
wire n_9076;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6951;
wire n_6963;
wire n_1581;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_375;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_5355;
wire n_6284;
wire n_998;
wire n_3592;
wire n_5321;
wire n_7454;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_8473;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_8351;
wire n_5915;
wire n_7276;
wire n_174;
wire n_6379;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_925;
wire n_7753;
wire n_6834;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_8948;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_719;
wire n_7541;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_7913;
wire n_8020;
wire n_7946;
wire n_8944;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_9275;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_6471;
wire n_6949;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_6760;
wire n_2940;
wire n_548;
wire n_3427;
wire n_8875;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_9102;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_2491;
wire n_7920;
wire n_1931;
wire n_5559;
wire n_8649;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_1820;
wire n_7841;
wire n_7324;
wire n_7160;
wire n_8205;
wire n_6046;
wire n_7054;
wire n_1233;
wire n_4493;
wire n_8975;
wire n_6055;
wire n_7161;
wire n_9004;
wire n_1808;
wire n_6364;
wire n_8919;
wire n_6091;
wire n_6348;
wire n_1635;
wire n_8440;
wire n_1704;
wire n_4896;
wire n_8041;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_886;
wire n_7837;
wire n_359;
wire n_6788;
wire n_1308;
wire n_6144;
wire n_1451;
wire n_1487;
wire n_675;
wire n_9200;
wire n_5528;
wire n_7806;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_8076;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_8757;
wire n_1355;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_8897;
wire n_7676;
wire n_8177;
wire n_2334;
wire n_5467;
wire n_7241;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_9207;
wire n_1916;
wire n_6285;
wire n_610;
wire n_7644;
wire n_4602;
wire n_1713;
wire n_7816;
wire n_8829;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_7430;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_8638;
wire n_1515;
wire n_817;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_7269;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_9176;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_214;
wire n_4103;
wire n_2529;
wire n_8101;
wire n_2374;
wire n_5439;
wire n_8687;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_137;
wire n_8721;
wire n_1366;
wire n_8749;
wire n_3938;
wire n_8937;
wire n_2278;
wire n_7067;
wire n_6272;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_7879;
wire n_8730;
wire n_6607;
wire n_4439;
wire n_520;
wire n_870;
wire n_4985;
wire n_9000;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_8503;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_9139;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_8315;
wire n_1961;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_2844;
wire n_8197;
wire n_402;
wire n_1979;
wire n_6616;
wire n_6719;
wire n_829;
wire n_4814;
wire n_8019;
wire n_8801;
wire n_339;
wire n_6178;
wire n_8707;
wire n_6677;
wire n_2221;
wire n_7875;
wire n_5502;
wire n_8962;
wire n_8931;
wire n_8248;
wire n_1283;
wire n_7550;
wire n_8554;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_2442;
wire n_7238;
wire n_6862;
wire n_8501;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_7292;
wire n_242;
wire n_645;
wire n_7804;
wire n_5098;
wire n_721;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_6443;
wire n_1276;
wire n_8263;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_7248;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_8040;
wire n_5466;
wire n_1528;
wire n_6941;
wire n_7239;
wire n_6552;
wire n_7826;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_8102;
wire n_3999;
wire n_518;
wire n_8196;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_8822;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_7971;
wire n_8885;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_8474;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_1636;
wire n_4597;
wire n_9043;
wire n_8152;
wire n_8269;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_6531;
wire n_3571;
wire n_238;
wire n_4576;
wire n_7577;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_8144;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_7513;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_7812;
wire n_5330;
wire n_6935;
wire n_1560;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_8058;
wire n_8909;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_9242;
wire n_6386;
wire n_3728;
wire n_2722;
wire n_6596;
wire n_612;
wire n_333;
wire n_5107;
wire n_7165;
wire n_512;
wire n_4680;
wire n_5067;
wire n_6830;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_9005;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_6510;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_6781;
wire n_7667;
wire n_4593;
wire n_8024;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_461;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_8107;
wire n_2981;
wire n_225;
wire n_1006;
wire n_546;
wire n_4995;
wire n_1159;
wire n_5873;
wire n_6514;
wire n_4498;
wire n_772;
wire n_6741;
wire n_1245;
wire n_6434;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_3429;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_6593;
wire n_676;
wire n_7827;
wire n_3758;
wire n_7631;
wire n_8748;
wire n_8452;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_8742;
wire n_3777;
wire n_8393;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_212;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_8122;
wire n_2426;
wire n_652;
wire n_6947;
wire n_8403;
wire n_8912;
wire n_4850;
wire n_9154;
wire n_1260;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_798;
wire n_8740;
wire n_5574;
wire n_8310;
wire n_3391;
wire n_5877;
wire n_912;
wire n_6375;
wire n_460;
wire n_7781;
wire n_4786;
wire n_6042;
wire n_8238;
wire n_5203;
wire n_7908;
wire n_8296;
wire n_7091;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_3159;
wire n_6315;
wire n_7855;
wire n_8850;
wire n_2855;
wire n_794;
wire n_2848;
wire n_7886;
wire n_7675;
wire n_6775;
wire n_8943;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_8993;
wire n_9205;
wire n_288;
wire n_1292;
wire n_7774;
wire n_8634;
wire n_8831;
wire n_6970;
wire n_1026;
wire n_6948;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_8676;
wire n_2202;
wire n_306;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_5408;
wire n_8758;
wire n_5812;
wire n_5540;
wire n_7381;
wire n_5804;
wire n_9007;
wire n_8544;
wire n_3240;
wire n_7999;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_9020;
wire n_9260;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_1079;
wire n_5200;
wire n_9235;
wire n_3393;
wire n_8652;
wire n_9112;
wire n_2836;
wire n_7873;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_5992;
wire n_8646;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_9133;
wire n_5684;
wire n_1399;
wire n_7228;
wire n_5981;
wire n_7784;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_8999;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_7713;
wire n_6623;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_1226;
wire n_2224;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_8031;
wire n_3257;
wire n_5737;
wire n_9125;
wire n_8015;
wire n_8412;
wire n_425;
wire n_3730;
wire n_8439;
wire n_8575;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_8499;
wire n_6390;
wire n_7640;
wire n_2302;
wire n_6799;
wire n_8772;
wire n_3014;
wire n_7912;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_8557;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_397;
wire n_3375;
wire n_2768;
wire n_351;
wire n_155;
wire n_3760;
wire n_5661;
wire n_7641;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_8815;
wire n_7949;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_8679;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_1020;
wire n_7764;
wire n_8446;
wire n_9163;
wire n_172;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_8789;
wire n_8128;
wire n_7520;
wire n_5314;
wire n_7616;
wire n_8359;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_6271;
wire n_7235;
wire n_2511;
wire n_564;
wire n_6572;
wire n_9224;
wire n_3981;
wire n_7271;
wire n_9055;
wire n_2681;
wire n_7222;
wire n_8678;
wire n_1689;
wire n_8605;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_345;
wire n_6930;
wire n_2335;
wire n_5482;
wire n_9145;
wire n_3215;
wire n_8443;
wire n_8525;
wire n_1401;
wire n_3138;
wire n_8312;
wire n_776;
wire n_2860;
wire n_8901;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_130;
wire n_6387;
wire n_466;
wire n_4201;
wire n_346;
wire n_6470;
wire n_7206;
wire n_8869;
wire n_552;
wire n_5287;
wire n_8272;
wire n_4719;
wire n_5651;
wire n_264;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_7383;
wire n_3994;
wire n_4636;
wire n_6826;
wire n_3185;
wire n_4983;
wire n_1217;
wire n_327;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_8870;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_8178;
wire n_5524;
wire n_7854;
wire n_926;
wire n_2296;
wire n_5735;
wire n_7959;
wire n_8234;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_7897;
wire n_186;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_8488;
wire n_2241;
wire n_6865;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_7132;
wire n_1570;
wire n_7533;
wire n_3377;
wire n_6722;
wire n_1518;
wire n_6420;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_855;
wire n_8862;
wire n_2059;
wire n_8184;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_1287;
wire n_1611;
wire n_120;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_6981;
wire n_7776;
wire n_4818;
wire n_8001;
wire n_8695;
wire n_7436;
wire n_8767;
wire n_8571;
wire n_7020;
wire n_8064;
wire n_5935;
wire n_6696;
wire n_4916;
wire n_8472;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_6045;
wire n_529;
wire n_1899;
wire n_5934;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_7978;
wire n_5488;
wire n_9099;
wire n_1105;
wire n_6900;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_8787;
wire n_8131;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_7694;
wire n_8771;
wire n_9245;
wire n_5832;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_983;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_699;
wire n_3542;
wire n_301;
wire n_3263;
wire n_5891;
wire n_8150;
wire n_2523;
wire n_1945;
wire n_9168;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_9074;
wire n_3222;
wire n_325;
wire n_1740;
wire n_5016;
wire n_4616;
wire n_6011;
wire n_7465;
wire n_5470;
wire n_8917;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_729;
wire n_8230;
wire n_6222;
wire n_2218;
wire n_8352;
wire n_1122;
wire n_7760;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_6969;
wire n_390;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_8914;
wire n_8821;
wire n_8465;
wire n_6587;
wire n_6688;
wire n_8360;
wire n_6505;
wire n_5362;
wire n_8209;
wire n_388;
wire n_8986;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_7629;
wire n_6987;
wire n_877;
wire n_3995;
wire n_7567;
wire n_8743;
wire n_8963;
wire n_9191;
wire n_3908;
wire n_6453;
wire n_9114;
wire n_6308;
wire n_1055;
wire n_8396;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_8514;
wire n_8550;
wire n_1089;
wire n_7449;
wire n_8151;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_3216;
wire n_2555;
wire n_3568;
wire n_2708;
wire n_6187;
wire n_735;
wire n_6597;
wire n_4844;
wire n_6220;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_7479;
wire n_7882;
wire n_1649;
wire n_2470;
wire n_7517;
wire n_1297;
wire n_3551;
wire n_417;
wire n_1708;
wire n_5037;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_5189;
wire n_4677;
wire n_8070;
wire n_4525;
wire n_8866;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_7878;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_278;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_842;
wire n_148;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_8797;
wire n_6547;
wire n_7177;
wire n_7902;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_476;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_8054;
wire n_982;
wire n_3791;
wire n_915;
wire n_6478;
wire n_2008;
wire n_454;
wire n_298;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_8841;
wire n_9084;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_6906;
wire n_403;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_606;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_7818;
wire n_509;
wire n_7645;
wire n_5385;
wire n_7482;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_8618;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_8538;
wire n_3582;
wire n_8590;
wire n_7907;
wire n_9204;
wire n_8970;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_3459;
wire n_2576;
wire n_8791;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_521;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_7862;
wire n_9130;
wire n_3735;
wire n_8703;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_1513;
wire n_1527;
wire n_3656;
wire n_7721;
wire n_4524;
wire n_9209;
wire n_8061;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_8754;
wire n_8864;
wire n_5941;
wire n_4891;
wire n_8837;
wire n_2629;
wire n_3369;
wire n_8915;
wire n_1257;
wire n_1954;
wire n_8784;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_9086;
wire n_1897;
wire n_8768;
wire n_6999;
wire n_8086;
wire n_8072;
wire n_9014;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_7539;
wire n_9010;
wire n_6440;
wire n_4977;
wire n_8774;
wire n_2492;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_3425;
wire n_2939;
wire n_4876;
wire n_241;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_9044;
wire n_2912;
wire n_5936;
wire n_8307;
wire n_595;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_1757;
wire n_8470;
wire n_1950;
wire n_2264;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_7830;
wire n_8050;
wire n_3124;
wire n_3811;
wire n_295;
wire n_4200;
wire n_190;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_463;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_469;
wire n_9261;
wire n_726;
wire n_5504;
wire n_878;
wire n_7348;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_8010;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_6464;
wire n_8802;
wire n_8950;
wire n_5129;
wire n_806;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_8603;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_1616;
wire n_7935;
wire n_2416;
wire n_8143;
wire n_2064;
wire n_3640;
wire n_9271;
wire n_5663;
wire n_5161;
wire n_7933;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_349;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_6850;
wire n_1505;
wire n_2408;
wire n_7743;
wire n_5389;
wire n_4764;
wire n_4990;
wire n_2986;
wire n_8584;
wire n_949;
wire n_2454;
wire n_9101;
wire n_6550;
wire n_6656;
wire n_8153;
wire n_6972;
wire n_3591;
wire n_8574;
wire n_198;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_7043;
wire n_7986;
wire n_3317;
wire n_8049;
wire n_7266;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_554;
wire n_4420;
wire n_7996;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_354;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_8509;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_594;
wire n_7035;
wire n_4173;
wire n_8354;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_422;
wire n_1269;
wire n_8277;
wire n_7442;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_8583;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_8681;
wire n_6258;
wire n_1288;
wire n_8644;
wire n_7939;
wire n_7715;
wire n_2173;
wire n_3982;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_8609;
wire n_1143;
wire n_9144;
wire n_3973;
wire n_8052;
wire n_4799;
wire n_8733;
wire n_8082;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_7699;
wire n_1153;
wire n_9273;
wire n_271;
wire n_465;
wire n_9196;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_9029;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_562;
wire n_2020;
wire n_7580;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_510;
wire n_5911;
wire n_7340;
wire n_8080;
wire n_256;
wire n_3600;
wire n_7303;
wire n_1023;
wire n_8819;
wire n_914;
wire n_7870;
wire n_689;
wire n_7568;
wire n_6139;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_8487;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3395;
wire n_3011;
wire n_2820;
wire n_497;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_455;
wire n_588;
wire n_638;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_8382;
wire n_1417;
wire n_3096;
wire n_8517;
wire n_7207;
wire n_8827;
wire n_9075;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_8906;
wire n_1603;
wire n_5841;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_8203;
wire n_413;
wire n_2935;
wire n_4246;
wire n_715;
wire n_7618;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_8340;
wire n_4754;
wire n_1534;
wire n_8268;
wire n_8171;
wire n_1290;
wire n_4375;
wire n_617;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_8008;
wire n_7633;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_8553;
wire n_2592;
wire n_8824;
wire n_3490;
wire n_7280;
wire n_8369;
wire n_962;
wire n_5043;
wire n_7339;
wire n_7597;
wire n_8884;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_9225;
wire n_4183;
wire n_7768;
wire n_918;
wire n_1968;
wire n_5645;
wire n_639;
wire n_6455;
wire n_673;
wire n_5020;
wire n_2842;
wire n_7615;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_8271;
wire n_9091;
wire n_3720;
wire n_6183;
wire n_8392;
wire n_8309;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_8874;
wire n_8228;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_8483;
wire n_6003;
wire n_5443;
wire n_8133;
wire n_7612;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_8172;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_5631;
wire n_3481;
wire n_280;
wire n_6994;
wire n_7401;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_9252;
wire n_6185;
wire n_8344;
wire n_692;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_223;
wire n_2150;
wire n_8738;
wire n_8936;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_8226;
wire n_6695;
wire n_7529;
wire n_3354;
wire n_6501;
wire n_5608;
wire n_2204;
wire n_9148;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_6467;
wire n_2231;
wire n_4212;
wire n_622;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_8088;
wire n_5702;
wire n_8930;
wire n_9155;
wire n_8662;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_9046;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_8783;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_8663;
wire n_5277;
wire n_792;
wire n_1262;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_6213;
wire n_1579;
wire n_8364;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_8490;
wire n_8981;
wire n_229;
wire n_9129;
wire n_923;
wire n_1124;
wire n_7872;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_7958;
wire n_2282;
wire n_4605;
wire n_8118;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_8671;
wire n_7101;
wire n_8785;
wire n_1204;
wire n_7843;
wire n_994;
wire n_2428;
wire n_9047;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_7578;
wire n_3410;
wire n_5415;
wire n_856;
wire n_7261;
wire n_8982;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_6993;
wire n_508;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_8100;
wire n_1858;
wire n_353;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_8522;
wire n_1361;
wire n_8381;
wire n_8835;
wire n_6767;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6558;
wire n_6755;
wire n_9108;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_7263;
wire n_3782;
wire n_1317;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_7688;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7925;
wire n_7310;
wire n_294;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_7585;
wire n_8356;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_7772;
wire n_8736;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_8918;
wire n_2402;
wire n_1458;
wire n_679;
wire n_220;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_9022;
wire n_7514;
wire n_1550;
wire n_1358;
wire n_8616;
wire n_1200;
wire n_6105;
wire n_387;
wire n_826;
wire n_5512;
wire n_7738;
wire n_2808;
wire n_2344;
wire n_8838;
wire n_8908;
wire n_3520;
wire n_2392;
wire n_7609;
wire n_9161;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_8607;
wire n_607;
wire n_8213;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_8436;
wire n_7282;
wire n_372;
wire n_8551;
wire n_2770;
wire n_4550;
wire n_9238;
wire n_4347;
wire n_7921;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_9248;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_7489;
wire n_9056;
wire n_6331;
wire n_5308;
wire n_9106;
wire n_311;
wire n_4434;
wire n_5068;
wire n_7863;
wire n_6493;
wire n_7363;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_7968;
wire n_6023;
wire n_7820;
wire n_8437;
wire n_269;
wire n_816;
wire n_7833;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_7750;
wire n_5057;
wire n_446;
wire n_9071;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_7588;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_7697;
wire n_5887;
wire n_7808;
wire n_3068;
wire n_1629;
wire n_9027;
wire n_7603;
wire n_1094;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_8704;
wire n_3002;
wire n_8984;
wire n_7192;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_8613;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_8012;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_8881;
wire n_5531;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_7988;
wire n_550;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_8763;
wire n_6450;
wire n_1152;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_671;
wire n_8387;
wire n_8105;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_7943;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_7377;
wire n_8900;
wire n_4392;
wire n_3103;
wire n_488;
wire n_6064;
wire n_8353;
wire n_505;
wire n_9051;
wire n_2048;
wire n_7723;
wire n_498;
wire n_3028;
wire n_4691;
wire n_7904;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_684;
wire n_5461;
wire n_9098;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_8323;
wire n_6164;
wire n_8711;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_8731;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_8597;
wire n_2515;
wire n_6330;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_838;
wire n_1941;
wire n_7045;
wire n_175;
wire n_3637;
wire n_8534;
wire n_1017;
wire n_8655;
wire n_9210;
wire n_734;
wire n_4893;
wire n_2240;
wire n_7777;
wire n_8302;
wire n_4258;
wire n_5756;
wire n_310;
wire n_8496;
wire n_7693;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_8078;
wire n_2097;
wire n_662;
wire n_3461;
wire n_7682;
wire n_7300;
wire n_939;
wire n_1410;
wire n_2297;
wire n_6861;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_7558;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_572;
wire n_9166;
wire n_8103;
wire n_8719;
wire n_1983;
wire n_7798;
wire n_8879;
wire n_4767;
wire n_8969;
wire n_9141;
wire n_4569;
wire n_948;
wire n_448;
wire n_6528;
wire n_8896;
wire n_3820;
wire n_5144;
wire n_6895;
wire n_3072;
wire n_8335;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_6472;
wire n_3763;
wire n_933;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_492;
wire n_252;
wire n_5183;
wire n_2585;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_8462;
wire n_3228;
wire n_8834;
wire n_8286;
wire n_8417;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_8964;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_7672;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_389;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_8247;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_8639;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_9160;
wire n_5751;
wire n_626;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_7712;
wire n_6885;
wire n_7681;
wire n_5039;
wire n_1818;
wire n_6613;
wire n_6580;
wire n_8566;
wire n_8727;
wire n_4265;
wire n_8482;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_7491;
wire n_265;
wire n_1583;
wire n_8599;
wire n_4612;
wire n_5997;
wire n_8781;
wire n_5375;
wire n_5438;
wire n_9167;
wire n_7150;
wire n_7954;
wire n_7974;
wire n_1264;
wire n_6530;
wire n_6602;
wire n_7915;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_6135;
wire n_246;
wire n_8839;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_8365;
wire n_1102;
wire n_2239;
wire n_6942;
wire n_7860;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_7357;
wire n_8112;
wire n_8489;
wire n_8859;
wire n_8060;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_8244;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_8096;
wire n_7336;
wire n_5932;
wire n_289;
wire n_6598;
wire n_6795;
wire n_6121;
wire n_457;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_8346;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_2152;
wire n_8367;
wire n_2517;
wire n_4696;
wire n_4967;
wire n_9113;
wire n_3484;
wire n_6001;
wire n_411;
wire n_4971;
wire n_2095;
wire n_7493;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_3041;
wire n_357;
wire n_2797;
wire n_412;
wire n_5823;
wire n_8658;
wire n_8898;
wire n_1421;
wire n_2423;
wire n_2208;
wire n_5944;
wire n_5422;
wire n_8905;
wire n_9222;
wire n_6989;
wire n_8237;
wire n_8145;
wire n_6299;
wire n_7424;
wire n_5246;
wire n_8562;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_573;
wire n_2823;
wire n_7273;
wire n_7901;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_7149;
wire n_589;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_8211;
wire n_3268;
wire n_2559;
wire n_8537;
wire n_8946;
wire n_5616;
wire n_1383;
wire n_603;
wire n_8055;
wire n_373;
wire n_4259;
wire n_5870;
wire n_7909;
wire n_2030;
wire n_6053;
wire n_850;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_245;
wire n_319;
wire n_6758;
wire n_2407;
wire n_690;
wire n_5367;
wire n_9069;
wire n_525;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_8332;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_7601;
wire n_8998;
wire n_1837;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_189;
wire n_8157;
wire n_2006;
wire n_4953;
wire n_8484;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_7596;
wire n_5294;
wire n_8161;
wire n_5570;
wire n_6411;
wire n_2731;
wire n_3703;
wire n_5670;
wire n_5411;
wire n_1246;
wire n_9211;
wire n_5265;
wire n_5955;
wire n_7549;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_8692;
wire n_3435;
wire n_410;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_9243;
wire n_6918;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_8812;
wire n_568;
wire n_8682;
wire n_4796;
wire n_8290;
wire n_1088;
wire n_7138;
wire n_766;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_7976;
wire n_377;
wire n_2750;
wire n_8890;
wire n_2547;
wire n_8747;
wire n_7617;
wire n_279;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_8062;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_7700;
wire n_8275;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_8667;
wire n_3220;
wire n_4581;
wire n_9192;
wire n_6008;
wire n_500;
wire n_665;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_9134;
wire n_3679;
wire n_738;
wire n_5575;
wire n_6654;
wire n_7661;
wire n_672;
wire n_4968;
wire n_7801;
wire n_8807;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_7876;
wire n_2735;
wire n_953;
wire n_4214;
wire n_143;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_557;
wire n_3419;
wire n_7323;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_6517;
wire n_795;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_9127;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_8048;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_7929;
wire n_486;
wire n_2782;
wire n_569;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_8212;
wire n_4950;
wire n_1650;
wire n_7755;
wire n_6504;
wire n_4176;
wire n_9078;
wire n_7556;
wire n_222;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_7216;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_8043;
wire n_8223;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_8159;
wire n_5845;
wire n_8868;
wire n_4608;
wire n_6691;
wire n_432;
wire n_293;
wire n_3948;
wire n_4839;
wire n_9174;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_9132;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_206;
wire n_2332;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_611;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_136;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_300;
wire n_6025;
wire n_3049;
wire n_8434;
wire n_3634;
wire n_5436;
wire n_7962;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_8608;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_376;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_8656;
wire n_3861;
wire n_5096;
wire n_9183;
wire n_2043;
wire n_6771;
wire n_7905;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_9117;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_7476;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_8249;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_9062;
wire n_209;
wire n_5240;
wire n_5718;
wire n_1461;
wire n_7208;
wire n_5503;
wire n_7718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_6567;
wire n_503;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_9001;
wire n_7290;
wire n_6868;
wire n_5131;
wire n_9081;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_9156;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_8717;
wire n_5174;
wire n_9024;
wire n_9198;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_380;
wire n_3119;
wire n_6671;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_7632;
wire n_4394;
wire n_257;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_8842;
wire n_475;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_8073;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_577;
wire n_5610;
wire n_407;
wire n_8576;
wire n_916;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_1555;
wire n_8799;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_7265;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_8181;
wire n_5808;
wire n_1182;
wire n_6527;
wire n_4594;
wire n_8447;
wire n_8045;
wire n_7289;
wire n_7538;
wire n_2748;
wire n_4642;
wire n_6913;
wire n_1376;
wire n_7473;
wire n_7242;
wire n_9253;
wire n_6533;
wire n_513;
wire n_179;
wire n_7164;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_8022;
wire n_3544;
wire n_6845;
wire n_5300;
wire n_8227;
wire n_7853;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_436;
wire n_5770;
wire n_7483;
wire n_8756;
wire n_5710;
wire n_324;
wire n_1491;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_1083;
wire n_274;
wire n_5333;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_8604;
wire n_8809;
wire n_8976;
wire n_3510;
wire n_7046;
wire n_7834;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_8940;
wire n_5008;
wire n_1312;
wire n_9077;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_563;
wire n_2219;
wire n_8844;
wire n_6148;
wire n_8995;
wire n_2100;
wire n_8255;
wire n_3666;
wire n_5538;
wire n_990;
wire n_6357;
wire n_867;
wire n_8216;
wire n_8693;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_9123;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_7811;
wire n_8669;
wire n_4285;
wire n_7097;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_9177;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_7880;
wire n_712;
wire n_8769;
wire n_909;
wire n_6713;
wire n_8149;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_7851;
wire n_2220;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_6108;
wire n_7664;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_7332;
wire n_8990;
wire n_5862;
wire n_471;
wire n_7477;
wire n_1914;
wire n_8208;
wire n_2253;
wire n_7468;
wire n_5886;
wire n_7714;
wire n_7899;
wire n_8710;
wire n_6415;
wire n_8479;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_8512;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_9087;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_7845;
wire n_347;
wire n_2434;
wire n_183;
wire n_1234;
wire n_3936;
wire n_479;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_9079;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_7858;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_6392;
wire n_6513;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_9197;
wire n_1237;
wire n_6720;
wire n_5883;
wire n_9140;
wire n_8401;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_370;
wire n_7680;
wire n_5630;
wire n_6666;
wire n_286;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_6815;
wire n_9203;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_8450;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_7710;
wire n_8788;
wire n_5394;
wire n_8324;
wire n_5975;
wire n_4242;
wire n_4751;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_9057;
wire n_3300;
wire n_7061;
wire n_8104;
wire n_7066;
wire n_9068;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_8014;
wire n_4122;
wire n_6661;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_8623;
wire n_4952;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_8651;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_9257;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_7783;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_9049;
wire n_487;
wire n_4728;
wire n_7171;
wire n_7990;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_7003;
wire n_8137;
wire n_2187;
wire n_1413;
wire n_8413;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_158;
wire n_3882;
wire n_3916;
wire n_6922;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_405;
wire n_3332;
wire n_8300;
wire n_8069;
wire n_7501;
wire n_320;
wire n_6432;
wire n_7984;
wire n_2055;
wire n_2998;
wire n_7366;
wire n_1423;
wire n_8173;
wire n_4359;
wire n_481;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_7589;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_218;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_1798;
wire n_8091;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_6699;
wire n_547;
wire n_439;
wire n_677;
wire n_3983;
wire n_9067;
wire n_8254;
wire n_703;
wire n_8400;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_7511;
wire n_326;
wire n_227;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_9033;
wire n_6957;
wire n_5074;
wire n_7917;
wire n_3788;
wire n_3939;
wire n_590;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_8368;
wire n_6694;
wire n_545;
wire n_9247;
wire n_2496;
wire n_3260;
wire n_8463;
wire n_536;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_1602;
wire n_7422;
wire n_3139;
wire n_8889;
wire n_427;
wire n_3801;
wire n_5681;
wire n_9244;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_9195;
wire n_8322;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_8987;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_7621;
wire n_8274;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_163;
wire n_2716;
wire n_6441;
wire n_7158;
wire n_7572;
wire n_314;
wire n_2944;
wire n_3439;
wire n_2780;
wire n_1120;
wire n_7500;
wire n_1202;
wire n_4084;
wire n_627;
wire n_7985;
wire n_1371;
wire n_4240;
wire n_8657;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_233;
wire n_8954;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_8311;
wire n_5748;
wire n_4393;
wire n_321;
wire n_6662;
wire n_7494;
wire n_9088;
wire n_3984;
wire n_1586;
wire n_8728;
wire n_1431;
wire n_8994;
wire n_4389;
wire n_6433;
wire n_1763;
wire n_8398;
wire n_6200;
wire n_5641;
wire n_8407;
wire n_8071;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_8528;
wire n_9227;
wire n_5657;
wire n_8475;
wire n_297;
wire n_2379;
wire n_3579;
wire n_9072;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_9054;
wire n_4551;
wire n_178;
wire n_551;
wire n_4521;
wire n_6956;
wire n_7587;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_7704;
wire n_5420;
wire n_6497;
wire n_8511;
wire n_7865;
wire n_2283;
wire n_5206;
wire n_582;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_534;
wire n_2508;
wire n_3186;
wire n_6701;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_8867;
wire n_3417;
wire n_8246;
wire n_560;
wire n_8558;
wire n_890;
wire n_3626;
wire n_451;
wire n_4598;
wire n_4464;
wire n_8925;
wire n_5106;
wire n_7881;
wire n_9147;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_8641;
wire n_2493;
wire n_5080;
wire n_535;
wire n_4565;
wire n_7032;
wire n_3392;
wire n_1800;
wire n_7198;
wire n_6884;
wire n_7752;
wire n_5081;
wire n_8201;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_7953;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_8046;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_8414;
wire n_3024;
wire n_8292;
wire n_5567;
wire n_9138;
wire n_5406;
wire n_8647;
wire n_6362;
wire n_9213;
wire n_4328;
wire n_8543;
wire n_1854;
wire n_666;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_8331;
wire n_999;
wire n_2280;
wire n_8317;
wire n_7126;
wire n_5867;
wire n_456;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_7496;
wire n_6430;
wire n_9179;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_342;
wire n_5602;
wire n_2035;
wire n_7196;
wire n_4928;
wire n_2614;
wire n_7360;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_6678;
wire n_7982;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_8174;
wire n_8187;
wire n_8929;
wire n_4436;
wire n_5822;
wire n_5786;
wire n_3586;
wire n_8846;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_6385;
wire n_1668;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_8032;
wire n_5417;
wire n_4545;
wire n_8200;
wire n_4758;
wire n_1161;
wire n_8036;
wire n_5713;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_9190;
wire n_8586;
wire n_8524;
wire n_618;
wire n_1191;
wire n_4535;
wire n_7518;
wire n_8828;
wire n_4385;
wire n_7779;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_7575;
wire n_2337;
wire n_7073;
wire n_8092;
wire n_1786;
wire n_6309;
wire n_8370;
wire n_3732;
wire n_9109;
wire n_211;
wire n_1804;
wire n_408;
wire n_8135;
wire n_6519;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_592;
wire n_4558;
wire n_1318;
wire n_8764;
wire n_1632;
wire n_1769;
wire n_7349;
wire n_1929;
wire n_8502;
wire n_4319;
wire n_6585;
wire n_7786;
wire n_9021;
wire n_8454;
wire n_2929;
wire n_4358;
wire n_9122;
wire n_1526;
wire n_7579;
wire n_7122;
wire n_4874;
wire n_180;
wire n_2656;
wire n_4904;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_640;
wire n_1733;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_7624;
wire n_1807;
wire n_1123;
wire n_8776;
wire n_2857;
wire n_8564;
wire n_8343;
wire n_7828;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_8718;
wire n_752;
wire n_985;
wire n_5506;
wire n_7543;
wire n_5475;
wire n_8042;
wire n_7727;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_9013;
wire n_5431;
wire n_8379;
wire n_643;
wire n_8034;
wire n_226;
wire n_7778;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_7019;
wire n_682;
wire n_9126;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_8441;
wire n_1429;
wire n_2353;
wire n_7702;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_686;
wire n_1154;
wire n_584;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_6685;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_8569;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_8592;
wire n_8865;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_7952;
wire n_7347;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_7791;
wire n_6971;
wire n_8362;
wire n_3336;
wire n_8632;
wire n_7739;
wire n_396;
wire n_7945;
wire n_9045;
wire n_8361;
wire n_7656;
wire n_5903;
wire n_7199;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_9159;
wire n_8561;
wire n_6549;
wire n_725;
wire n_8611;
wire n_8410;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_6683;
wire n_3067;
wire n_154;
wire n_3809;
wire n_4921;
wire n_473;
wire n_1852;
wire n_801;
wire n_5912;
wire n_5745;
wire n_7923;
wire n_6086;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_8878;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_272;
wire n_8492;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_8888;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_7610;
wire n_7107;
wire n_4561;
wire n_1541;
wire n_597;
wire n_3291;
wire n_7456;
wire n_8095;
wire n_7369;
wire n_1472;
wire n_1050;
wire n_7548;
wire n_2578;
wire n_152;
wire n_1201;
wire n_8735;
wire n_7598;
wire n_1185;
wire n_2475;
wire n_7250;
wire n_8808;
wire n_9201;
wire n_8902;
wire n_7823;
wire n_8833;
wire n_4715;
wire n_6157;
wire n_8796;
wire n_2715;
wire n_335;
wire n_2665;
wire n_4879;
wire n_344;
wire n_8794;
wire n_5044;
wire n_210;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_9274;
wire n_8549;
wire n_6676;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_224;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_7525;
wire n_4418;
wire n_7924;
wire n_3341;
wire n_9232;
wire n_8690;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_8593;
wire n_276;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4412;
wire n_4151;
wire n_2036;
wire n_6923;
wire n_7649;
wire n_843;
wire n_8195;
wire n_8009;
wire n_8588;
wire n_3358;
wire n_6704;
wire n_7634;
wire n_9090;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_7406;
wire n_4682;
wire n_1128;
wire n_6673;
wire n_2419;
wire n_2330;
wire n_6534;
wire n_8805;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_1440;
wire n_6246;
wire n_1370;
wire n_305;
wire n_5005;
wire n_6126;
wire n_7372;
wire n_8596;
wire n_1549;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_7844;
wire n_5207;
wire n_7934;
wire n_361;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_7009;
wire n_5474;
wire n_3376;
wire n_181;
wire n_9121;
wire n_7371;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_683;
wire n_7463;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_9158;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_660;
wire n_464;
wire n_4413;
wire n_8627;
wire n_1210;
wire n_3307;
wire n_8945;
wire n_9142;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_9216;
wire n_9189;
wire n_6723;
wire n_7398;
wire n_1038;
wire n_3723;
wire n_7941;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_8858;
wire n_414;
wire n_571;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_8916;
wire n_613;
wire n_1022;
wire n_5465;
wire n_171;
wire n_8745;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_8169;
wire n_6184;
wire n_8018;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_7083;
wire n_316;
wire n_125;
wire n_1973;
wire n_1444;
wire n_820;
wire n_8260;
wire n_254;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_7701;
wire n_8688;
wire n_7969;
wire n_8279;
wire n_4384;
wire n_8793;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_6312;
wire n_7683;
wire n_532;
wire n_2154;
wire n_7669;
wire n_1986;
wire n_8298;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_8023;
wire n_7330;
wire n_6007;
wire n_621;
wire n_6734;
wire n_6535;
wire n_8053;
wire n_8059;
wire n_1772;
wire n_6879;
wire n_493;
wire n_1311;
wire n_3106;
wire n_7190;
wire n_6208;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_7692;
wire n_697;
wire n_4620;
wire n_6255;
wire n_6457;
wire n_5397;
wire n_9272;
wire n_4924;
wire n_4044;
wire n_8372;
wire n_6270;
wire n_2305;
wire n_8737;
wire n_5996;
wire n_880;
wire n_5566;
wire n_3304;
wire n_7288;
wire n_4388;
wire n_7362;
wire n_7082;
wire n_7237;
wire n_8988;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_739;
wire n_1028;
wire n_530;
wire n_8723;
wire n_9050;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_7042;
wire n_8419;
wire n_2809;
wire n_5652;
wire n_8893;
wire n_975;
wire n_1645;
wire n_5805;
wire n_7304;
wire n_932;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_8077;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_7754;
wire n_8826;
wire n_3178;
wire n_268;
wire n_7023;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_8959;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_7981;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_191;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_8712;
wire n_1011;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_8109;
wire n_116;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_7378;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_7877;
wire n_7787;
wire n_7836;
wire n_8515;
wire n_8725;
wire n_8007;
wire n_2387;
wire n_4318;
wire n_332;
wire n_8910;
wire n_5227;
wire n_830;
wire n_5902;
wire n_987;
wire n_2510;
wire n_9164;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_8301;
wire n_6764;
wire n_7871;
wire n_541;
wire n_499;
wire n_2639;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_8892;
wire n_5386;
wire n_1167;
wire n_6215;
wire n_4554;
wire n_7571;
wire n_8252;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_6955;
wire n_7563;
wire n_5952;
wire n_7180;
wire n_2086;
wire n_1926;
wire n_8972;
wire n_8494;
wire n_6569;
wire n_1630;
wire n_7919;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_8278;
wire n_443;
wire n_3431;
wire n_8180;
wire n_3355;
wire n_7031;
wire n_1738;
wire n_5716;
wire n_8941;
wire n_8891;
wire n_406;
wire n_3897;
wire n_7103;
wire n_139;
wire n_6605;
wire n_1735;
wire n_391;
wire n_5888;
wire n_9266;
wire n_4005;
wire n_8270;
wire n_8231;
wire n_4181;
wire n_2543;
wire n_2597;
wire n_1077;
wire n_2321;
wire n_6832;
wire n_5980;
wire n_8683;
wire n_956;
wire n_765;
wire n_4092;
wire n_122;
wire n_4875;
wire n_7771;
wire n_8903;
wire n_4255;
wire n_2758;
wire n_385;
wire n_6544;
wire n_8810;
wire n_6469;
wire n_5036;
wire n_1271;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_399;
wire n_7130;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_8932;
wire n_8264;
wire n_2471;
wire n_7134;
wire n_3042;
wire n_8288;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_1551;
wire n_5271;
wire n_4849;
wire n_2039;
wire n_7133;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_3838;
wire n_6651;
wire n_6289;
wire n_9255;
wire n_8882;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_8388;
wire n_5445;
wire n_2734;
wire n_8067;
wire n_8385;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_8670;
wire n_4504;
wire n_3598;
wire n_7706;
wire n_7813;
wire n_4917;
wire n_8142;
wire n_2420;
wire n_7992;
wire n_9085;
wire n_7643;
wire n_153;
wire n_648;
wire n_6836;
wire n_3273;
wire n_9120;
wire n_2918;
wire n_6595;
wire n_835;
wire n_9136;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_401;
wire n_7628;
wire n_1792;
wire n_5628;
wire n_504;
wire n_5245;
wire n_2062;
wire n_483;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_8224;
wire n_5472;
wire n_6035;
wire n_9042;
wire n_839;
wire n_1754;
wire n_7236;
wire n_9239;
wire n_4833;
wire n_3394;
wire n_6405;
wire n_8345;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_8614;
wire n_8242;
wire n_6786;
wire n_4564;
wire n_8299;
wire n_1848;
wire n_9131;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_9060;
wire n_3581;
wire n_8110;
wire n_5072;
wire n_8529;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_8951;
wire n_2260;
wire n_323;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_8700;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_7519;
wire n_7802;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_7457;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_6416;
wire n_654;
wire n_2933;
wire n_8468;
wire n_9031;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_8933;
wire n_6214;
wire n_3952;
wire n_8636;
wire n_9006;
wire n_9221;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_7049;
wire n_7884;
wire n_6945;
wire n_8378;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_7749;
wire n_7592;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_539;
wire n_8283;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_7914;
wire n_1866;
wire n_8860;
wire n_2664;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_4390;
wire n_459;
wire n_1782;
wire n_7892;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4609;
wire n_4361;
wire n_7325;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_723;
wire n_1393;
wire n_7674;
wire n_8686;
wire n_6175;
wire n_6445;
wire n_8563;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_8493;
wire n_6198;
wire n_5172;
wire n_881;
wire n_1019;
wire n_1477;
wire n_6499;
wire n_1982;
wire n_7983;
wire n_641;
wire n_5311;
wire n_8765;
wire n_910;
wire n_290;
wire n_5164;
wire n_4964;
wire n_9153;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_217;
wire n_7361;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_201;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_8653;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_8601;
wire n_1043;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_255;
wire n_2869;
wire n_8333;
wire n_9097;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_1613;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_196;
wire n_3244;
wire n_1779;
wire n_3112;
wire n_954;
wire n_2562;
wire n_2051;
wire n_3196;
wire n_231;
wire n_8708;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_664;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_8659;
wire n_6732;
wire n_8759;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_544;
wire n_7646;
wire n_3779;
wire n_599;
wire n_6982;
wire n_537;
wire n_1063;
wire n_7291;
wire n_8790;
wire n_991;
wire n_2275;
wire n_7668;
wire n_7435;
wire n_4606;
wire n_8832;
wire n_8305;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_8453;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_583;
wire n_1000;
wire n_313;
wire n_4868;
wire n_7017;
wire n_378;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_4465;
wire n_8127;
wire n_2596;
wire n_5217;
wire n_8337;
wire n_9115;
wire n_3986;
wire n_7861;
wire n_3725;
wire n_5558;
wire n_472;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_7889;
wire n_208;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_4852;
wire n_275;
wire n_7554;
wire n_3202;
wire n_8508;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_7648;
wire n_8968;
wire n_147;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_7653;
wire n_6400;
wire n_1644;
wire n_7846;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_8347;
wire n_131;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_250;
wire n_773;
wire n_5135;
wire n_7551;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_718;
wire n_1434;
wire n_8093;
wire n_8899;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_7737;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_523;
wire n_1662;
wire n_8481;
wire n_3249;
wire n_3483;
wire n_6851;
wire n_6621;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_7606;
wire n_7420;
wire n_8115;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_484;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_1574;
wire n_3033;
wire n_893;
wire n_9182;
wire n_1582;
wire n_8182;
wire n_1981;
wire n_2824;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_796;
wire n_127;
wire n_531;
wire n_1374;
wire n_2089;
wire n_7896;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_5900;
wire n_8629;
wire n_8186;
wire n_7319;
wire n_1486;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_9246;
wire n_4342;
wire n_691;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_8233;
wire n_4382;
wire n_4085;
wire n_423;
wire n_2509;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_8282;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_5851;
wire n_7516;
wire n_6928;
wire n_6317;
wire n_6707;
wire n_7244;
wire n_187;
wire n_1463;
wire n_4626;
wire n_7625;
wire n_8750;
wire n_4997;
wire n_8183;
wire n_5065;
wire n_9104;
wire n_6806;
wire n_924;
wire n_7991;
wire n_781;
wire n_8637;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_8792;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_7857;
wire n_7970;
wire n_1706;
wire n_2461;
wire n_8258;
wire n_3719;
wire n_117;
wire n_7154;
wire n_524;
wire n_1214;
wire n_634;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_8390;
wire n_8416;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_8696;
wire n_9185;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_7175;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_7163;
wire n_3797;
wire n_1836;
wire n_7027;
wire n_3416;
wire n_8552;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_7964;
wire n_5749;
wire n_6320;
wire n_6316;
wire n_8619;
wire n_419;
wire n_7068;
wire n_2908;
wire n_8594;
wire n_270;
wire n_4106;
wire n_285;
wire n_2156;
wire n_1184;
wire n_202;
wire n_8162;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_7327;
wire n_1277;
wire n_1746;
wire n_6610;
wire n_1062;
wire n_5998;
wire n_8318;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_167;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_8425;
wire n_6752;
wire n_6959;
wire n_6250;
wire n_3283;
wire n_259;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_7864;
wire n_3451;
wire n_8051;
wire n_4734;
wire n_6675;
wire n_7955;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_9039;
wire n_7384;
wire n_267;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_5678;
wire n_6561;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_7512;
wire n_1718;
wire n_7814;
wire n_8389;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_200;
wire n_2539;
wire n_8620;
wire n_5555;
wire n_2078;
wire n_8886;
wire n_1145;
wire n_7152;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_8202;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_7223;
wire n_5251;
wire n_1314;
wire n_8755;
wire n_1512;
wire n_8668;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_8979;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_7761;
wire n_8141;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_8199;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_8004;
wire n_8383;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_7437;
wire n_6489;
wire n_9023;
wire n_5310;
wire n_2769;
wire n_8895;
wire n_438;
wire n_8680;
wire n_1548;
wire n_4987;
wire n_6714;
wire n_8394;
wire n_440;
wire n_7849;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_7417;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_2902;
wire n_6245;
wire n_6030;
wire n_4360;
wire n_1544;
wire n_6620;
wire n_6791;
wire n_4540;
wire n_9220;
wire n_6821;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_8198;
wire n_1354;
wire n_8665;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_7859;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_491;
wire n_1595;
wire n_8017;
wire n_1142;
wire n_5477;
wire n_260;
wire n_2727;
wire n_942;
wire n_7523;
wire n_5234;
wire n_1416;
wire n_6890;
wire n_9184;
wire n_7559;
wire n_9037;
wire n_7576;
wire n_6988;
wire n_8303;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_8000;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_7769;
wire n_9193;
wire n_7257;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_8852;
wire n_5007;
wire n_8709;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_9218;
wire n_4357;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_287;
wire n_3191;
wire n_1716;
wire n_302;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_8782;
wire n_7081;
wire n_7742;
wire n_5253;
wire n_3588;
wire n_355;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_9162;
wire n_135;
wire n_3095;
wire n_947;
wire n_7341;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_4775;
wire n_6256;
wire n_482;
wire n_2620;
wire n_1833;
wire n_8716;
wire n_1691;
wire n_8250;
wire n_7264;
wire n_7842;
wire n_2499;
wire n_2549;
wire n_6648;
wire n_7492;
wire n_804;
wire n_6649;
wire n_8714;
wire n_1656;
wire n_8357;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_3885;
wire n_955;
wire n_8466;
wire n_4264;
wire n_5954;
wire n_9015;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_514;
wire n_6431;
wire n_418;
wire n_8589;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_8266;
wire n_3839;
wire n_8587;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_8876;
wire n_9214;
wire n_4206;
wire n_4099;
wire n_2415;
wire n_8922;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_9070;
wire n_8498;
wire n_4794;
wire n_4843;
wire n_669;
wire n_5580;
wire n_5215;
wire n_337;
wire n_437;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_8457;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_8267;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_615;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_517;
wire n_8124;
wire n_3604;
wire n_8545;
wire n_5430;
wire n_6041;
wire n_8526;
wire n_824;
wire n_159;
wire n_8319;
wire n_7997;
wire n_5659;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_144;
wire n_3792;
wire n_7950;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_8581;
wire n_8214;
wire n_7793;
wire n_9053;
wire n_8516;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_470;
wire n_3021;
wire n_8989;
wire n_7746;
wire n_477;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_7570;
wire n_2898;
wire n_1825;
wire n_6912;
wire n_3567;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_9217;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_1731;
wire n_799;
wire n_7894;
wire n_1147;
wire n_7957;
wire n_8262;
wire n_2378;
wire n_5530;
wire n_6718;
wire n_8289;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_7121;
wire n_7531;
wire n_6410;
wire n_356;
wire n_6473;
wire n_8087;
wire n_4056;
wire n_4806;
wire n_7961;
wire n_1674;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4723;
wire n_4484;
wire n_2142;
wire n_8863;
wire n_4517;
wire n_2896;
wire n_8701;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_9237;
wire n_2311;
wire n_6857;
wire n_8705;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_6975;
wire n_7763;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_205;
wire n_7703;
wire n_7928;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_8722;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_713;
wire n_3179;
wire n_598;
wire n_6622;
wire n_7665;
wire n_5522;
wire n_3889;
wire n_7677;
wire n_5262;
wire n_4836;
wire n_3262;
wire n_5319;
wire n_927;
wire n_7469;
wire n_261;
wire n_3699;
wire n_6118;
wire n_706;
wire n_2120;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_1419;
wire n_8622;
wire n_3816;
wire n_8099;
wire n_8729;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_4207;
wire n_8085;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_348;
wire n_9173;
wire n_2312;
wire n_7203;
wire n_8947;
wire n_7797;
wire n_1826;
wire n_9267;
wire n_5943;
wire n_6556;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_7128;
wire n_5335;
wire n_1259;
wire n_6365;
wire n_8459;
wire n_7111;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_8478;
wire n_5284;
wire n_8786;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_8887;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_8851;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_8540;
wire n_8276;
wire n_7284;
wire n_3615;
wire n_5516;
wire n_7057;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_9152;
wire n_8706;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_145;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_8532;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_7278;
wire n_9103;
wire n_9111;
wire n_6772;
wire n_7088;
wire n_7799;
wire n_5698;
wire n_5731;
wire n_8871;
wire n_4007;
wire n_1456;
wire n_8433;
wire n_9065;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_7048;
wire n_7979;
wire n_6617;
wire n_553;
wire n_7725;
wire n_814;
wire n_578;
wire n_5120;
wire n_3572;
wire n_8371;
wire n_2975;
wire n_2399;
wire n_8547;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_8467;
wire n_647;
wire n_2027;
wire n_2932;
wire n_8409;
wire n_6217;
wire n_600;
wire n_3118;
wire n_9157;
wire n_5560;
wire n_9170;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_6777;
wire n_502;
wire n_8640;
wire n_5455;
wire n_6742;
wire n_1467;
wire n_7447;
wire n_5209;
wire n_247;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_8431;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_8415;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_6479;
wire n_5099;
wire n_681;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_7365;
wire n_3443;
wire n_8329;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_5022;
wire n_8089;
wire n_9208;
wire n_6370;
wire n_9223;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_3009;
wire n_8633;
wire n_777;
wire n_7095;
wire n_7390;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_920;
wire n_8541;
wire n_8762;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_1132;
wire n_8125;
wire n_501;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_9226;
wire n_6712;
wire n_7530;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_7471;
wire n_6465;
wire n_221;
wire n_8188;
wire n_5673;
wire n_861;
wire n_8615;
wire n_5814;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_8011;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_8923;
wire n_281;
wire n_3326;
wire n_8624;
wire n_262;
wire n_8222;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_8206;
wire n_6515;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_8065;
wire n_527;
wire n_2949;
wire n_7008;
wire n_6468;
wire n_7709;
wire n_4269;
wire n_1927;
wire n_7540;
wire n_7581;
wire n_343;
wire n_1222;
wire n_7139;
wire n_8935;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_7782;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_8155;
wire n_2449;
wire n_4428;
wire n_745;
wire n_6483;
wire n_1572;
wire n_7770;
wire n_8397;
wire n_8568;
wire n_4463;
wire n_5357;
wire n_8175;
wire n_7173;
wire n_3648;
wire n_9254;
wire n_6810;
wire n_6576;
wire n_1975;
wire n_5421;
wire n_9083;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_8026;
wire n_6667;
wire n_9175;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_8974;
wire n_6305;
wire n_8836;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_8168;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_7751;
wire n_7951;
wire n_657;
wire n_7060;
wire n_3924;
wire n_3997;
wire n_8873;
wire n_7591;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_6750;
wire n_7444;
wire n_7911;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_2306;
wire n_7790;
wire n_2071;
wire n_7426;
wire n_430;
wire n_4400;
wire n_3953;
wire n_7502;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_6855;
wire n_8170;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_5768;
wire n_1342;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_8120;
wire n_9116;
wire n_8825;
wire n_852;
wire n_9169;
wire n_2916;
wire n_7252;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_4192;
wire n_8003;
wire n_9215;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_8395;
wire n_3400;
wire n_5972;
wire n_7065;
wire n_1466;
wire n_8083;
wire n_6177;
wire n_8057;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_9259;
wire n_5146;
wire n_7367;
wire n_8164;
wire n_7405;
wire n_7267;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_8877;
wire n_1329;
wire n_6825;
wire n_7614;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_134;
wire n_4035;
wire n_9150;
wire n_6952;
wire n_1480;
wire n_3670;
wire n_8366;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_8476;
wire n_1605;
wire n_3060;
wire n_6218;
wire n_7685;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_157;
wire n_7619;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_624;
wire n_5577;
wire n_876;
wire n_9100;
wire n_5872;
wire n_7883;
wire n_6692;
wire n_5017;
wire n_8854;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_9262;
wire n_5976;
wire n_4717;
wire n_9249;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_602;
wire n_854;
wire n_8256;
wire n_2091;
wire n_393;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_7270;
wire n_1658;
wire n_1072;
wire n_8621;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_8577;
wire n_9019;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_7731;
wire n_6626;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_7034;
wire n_8654;
wire n_3694;
wire n_6854;
wire n_7940;
wire n_771;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_421;
wire n_3702;
wire n_5930;
wire n_8952;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_7537;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_7458;
wire n_1824;
wire n_7740;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_819;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_3543;
wire n_8421;
wire n_7179;
wire n_1776;
wire n_3448;
wire n_7433;
wire n_4279;
wire n_605;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_6334;
wire n_6257;
wire n_4152;
wire n_6874;
wire n_8911;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_8971;
wire n_7015;
wire n_6355;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_7987;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_9009;
wire n_2368;
wire n_6377;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_7272;
wire n_8215;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_151;
wire n_7906;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_7765;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_8949;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_6511;
wire n_7815;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_8983;
wire n_4969;
wire n_8121;
wire n_5252;
wire n_5777;
wire n_8942;
wire n_7785;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_566;
wire n_7728;
wire n_8280;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_169;
wire n_7181;
wire n_173;
wire n_2796;
wire n_858;
wire n_5393;
wire n_8328;
wire n_4817;
wire n_8861;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_8427;
wire n_2136;
wire n_433;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_253;
wire n_928;
wire n_3769;
wire n_7825;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_128;
wire n_7916;
wire n_3055;
wire n_8194;
wire n_420;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_748;
wire n_7903;
wire n_7089;
wire n_1045;
wire n_8217;
wire n_1881;
wire n_2635;
wire n_7604;
wire n_7647;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_330;
wire n_5868;
wire n_6417;
wire n_328;
wire n_368;
wire n_8285;
wire n_7145;
wire n_8521;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_9178;
wire n_7803;
wire n_2713;
wire n_1422;
wire n_8448;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_5104;
wire n_6961;
wire n_576;
wire n_8732;
wire n_511;
wire n_7622;
wire n_429;
wire n_7839;
wire n_6792;
wire n_7720;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_8136;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_8420;
wire n_141;
wire n_4430;
wire n_8386;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_1356;
wire n_6831;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_312;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_7809;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_623;
wire n_3509;
wire n_8746;
wire n_1403;
wire n_5395;
wire n_453;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_8857;
wire n_543;
wire n_6986;
wire n_3456;
wire n_4532;
wire n_236;
wire n_601;
wire n_7564;
wire n_628;
wire n_5863;
wire n_8185;
wire n_8313;
wire n_6633;
wire n_3790;
wire n_7775;
wire n_907;
wire n_7118;
wire n_9234;
wire n_7960;
wire n_6152;
wire n_5734;
wire n_8281;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_7636;
wire n_4341;
wire n_1694;
wire n_6925;
wire n_7186;
wire n_593;
wire n_8766;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_5480;
wire n_4650;
wire n_6428;
wire n_609;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_8066;
wire n_7666;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_7967;
wire n_5977;
wire n_519;
wire n_8314;
wire n_384;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_9064;
wire n_3409;
wire n_4381;
wire n_8239;
wire n_9092;
wire n_3583;
wire n_4316;
wire n_7301;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_8497;
wire n_1157;
wire n_7262;
wire n_234;
wire n_5959;
wire n_8210;
wire n_8056;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_7584;
wire n_7748;
wire n_1789;
wire n_9066;
wire n_763;
wire n_6301;
wire n_2174;
wire n_540;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_1687;
wire n_4703;
wire n_6282;
wire n_4934;
wire n_7686;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_395;
wire n_6737;
wire n_1587;
wire n_213;
wire n_2340;
wire n_4804;
wire n_8404;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_6459;
wire n_1427;
wire n_7670;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_8505;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_585;
wire n_1617;
wire n_2600;
wire n_8606;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_9059;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_3329;
wire n_3833;
wire n_2927;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_9002;
wire n_3402;
wire n_1621;
wire n_6448;
wire n_9229;
wire n_5186;
wire n_7930;
wire n_7487;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_580;
wire n_3664;
wire n_4218;
wire n_434;
wire n_4687;
wire n_7077;
wire n_394;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_8518;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_5604;
wire n_3470;
wire n_243;
wire n_7663;
wire n_8350;
wire n_8741;
wire n_5221;
wire n_7024;
wire n_1407;
wire n_8148;
wire n_8408;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_8236;
wire n_7214;
wire n_8806;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_8295;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_7977;
wire n_121;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_8167;
wire n_8377;
wire n_3989;
wire n_7652;
wire n_4644;
wire n_8956;
wire n_4752;
wire n_8673;
wire n_4746;
wire n_7566;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_8760;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_322;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_558;
wire n_5325;
wire n_4231;
wire n_8960;
wire n_8957;
wire n_9008;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_653;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_8207;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_556;
wire n_170;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_1471;
wire n_6212;
wire n_3440;
wire n_9194;
wire n_6816;
wire n_8904;
wire n_3658;
wire n_7374;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_7678;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_7975;
wire n_8451;
wire n_6089;
wire n_591;
wire n_5634;
wire n_5133;
wire n_7553;
wire n_8527;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_1625;
wire n_7086;
wire n_5689;
wire n_7732;
wire n_7891;
wire n_9089;
wire n_4578;
wire n_318;
wire n_8840;
wire n_5644;
wire n_9137;
wire n_3644;
wire n_8038;
wire n_8190;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_528;
wire n_9080;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_9151;
wire n_8179;
wire n_7038;
wire n_7994;
wire n_4470;
wire n_4187;
wire n_8287;
wire n_1904;
wire n_8111;
wire n_8341;
wire n_8830;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_7345;
wire n_8308;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_631;
wire n_8021;
wire n_1170;
wire n_2724;
wire n_8965;
wire n_2258;
wire n_7041;
wire n_6717;
wire n_7593;
wire n_8265;
wire n_898;
wire n_6881;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_5343;
wire n_6672;
wire n_7757;
wire n_1093;
wire n_8251;
wire n_7866;
wire n_6518;
wire n_7334;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_8773;
wire n_5947;
wire n_6242;
wire n_336;
wire n_6601;
wire n_8570;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_668;
wire n_8579;
wire n_2111;
wire n_3743;
wire n_8079;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_8506;
wire n_8973;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_8291;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_7758;
wire n_8320;
wire n_8635;
wire n_4472;
wire n_9118;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_291;
wire n_5180;
wire n_1640;
wire n_8375;
wire n_2973;
wire n_8612;
wire n_8778;
wire n_5893;
wire n_2710;
wire n_7705;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_9018;
wire n_5025;
wire n_2397;
wire n_8872;
wire n_240;
wire n_369;
wire n_7333;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_8006;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_8491;
wire n_8218;
wire n_1212;
wire n_7337;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_7439;
wire n_4371;
wire n_188;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_7210;
wire n_7744;
wire n_3898;
wire n_694;
wire n_6228;
wire n_6702;
wire n_7358;
wire n_8240;
wire n_4749;
wire n_7707;
wire n_5924;
wire n_1845;
wire n_7733;
wire n_921;
wire n_5545;
wire n_8458;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_8853;
wire n_5083;
wire n_7684;
wire n_3253;
wire n_8306;
wire n_2088;
wire n_1275;
wire n_6997;
wire n_4238;
wire n_6371;
wire n_904;
wire n_7673;
wire n_2005;
wire n_1696;
wire n_7187;
wire n_8013;
wire n_2108;
wire n_3824;
wire n_8342;
wire n_2246;
wire n_7313;
wire n_5899;
wire n_9012;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_3203;
wire n_383;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_6264;
wire n_5782;
wire n_8119;
wire n_9264;
wire n_630;
wire n_4168;
wire n_1369;
wire n_8582;
wire n_7036;
wire n_4298;
wire n_7370;
wire n_7931;
wire n_4743;
wire n_8445;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_8044;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_8363;
wire n_8464;
wire n_8921;
wire n_235;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_7480;
wire n_8843;
wire n_371;
wire n_5185;
wire n_8405;
wire n_2964;
wire n_8376;
wire n_308;
wire n_5032;
wire n_6990;
wire n_865;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_1041;
wire n_2451;
wire n_8694;
wire n_2913;
wire n_8848;
wire n_6288;
wire n_993;
wire n_1862;
wire n_3752;
wire n_8752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_8625;
wire n_8894;
wire n_7380;
wire n_2839;
wire n_8813;
wire n_3237;
wire n_7708;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_8430;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_8770;
wire n_6277;
wire n_8426;
wire n_5115;
wire n_7376;
wire n_8411;
wire n_902;
wire n_8817;
wire n_8461;
wire n_1723;
wire n_3918;
wire n_9230;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_596;
wire n_6409;
wire n_4095;
wire n_8391;
wire n_8507;
wire n_1310;
wire n_5927;
wire n_8691;
wire n_9188;
wire n_4485;
wire n_9032;
wire n_7657;
wire n_6388;
wire n_574;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_8967;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_9231;
wire n_6864;
wire n_1516;
wire n_4890;
wire n_8084;
wire n_8856;
wire n_2485;
wire n_6679;
wire n_8631;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_8219;
wire n_5507;
wire n_195;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_7504;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_8428;
wire n_9172;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_8338;
wire n_1631;
wire n_7602;
wire n_9180;
wire n_9017;
wire n_156;
wire n_9269;
wire n_6566;
wire n_9026;
wire n_1794;
wire n_5696;
wire n_7998;
wire n_8666;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_204;
wire n_7557;
wire n_3772;
wire n_7408;
wire n_2891;
wire n_496;
wire n_4335;
wire n_7026;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_7394;
wire n_263;
wire n_4516;
wire n_5235;
wire n_360;
wire n_1129;
wire n_7627;
wire n_6436;
wire n_1464;
wire n_7719;
wire n_2798;
wire n_7450;
wire n_165;
wire n_3217;
wire n_8938;
wire n_6081;
wire n_1249;
wire n_329;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_340;
wire n_3201;
wire n_7462;
wire n_7780;
wire n_3503;
wire n_8523;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_177;
wire n_364;
wire n_258;
wire n_7582;
wire n_5521;
wire n_431;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_8924;
wire n_2965;
wire n_4955;
wire n_7555;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_447;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_8380;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_841;
wire n_3204;
wire n_7451;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_5258;

INVx2_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_57),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_15),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_21),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_16),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_36),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_54),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_82),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_52),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_78),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_27),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_33),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_11),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_11),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_103),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_68),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_74),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_50),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_25),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_76),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_41),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_65),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_25),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_62),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_48),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_12),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_13),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_48),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_29),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_110),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_34),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_99),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_31),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_79),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_81),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_1),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_26),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_64),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_4),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_39),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_13),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_55),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_21),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_40),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_1),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_26),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_59),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_53),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_23),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_60),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_69),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_91),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_72),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_8),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_51),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_102),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_43),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_45),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_105),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_101),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_39),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_33),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_36),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_85),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_53),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_86),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_37),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_67),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_30),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_14),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_52),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_0),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_27),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_18),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_17),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_5),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_4),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_18),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_46),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_93),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_94),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_104),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_111),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_32),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_15),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_41),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_70),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_106),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_49),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_22),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_63),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_49),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_20),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_19),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_7),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_37),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_12),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_L g229 ( 
.A(n_134),
.B(n_0),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_133),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_129),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_138),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_L g233 ( 
.A(n_134),
.B(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_127),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_153),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_120),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_153),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_133),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_153),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_153),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_153),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_125),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_131),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_153),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_127),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_146),
.Y(n_251)
);

INVxp33_ASAP7_75t_SL g252 ( 
.A(n_123),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_146),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_123),
.B(n_2),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_134),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_150),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_135),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_186),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_150),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_239),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_251),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_241),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_247),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_116),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_230),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_251),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_248),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_243),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_254),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_253),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_252),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_117),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_252),
.Y(n_281)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_254),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_242),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_254),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_255),
.Y(n_290)
);

INVxp33_ASAP7_75t_SL g291 ( 
.A(n_255),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_235),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_235),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_235),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_253),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_256),
.Y(n_298)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_115),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_256),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

AND2x4_ASAP7_75t_SL g303 ( 
.A(n_268),
.B(n_204),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_233),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_256),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_259),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_259),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_233),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_284),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_261),
.A2(n_259),
.B(n_250),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_270),
.B(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

OAI22x1_ASAP7_75t_R g314 ( 
.A1(n_277),
.A2(n_183),
.B1(n_142),
.B2(n_220),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_265),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_283),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

OA21x2_ASAP7_75t_L g326 ( 
.A1(n_286),
.A2(n_245),
.B(n_244),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_266),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_250),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_282),
.A2(n_229),
.B1(n_162),
.B2(n_140),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_278),
.B(n_229),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_228),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_297),
.A2(n_140),
.B1(n_227),
.B2(n_226),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_296),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_298),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_277),
.A2(n_171),
.B1(n_225),
.B2(n_224),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_295),
.B(n_186),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_295),
.B(n_215),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_267),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_295),
.B(n_215),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_279),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_268),
.B(n_228),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_293),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_268),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_267),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_268),
.Y(n_357)
);

OA21x2_ASAP7_75t_L g358 ( 
.A1(n_280),
.A2(n_246),
.B(n_245),
.Y(n_358)
);

BUFx12f_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_280),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_289),
.A2(n_197),
.B1(n_175),
.B2(n_174),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_268),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_276),
.B(n_215),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_276),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_L g365 ( 
.A(n_272),
.B(n_119),
.Y(n_365)
);

NAND2x1_ASAP7_75t_L g366 ( 
.A(n_289),
.B(n_250),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_281),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_269),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_269),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_275),
.B(n_228),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_260),
.A2(n_154),
.B1(n_136),
.B2(n_144),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_275),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_260),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_262),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_262),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_292),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_294),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_294),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_264),
.B(n_139),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_294),
.Y(n_381)
);

XNOR2x2_ASAP7_75t_L g382 ( 
.A(n_297),
.B(n_118),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_294),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_294),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_290),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_294),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_261),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_261),
.A2(n_246),
.B(n_245),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_261),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_290),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_263),
.B(n_231),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_264),
.B(n_118),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_L g393 ( 
.A(n_265),
.B(n_126),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_268),
.B(n_147),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_294),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_260),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_290),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_292),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_264),
.B(n_122),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_264),
.B(n_139),
.Y(n_400)
);

NOR2x1_ASAP7_75t_L g401 ( 
.A(n_296),
.B(n_178),
.Y(n_401)
);

CKINVDCx8_ASAP7_75t_R g402 ( 
.A(n_265),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_261),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_264),
.B(n_231),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_282),
.A2(n_170),
.B1(n_169),
.B2(n_168),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_264),
.B(n_231),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_261),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_294),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_292),
.B(n_115),
.Y(n_409)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_292),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_260),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_294),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_261),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_261),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_261),
.A2(n_249),
.B(n_246),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_294),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_316),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_327),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_301),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_302),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_359),
.B(n_234),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_301),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_359),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_402),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_313),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_402),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_411),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_313),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_373),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_396),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_352),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_315),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_307),
.B(n_234),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_322),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_315),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_322),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_385),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_302),
.Y(n_438)
);

AND2x2_ASAP7_75t_SL g439 ( 
.A(n_303),
.B(n_115),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_332),
.B(n_178),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_317),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_335),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_385),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_353),
.A2(n_336),
.B1(n_308),
.B2(n_304),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_317),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_335),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_319),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_319),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_320),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_R g450 ( 
.A(n_365),
.B(n_130),
.Y(n_450)
);

OR2x6_ASAP7_75t_L g451 ( 
.A(n_366),
.B(n_234),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_390),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_390),
.Y(n_453)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_314),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_397),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_397),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_372),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_372),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_361),
.A2(n_202),
.B1(n_180),
.B2(n_165),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_372),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_314),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_372),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_342),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_372),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_372),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_303),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_303),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_R g468 ( 
.A(n_393),
.B(n_132),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_367),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_357),
.B(n_167),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_367),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_371),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_309),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_320),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_374),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_323),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_374),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_375),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_375),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_302),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_323),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_329),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_321),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_376),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_382),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_323),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_R g487 ( 
.A(n_309),
.B(n_137),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_SL g488 ( 
.A(n_357),
.B(n_151),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_377),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_382),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_335),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_336),
.B(n_339),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_338),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_368),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_321),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_368),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_368),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_R g498 ( 
.A(n_362),
.B(n_143),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_369),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_369),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_369),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_370),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_325),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_405),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_364),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_340),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_364),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_346),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_363),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_334),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_307),
.B(n_236),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_R g512 ( 
.A(n_362),
.B(n_145),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_R g513 ( 
.A(n_345),
.B(n_148),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_300),
.B(n_236),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_363),
.Y(n_515)
);

CKINVDCx6p67_ASAP7_75t_R g516 ( 
.A(n_363),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_363),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_357),
.B(n_167),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_370),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_345),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_345),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_300),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_325),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_348),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_R g525 ( 
.A(n_304),
.B(n_152),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_306),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_302),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_310),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_345),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_345),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_328),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_345),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_R g533 ( 
.A(n_304),
.B(n_156),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_348),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_338),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_348),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_310),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_354),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_354),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_354),
.B(n_158),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_350),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_350),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_R g543 ( 
.A(n_357),
.B(n_155),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_356),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_348),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_356),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_306),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_353),
.A2(n_176),
.B1(n_184),
.B2(n_196),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_349),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_344),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_339),
.B(n_164),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_328),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_360),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_337),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_343),
.B(n_181),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_360),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_337),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_333),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_391),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_333),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_344),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_310),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_391),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_392),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_330),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_349),
.B(n_236),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_392),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_392),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_330),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_387),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_344),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_392),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_387),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_338),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_399),
.B(n_122),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_330),
.Y(n_576)
);

AOI21x1_ASAP7_75t_L g577 ( 
.A1(n_389),
.A2(n_249),
.B(n_217),
.Y(n_577)
);

BUFx6f_ASAP7_75t_SL g578 ( 
.A(n_349),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_302),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_349),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_399),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_389),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_351),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_351),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_403),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_351),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_403),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_336),
.B(n_176),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_351),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_394),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_336),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_338),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_399),
.B(n_304),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_308),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_R g595 ( 
.A(n_357),
.B(n_157),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_407),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_407),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_308),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_308),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_338),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_399),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_343),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_SL g603 ( 
.A(n_357),
.B(n_191),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_R g604 ( 
.A(n_358),
.B(n_355),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_302),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_R g606 ( 
.A(n_338),
.B(n_159),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_347),
.B(n_184),
.Y(n_607)
);

AND3x2_ASAP7_75t_L g608 ( 
.A(n_347),
.B(n_124),
.C(n_198),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_347),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_341),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_341),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_R g612 ( 
.A(n_380),
.B(n_160),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_341),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_400),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_378),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_299),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_377),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_305),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_413),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_404),
.Y(n_620)
);

AOI21x1_ASAP7_75t_L g621 ( 
.A1(n_413),
.A2(n_249),
.B(n_206),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_414),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_414),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_406),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_378),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_299),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_299),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_299),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_378),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_299),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_401),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_299),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_377),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_379),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_299),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_366),
.B(n_193),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_318),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_299),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_409),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_379),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_401),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_379),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_381),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_381),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_312),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_381),
.Y(n_646)
);

CKINVDCx16_ASAP7_75t_R g647 ( 
.A(n_409),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_324),
.Y(n_648)
);

NOR2xp67_ASAP7_75t_L g649 ( 
.A(n_355),
.B(n_237),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_324),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_324),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_318),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_324),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_324),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_R g655 ( 
.A(n_398),
.B(n_355),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_324),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_331),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_318),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_331),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_383),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_383),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_331),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_331),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_331),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_358),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_331),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_383),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_384),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_358),
.Y(n_669)
);

NOR2xp67_ASAP7_75t_L g670 ( 
.A(n_384),
.B(n_237),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_409),
.Y(n_671)
);

CKINVDCx11_ASAP7_75t_R g672 ( 
.A(n_384),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_386),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_358),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_386),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_416),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_386),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_395),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_395),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_409),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_395),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_409),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_409),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_409),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_416),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_408),
.Y(n_686)
);

NOR2xp67_ASAP7_75t_L g687 ( 
.A(n_408),
.B(n_237),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_408),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_R g689 ( 
.A(n_398),
.B(n_163),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_410),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_442),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_618),
.B(n_409),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_442),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_L g694 ( 
.A(n_520),
.B(n_521),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_446),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_618),
.B(n_398),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_446),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_593),
.A2(n_490),
.B1(n_485),
.B2(n_601),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_491),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_620),
.B(n_398),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_491),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_614),
.B(n_410),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_434),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_419),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_422),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_616),
.Y(n_706)
);

NOR2x1p5_ASAP7_75t_L g707 ( 
.A(n_423),
.B(n_124),
.Y(n_707)
);

NAND3xp33_ASAP7_75t_L g708 ( 
.A(n_417),
.B(n_318),
.C(n_199),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_626),
.Y(n_709)
);

INVx5_ASAP7_75t_L g710 ( 
.A(n_616),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_620),
.B(n_412),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_425),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_616),
.Y(n_713)
);

BUFx4f_ASAP7_75t_L g714 ( 
.A(n_593),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_428),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_420),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_432),
.Y(n_717)
);

INVx5_ASAP7_75t_L g718 ( 
.A(n_671),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_435),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_614),
.B(n_410),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_535),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_624),
.B(n_412),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_430),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_441),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_418),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_445),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_591),
.B(n_318),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_469),
.B(n_410),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_624),
.B(n_412),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_417),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_447),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_690),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_420),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_591),
.B(n_601),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_448),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_528),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_449),
.Y(n_737)
);

INVx5_ASAP7_75t_L g738 ( 
.A(n_671),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_609),
.B(n_602),
.Y(n_739)
);

INVx5_ASAP7_75t_L g740 ( 
.A(n_671),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_524),
.B(n_318),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_439),
.A2(n_416),
.B1(n_204),
.B2(n_211),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_609),
.B(n_410),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_L g744 ( 
.A(n_529),
.B(n_200),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_592),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_564),
.A2(n_196),
.B1(n_206),
.B2(n_217),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_528),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_469),
.B(n_201),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_538),
.B(n_203),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_424),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_474),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_537),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_566),
.B(n_311),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_483),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_602),
.B(n_311),
.Y(n_755)
);

OAI21xp33_ASAP7_75t_SL g756 ( 
.A1(n_444),
.A2(n_415),
.B(n_198),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_476),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_424),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_439),
.A2(n_204),
.B1(n_211),
.B2(n_195),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_539),
.B(n_205),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_594),
.A2(n_204),
.B1(n_211),
.B2(n_195),
.Y(n_761)
);

NOR2x1p5_ASAP7_75t_L g762 ( 
.A(n_423),
.B(n_149),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_495),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_537),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_471),
.B(n_207),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_420),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_476),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_503),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_562),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_562),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_631),
.B(n_222),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_426),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_565),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_523),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_567),
.A2(n_223),
.B1(n_189),
.B2(n_185),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_645),
.B(n_149),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_420),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_535),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_440),
.B(n_610),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_574),
.Y(n_780)
);

INVx6_ASAP7_75t_L g781 ( 
.A(n_574),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_594),
.B(n_172),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_600),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_568),
.A2(n_190),
.B1(n_189),
.B2(n_166),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_426),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_565),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_610),
.B(n_161),
.Y(n_787)
);

BUFx10_ASAP7_75t_L g788 ( 
.A(n_429),
.Y(n_788)
);

XNOR2xp5_ASAP7_75t_L g789 ( 
.A(n_461),
.B(n_161),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_531),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_611),
.B(n_166),
.Y(n_791)
);

BUFx10_ASAP7_75t_L g792 ( 
.A(n_429),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_552),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_598),
.B(n_177),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_598),
.B(n_179),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_599),
.A2(n_211),
.B1(n_185),
.B2(n_190),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_534),
.B(n_238),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_569),
.Y(n_798)
);

XOR2xp5_ASAP7_75t_L g799 ( 
.A(n_427),
.B(n_326),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_566),
.B(n_238),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_569),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_600),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_599),
.B(n_572),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_626),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_536),
.B(n_238),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_581),
.A2(n_510),
.B1(n_506),
.B2(n_575),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_576),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_611),
.B(n_209),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_476),
.Y(n_809)
);

AND2x6_ASAP7_75t_L g810 ( 
.A(n_647),
.B(n_218),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_550),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_613),
.B(n_209),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_522),
.B(n_326),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_575),
.A2(n_214),
.B1(n_216),
.B2(n_219),
.Y(n_814)
);

CKINVDCx16_ASAP7_75t_R g815 ( 
.A(n_463),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_466),
.B(n_182),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_466),
.B(n_210),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_431),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_558),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_451),
.B(n_388),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_576),
.Y(n_821)
);

AND2x6_ASAP7_75t_L g822 ( 
.A(n_575),
.B(n_218),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_615),
.Y(n_823)
);

INVxp33_ASAP7_75t_L g824 ( 
.A(n_487),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_561),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_617),
.Y(n_826)
);

INVx6_ASAP7_75t_L g827 ( 
.A(n_617),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_526),
.A2(n_214),
.B1(n_216),
.B2(n_219),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_502),
.B(n_388),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_547),
.A2(n_128),
.B1(n_141),
.B2(n_213),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_481),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_627),
.Y(n_832)
);

INVx6_ASAP7_75t_L g833 ( 
.A(n_420),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_438),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_508),
.A2(n_128),
.B1(n_141),
.B2(n_213),
.Y(n_835)
);

INVx4_ASAP7_75t_L g836 ( 
.A(n_627),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_615),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_430),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_481),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_560),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_628),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_452),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_545),
.B(n_504),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_570),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_573),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_557),
.B(n_388),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_582),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_519),
.B(n_388),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_438),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_585),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_467),
.B(n_187),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_587),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_481),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_596),
.Y(n_854)
);

INVx4_ASAP7_75t_SL g855 ( 
.A(n_470),
.Y(n_855)
);

AND2x2_ASAP7_75t_SL g856 ( 
.A(n_680),
.B(n_326),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_559),
.B(n_326),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_580),
.B(n_415),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_597),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_619),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_571),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_584),
.B(n_221),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_457),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_613),
.B(n_212),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_514),
.B(n_192),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_622),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_457),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_514),
.B(n_433),
.Y(n_868)
);

AND2x2_ASAP7_75t_SL g869 ( 
.A(n_684),
.B(n_121),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_L g870 ( 
.A(n_459),
.B(n_188),
.C(n_213),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_623),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_456),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_467),
.B(n_173),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_584),
.B(n_2),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_625),
.Y(n_875)
);

OR2x6_ASAP7_75t_L g876 ( 
.A(n_451),
.B(n_173),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_458),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_586),
.B(n_3),
.Y(n_878)
);

BUFx10_ASAP7_75t_L g879 ( 
.A(n_578),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_458),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_629),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_643),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_634),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_438),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_433),
.B(n_3),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_482),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_643),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_438),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_678),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_586),
.B(n_5),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_460),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_511),
.B(n_6),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_589),
.B(n_6),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_589),
.B(n_173),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_678),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_640),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_642),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_578),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_511),
.B(n_7),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_436),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_R g901 ( 
.A(n_431),
.B(n_530),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_492),
.A2(n_578),
.B1(n_669),
.B2(n_674),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_563),
.B(n_141),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_628),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_641),
.B(n_9),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_551),
.B(n_9),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_644),
.Y(n_907)
);

INVxp67_ASAP7_75t_SL g908 ( 
.A(n_493),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_460),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_630),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_532),
.B(n_128),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_549),
.B(n_127),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_555),
.B(n_10),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_646),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_665),
.A2(n_121),
.B1(n_16),
.B2(n_17),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_462),
.Y(n_916)
);

INVx4_ASAP7_75t_SL g917 ( 
.A(n_470),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_473),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_509),
.B(n_121),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_486),
.Y(n_920)
);

BUFx8_ASAP7_75t_SL g921 ( 
.A(n_436),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_525),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_540),
.B(n_10),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_660),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_462),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_661),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_667),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_583),
.B(n_421),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_677),
.Y(n_929)
);

OR2x6_ASAP7_75t_L g930 ( 
.A(n_451),
.B(n_121),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_554),
.B(n_19),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_451),
.B(n_588),
.Y(n_932)
);

INVxp33_ASAP7_75t_SL g933 ( 
.A(n_437),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_516),
.A2(n_121),
.B1(n_22),
.B2(n_23),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_548),
.B(n_20),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_515),
.B(n_517),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_437),
.B(n_24),
.Y(n_937)
);

INVx5_ASAP7_75t_L g938 ( 
.A(n_438),
.Y(n_938)
);

CKINVDCx16_ASAP7_75t_R g939 ( 
.A(n_533),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_464),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_480),
.B(n_527),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_630),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_480),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_676),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_480),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_685),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_464),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_443),
.B(n_24),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_443),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_679),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_453),
.Y(n_951)
);

BUFx8_ASAP7_75t_SL g952 ( 
.A(n_453),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_516),
.A2(n_121),
.B1(n_30),
.B2(n_31),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_L g954 ( 
.A(n_505),
.B(n_28),
.C(n_32),
.Y(n_954)
);

AND2x6_ASAP7_75t_L g955 ( 
.A(n_486),
.B(n_56),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_681),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_486),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_686),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_507),
.B(n_28),
.Y(n_959)
);

INVx4_ASAP7_75t_SL g960 ( 
.A(n_470),
.Y(n_960)
);

BUFx4f_ASAP7_75t_L g961 ( 
.A(n_470),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_657),
.B(n_34),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_688),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_489),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_455),
.B(n_35),
.Y(n_965)
);

NOR3xp33_ASAP7_75t_L g966 ( 
.A(n_455),
.B(n_35),
.C(n_38),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_480),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_670),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_632),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_687),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_659),
.B(n_38),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_607),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_668),
.B(n_40),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_454),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_472),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_632),
.Y(n_976)
);

AND2x6_ASAP7_75t_L g977 ( 
.A(n_489),
.B(n_80),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_465),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_673),
.B(n_47),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_480),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_527),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_527),
.B(n_579),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_465),
.B(n_47),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_494),
.B(n_50),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_489),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_633),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_662),
.B(n_51),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_675),
.B(n_61),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_484),
.B(n_66),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_496),
.B(n_497),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_527),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_633),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_499),
.A2(n_71),
.B1(n_73),
.B2(n_75),
.Y(n_993)
);

AND2x6_ASAP7_75t_L g994 ( 
.A(n_633),
.B(n_83),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_577),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_621),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_527),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_663),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_541),
.B(n_87),
.Y(n_999)
);

INVxp67_ASAP7_75t_SL g1000 ( 
.A(n_579),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_579),
.Y(n_1001)
);

CKINVDCx6p67_ASAP7_75t_R g1002 ( 
.A(n_672),
.Y(n_1002)
);

BUFx4f_ASAP7_75t_L g1003 ( 
.A(n_470),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_664),
.B(n_88),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_579),
.Y(n_1005)
);

NAND2xp33_ASAP7_75t_SL g1006 ( 
.A(n_655),
.B(n_666),
.Y(n_1006)
);

BUFx4f_ASAP7_75t_L g1007 ( 
.A(n_470),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_500),
.A2(n_501),
.B1(n_553),
.B2(n_546),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_475),
.B(n_97),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_635),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_579),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_605),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_SL g1013 ( 
.A(n_477),
.B(n_112),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_542),
.B(n_556),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_450),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_544),
.B(n_98),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_478),
.B(n_100),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_479),
.B(n_590),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_605),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_605),
.Y(n_1020)
);

AO22x2_ASAP7_75t_L g1021 ( 
.A1(n_636),
.A2(n_608),
.B1(n_604),
.B2(n_590),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_605),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_605),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_648),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_650),
.B(n_651),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_653),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_635),
.B(n_639),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_612),
.B(n_656),
.Y(n_1028)
);

INVx5_ASAP7_75t_L g1029 ( 
.A(n_637),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_638),
.B(n_683),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_637),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_637),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_638),
.B(n_639),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_637),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_779),
.B(n_739),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_906),
.A2(n_649),
.B(n_488),
.C(n_603),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_868),
.B(n_797),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_933),
.B(n_654),
.Y(n_1038)
);

NAND2xp33_ASAP7_75t_SL g1039 ( 
.A(n_901),
.B(n_498),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_797),
.B(n_468),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_714),
.B(n_606),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_L g1042 ( 
.A(n_748),
.B(n_765),
.C(n_959),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_691),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_797),
.B(n_512),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_745),
.B(n_829),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_691),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_714),
.B(n_1014),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_714),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_933),
.B(n_683),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_805),
.B(n_513),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_1030),
.B(n_1027),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_SL g1052 ( 
.A(n_870),
.B(n_689),
.C(n_543),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_805),
.B(n_518),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_818),
.B(n_682),
.Y(n_1054)
);

NAND3xp33_ASAP7_75t_L g1055 ( 
.A(n_923),
.B(n_637),
.C(n_652),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_736),
.Y(n_1056)
);

AND2x6_ASAP7_75t_SL g1057 ( 
.A(n_1018),
.B(n_595),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_SL g1058 ( 
.A(n_750),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_818),
.B(n_682),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_1025),
.B(n_658),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_941),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_900),
.B(n_652),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_747),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1030),
.B(n_652),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_805),
.B(n_518),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_949),
.B(n_652),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_693),
.Y(n_1067)
);

NOR2xp67_ASAP7_75t_L g1068 ( 
.A(n_938),
.B(n_652),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_725),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_1030),
.B(n_1027),
.Y(n_1070)
);

AO221x1_ASAP7_75t_L g1071 ( 
.A1(n_1021),
.A2(n_518),
.B1(n_658),
.B2(n_784),
.C(n_775),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_1008),
.B(n_658),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_799),
.A2(n_518),
.B1(n_658),
.B2(n_698),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_693),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_990),
.B(n_658),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_747),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_728),
.B(n_518),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_702),
.B(n_518),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_703),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_720),
.B(n_787),
.Y(n_1080)
);

INVx6_ASAP7_75t_L g1081 ( 
.A(n_879),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_867),
.B(n_909),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_791),
.B(n_808),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_812),
.B(n_800),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_800),
.B(n_857),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_867),
.B(n_909),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_811),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_695),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_916),
.B(n_940),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_916),
.B(n_940),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_752),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_695),
.Y(n_1092)
);

NAND2x1_ASAP7_75t_L g1093 ( 
.A(n_941),
.B(n_982),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_944),
.B(n_946),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_938),
.B(n_1020),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_978),
.B(n_863),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_696),
.A2(n_700),
.B(n_1006),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_990),
.B(n_951),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_978),
.B(n_863),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_776),
.B(n_972),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_951),
.B(n_872),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_972),
.B(n_704),
.Y(n_1102)
);

INVxp33_ASAP7_75t_L g1103 ( 
.A(n_723),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_838),
.B(n_824),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_704),
.B(n_705),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_705),
.B(n_712),
.Y(n_1106)
);

AO22x2_ASAP7_75t_L g1107 ( 
.A1(n_799),
.A2(n_1021),
.B1(n_846),
.B2(n_848),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_SL g1108 ( 
.A(n_730),
.B(n_975),
.C(n_965),
.Y(n_1108)
);

NOR2x1p5_ASAP7_75t_L g1109 ( 
.A(n_1002),
.B(n_772),
.Y(n_1109)
);

NAND2xp33_ASAP7_75t_L g1110 ( 
.A(n_913),
.B(n_716),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_846),
.A2(n_731),
.B1(n_735),
.B2(n_712),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_697),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_877),
.B(n_880),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_877),
.B(n_880),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_752),
.Y(n_1115)
);

INVx8_ASAP7_75t_L g1116 ( 
.A(n_930),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_764),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_891),
.B(n_925),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_891),
.B(n_925),
.Y(n_1119)
);

INVx8_ASAP7_75t_L g1120 ( 
.A(n_930),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_857),
.B(n_753),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_731),
.B(n_735),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_697),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_737),
.B(n_751),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_737),
.B(n_751),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_930),
.B(n_932),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_764),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_754),
.B(n_763),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_947),
.B(n_730),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_947),
.B(n_772),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_699),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_769),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_SL g1133 ( 
.A(n_750),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_754),
.B(n_763),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_753),
.B(n_768),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_769),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_768),
.B(n_774),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_699),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_774),
.B(n_790),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_770),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_701),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_822),
.A2(n_878),
.B1(n_890),
.B2(n_874),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_701),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_770),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_773),
.Y(n_1145)
);

NOR3xp33_ASAP7_75t_L g1146 ( 
.A(n_954),
.B(n_966),
.C(n_862),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_773),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_875),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_875),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_790),
.B(n_793),
.Y(n_1150)
);

NAND2xp33_ASAP7_75t_L g1151 ( 
.A(n_716),
.B(n_733),
.Y(n_1151)
);

O2A1O1Ixp5_ASAP7_75t_L g1152 ( 
.A1(n_973),
.A2(n_979),
.B(n_727),
.C(n_892),
.Y(n_1152)
);

AO22x2_ASAP7_75t_L g1153 ( 
.A1(n_1021),
.A2(n_848),
.B1(n_829),
.B2(n_983),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_793),
.B(n_840),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_786),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_SL g1156 ( 
.A(n_750),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1006),
.A2(n_964),
.B(n_755),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_941),
.Y(n_1158)
);

INVx8_ASAP7_75t_L g1159 ( 
.A(n_930),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_886),
.B(n_1015),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_827),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_840),
.B(n_844),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1015),
.B(n_785),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_785),
.B(n_771),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_786),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_798),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_881),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_941),
.Y(n_1168)
);

NOR2xp67_ASAP7_75t_SL g1169 ( 
.A(n_938),
.B(n_1020),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_716),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1033),
.B(n_938),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_R g1172 ( 
.A(n_725),
.B(n_842),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_734),
.B(n_842),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_918),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_743),
.A2(n_1000),
.B(n_982),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_881),
.Y(n_1176)
);

BUFx12f_ASAP7_75t_L g1177 ( 
.A(n_758),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_883),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_893),
.B(n_922),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_827),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_998),
.B(n_1028),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_883),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_R g1183 ( 
.A(n_815),
.B(n_758),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_844),
.B(n_845),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1021),
.A2(n_810),
.B1(n_806),
.B2(n_822),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_845),
.B(n_847),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_798),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_L g1188 ( 
.A(n_938),
.B(n_1020),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_801),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_847),
.B(n_850),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_827),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_801),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_850),
.A2(n_854),
.B1(n_859),
.B2(n_852),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_897),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_807),
.Y(n_1195)
);

AO221x1_ASAP7_75t_L g1196 ( 
.A1(n_716),
.A2(n_884),
.B1(n_945),
.B2(n_888),
.C(n_943),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_827),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_843),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_998),
.B(n_928),
.Y(n_1199)
);

OAI22x1_ASAP7_75t_SL g1200 ( 
.A1(n_789),
.A2(n_921),
.B1(n_952),
.B2(n_1002),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_903),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_852),
.B(n_854),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_859),
.B(n_860),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_803),
.B(n_864),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_897),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_781),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_937),
.B(n_948),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_914),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_822),
.A2(n_935),
.B1(n_984),
.B2(n_905),
.Y(n_1209)
);

NOR2x1p5_ASAP7_75t_L g1210 ( 
.A(n_811),
.B(n_825),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_860),
.B(n_866),
.Y(n_1211)
);

NOR2x1p5_ASAP7_75t_L g1212 ( 
.A(n_825),
.B(n_861),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_866),
.B(n_871),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_810),
.A2(n_822),
.B1(n_759),
.B2(n_984),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_928),
.B(n_758),
.Y(n_1215)
);

OR2x6_ASAP7_75t_L g1216 ( 
.A(n_932),
.B(n_876),
.Y(n_1216)
);

BUFx8_ASAP7_75t_L g1217 ( 
.A(n_861),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_871),
.B(n_711),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_745),
.B(n_722),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_810),
.A2(n_822),
.B1(n_869),
.B2(n_902),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_813),
.B(n_715),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_807),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_821),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_732),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_928),
.B(n_1009),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_716),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_729),
.B(n_717),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_719),
.B(n_724),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_937),
.B(n_948),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_921),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_914),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_903),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_924),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1017),
.A2(n_692),
.B(n_756),
.C(n_1016),
.Y(n_1234)
);

AND2x6_ASAP7_75t_L g1235 ( 
.A(n_1033),
.B(n_706),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1009),
.B(n_1024),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_726),
.B(n_819),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_732),
.Y(n_1238)
);

NAND2xp33_ASAP7_75t_L g1239 ( 
.A(n_733),
.B(n_766),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1026),
.B(n_788),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_936),
.B(n_952),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_788),
.B(n_792),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_924),
.Y(n_1243)
);

NOR2xp67_ASAP7_75t_SL g1244 ( 
.A(n_1020),
.B(n_1029),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_926),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_865),
.B(n_814),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_989),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_926),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_788),
.B(n_792),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_929),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_749),
.B(n_760),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1020),
.B(n_1029),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_810),
.A2(n_822),
.B1(n_869),
.B2(n_939),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_989),
.B(n_873),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_823),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_792),
.B(n_782),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_999),
.A2(n_746),
.B(n_899),
.C(n_885),
.Y(n_1257)
);

NAND2xp33_ASAP7_75t_L g1258 ( 
.A(n_733),
.B(n_766),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_794),
.B(n_795),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_983),
.B(n_912),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_741),
.B(n_709),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_931),
.B(n_894),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_741),
.B(n_709),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_912),
.B(n_810),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_741),
.B(n_709),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_929),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_804),
.B(n_832),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_963),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_915),
.A2(n_1013),
.B1(n_810),
.B2(n_744),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_912),
.B(n_744),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_961),
.A2(n_1003),
.B(n_1007),
.C(n_988),
.Y(n_1271)
);

OAI221xp5_ASAP7_75t_L g1272 ( 
.A1(n_828),
.A2(n_974),
.B1(n_796),
.B2(n_953),
.C(n_934),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_835),
.A2(n_742),
.B1(n_830),
.B2(n_789),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_813),
.B(n_963),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_694),
.B(n_896),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_804),
.B(n_832),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_816),
.B(n_817),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_823),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_837),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_694),
.B(n_896),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_851),
.B(n_781),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_982),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_907),
.B(n_927),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_804),
.B(n_832),
.Y(n_1284)
);

INVxp67_ASAP7_75t_SL g1285 ( 
.A(n_908),
.Y(n_1285)
);

INVxp67_ASAP7_75t_L g1286 ( 
.A(n_962),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_971),
.A2(n_987),
.B(n_986),
.C(n_985),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_907),
.B(n_927),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_950),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_950),
.B(n_956),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_836),
.A2(n_976),
.B1(n_1010),
.B2(n_969),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_956),
.B(n_958),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_836),
.B(n_841),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_932),
.B(n_876),
.Y(n_1294)
);

NAND2xp33_ASAP7_75t_L g1295 ( 
.A(n_733),
.B(n_766),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_958),
.B(n_761),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_802),
.B(n_826),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_836),
.B(n_841),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_837),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_882),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_841),
.B(n_904),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_802),
.B(n_826),
.Y(n_1302)
);

OR2x6_ASAP7_75t_L g1303 ( 
.A(n_932),
.B(n_876),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_882),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_876),
.B(n_856),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_780),
.B(n_887),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_887),
.B(n_889),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_858),
.A2(n_762),
.B1(n_707),
.B2(n_820),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_968),
.A2(n_970),
.B1(n_856),
.B2(n_895),
.Y(n_1309)
);

OAI221xp5_ASAP7_75t_L g1310 ( 
.A1(n_993),
.A2(n_961),
.B1(n_1003),
.B2(n_1007),
.C(n_708),
.Y(n_1310)
);

NOR2x1p5_ASAP7_75t_L g1311 ( 
.A(n_904),
.B(n_910),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_889),
.B(n_895),
.Y(n_1312)
);

OAI221xp5_ASAP7_75t_L g1313 ( 
.A1(n_961),
.A2(n_1007),
.B1(n_1003),
.B2(n_968),
.C(n_970),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_904),
.B(n_910),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_858),
.B(n_982),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_985),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_733),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_781),
.B(n_1005),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_R g1319 ( 
.A(n_879),
.B(n_898),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_910),
.B(n_942),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_942),
.B(n_976),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_781),
.B(n_1011),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_942),
.B(n_969),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_721),
.B(n_783),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_879),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_721),
.B(n_783),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_858),
.B(n_820),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_986),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1005),
.B(n_1011),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_778),
.B(n_920),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_757),
.Y(n_1331)
);

NOR2x1p5_ASAP7_75t_L g1332 ( 
.A(n_969),
.B(n_976),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1010),
.A2(n_833),
.B1(n_1029),
.B2(n_920),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_757),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_778),
.B(n_920),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1031),
.B(n_1032),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1029),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_820),
.B(n_957),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_757),
.B(n_957),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1010),
.B(n_1029),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_767),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_767),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_767),
.B(n_957),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_766),
.B(n_943),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_820),
.A2(n_919),
.B1(n_994),
.B2(n_977),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_809),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1031),
.A2(n_1032),
.B(n_1004),
.C(n_853),
.Y(n_1347)
);

BUFx4f_ASAP7_75t_L g1348 ( 
.A(n_955),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_809),
.B(n_992),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_809),
.B(n_992),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_710),
.B(n_718),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_831),
.Y(n_1352)
);

BUFx5_ASAP7_75t_L g1353 ( 
.A(n_955),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_831),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_898),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_L g1356 ( 
.A1(n_995),
.A2(n_996),
.B(n_1023),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_831),
.B(n_853),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_766),
.B(n_945),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_839),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_SL g1360 ( 
.A(n_777),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_710),
.B(n_718),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_839),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_839),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_898),
.A2(n_911),
.B1(n_1023),
.B2(n_1022),
.Y(n_1364)
);

NAND2xp33_ASAP7_75t_L g1365 ( 
.A(n_777),
.B(n_849),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_853),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_992),
.B(n_997),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_995),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_777),
.B(n_888),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_777),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_996),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_777),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_834),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_833),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_834),
.B(n_943),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_834),
.B(n_943),
.Y(n_1376)
);

INVxp33_ASAP7_75t_L g1377 ( 
.A(n_980),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_980),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_981),
.A2(n_1034),
.B1(n_1022),
.B2(n_1019),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_981),
.A2(n_1034),
.B1(n_1019),
.B2(n_1012),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_997),
.B(n_1001),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_991),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_991),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_1001),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1012),
.A2(n_960),
.B1(n_917),
.B2(n_855),
.Y(n_1385)
);

NOR3xp33_ASAP7_75t_L g1386 ( 
.A(n_997),
.B(n_706),
.C(n_713),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_955),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_955),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_955),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_834),
.B(n_884),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_834),
.B(n_884),
.Y(n_1391)
);

INVx8_ASAP7_75t_L g1392 ( 
.A(n_955),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_849),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_833),
.B(n_884),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_855),
.B(n_917),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_849),
.B(n_884),
.Y(n_1396)
);

NAND3xp33_ASAP7_75t_SL g1397 ( 
.A(n_977),
.B(n_994),
.C(n_855),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_849),
.B(n_888),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_977),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_849),
.B(n_888),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_888),
.B(n_967),
.Y(n_1401)
);

NAND2xp33_ASAP7_75t_SL g1402 ( 
.A(n_943),
.B(n_967),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_945),
.B(n_967),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_945),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_855),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_945),
.B(n_967),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_967),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_833),
.B(n_960),
.Y(n_1408)
);

AOI221xp5_ASAP7_75t_L g1409 ( 
.A1(n_706),
.A2(n_713),
.B1(n_960),
.B2(n_917),
.C(n_738),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_713),
.B(n_710),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_917),
.B(n_960),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_977),
.B(n_994),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_977),
.B(n_994),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_710),
.B(n_718),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_977),
.B(n_994),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_710),
.B(n_718),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_994),
.A2(n_740),
.B(n_718),
.C(n_738),
.Y(n_1417)
);

AO22x2_ASAP7_75t_L g1418 ( 
.A1(n_738),
.A2(n_799),
.B1(n_382),
.B2(n_1021),
.Y(n_1418)
);

NOR2xp67_ASAP7_75t_L g1419 ( 
.A(n_738),
.B(n_740),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_738),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_740),
.B(n_593),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_740),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_740),
.A2(n_601),
.B1(n_868),
.B2(n_567),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_736),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_716),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_779),
.B(n_618),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_736),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_779),
.B(n_618),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_779),
.B(n_618),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_736),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_691),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_691),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1030),
.B(n_1027),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_779),
.B(n_618),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_799),
.A2(n_485),
.B1(n_490),
.B2(n_382),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_714),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_739),
.A2(n_601),
.B1(n_567),
.B2(n_568),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_736),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_691),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_779),
.B(n_618),
.Y(n_1440)
);

OAI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_748),
.A2(n_334),
.B1(n_959),
.B2(n_281),
.C(n_279),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_691),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_739),
.B(n_279),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_868),
.A2(n_601),
.B1(n_567),
.B2(n_568),
.Y(n_1444)
);

BUFx5_ASAP7_75t_L g1445 ( 
.A(n_955),
.Y(n_1445)
);

INVx8_ASAP7_75t_L g1446 ( 
.A(n_930),
.Y(n_1446)
);

INVxp67_ASAP7_75t_L g1447 ( 
.A(n_703),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_739),
.B(n_469),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_739),
.B(n_279),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_779),
.B(n_618),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_691),
.Y(n_1451)
);

NAND2xp33_ASAP7_75t_L g1452 ( 
.A(n_923),
.B(n_357),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_779),
.B(n_618),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_739),
.B(n_469),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_714),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_703),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_739),
.B(n_469),
.Y(n_1457)
);

O2A1O1Ixp5_ASAP7_75t_L g1458 ( 
.A1(n_923),
.A2(n_913),
.B(n_906),
.C(n_488),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1030),
.B(n_1027),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_739),
.B(n_279),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_739),
.B(n_469),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_799),
.A2(n_485),
.B1(n_490),
.B2(n_382),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_703),
.Y(n_1463)
);

OAI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_739),
.A2(n_601),
.B1(n_567),
.B2(n_568),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_739),
.B(n_279),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_739),
.B(n_279),
.Y(n_1466)
);

NAND2x1p5_ASAP7_75t_L g1467 ( 
.A(n_938),
.B(n_1020),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_714),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_868),
.A2(n_601),
.B1(n_567),
.B2(n_568),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_739),
.A2(n_601),
.B1(n_567),
.B2(n_568),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_739),
.B(n_469),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1030),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_714),
.B(n_593),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_779),
.B(n_618),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_779),
.B(n_618),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_739),
.B(n_279),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_691),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_799),
.A2(n_485),
.B1(n_490),
.B2(n_382),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_779),
.B(n_618),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_736),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1030),
.B(n_1027),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_779),
.B(n_618),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_941),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_SL g1484 ( 
.A(n_750),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_691),
.Y(n_1485)
);

NAND2xp33_ASAP7_75t_L g1486 ( 
.A(n_923),
.B(n_357),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_779),
.B(n_618),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_703),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_725),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_691),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_779),
.B(n_618),
.Y(n_1491)
);

INVxp67_ASAP7_75t_SL g1492 ( 
.A(n_1025),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_779),
.B(n_618),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_736),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_779),
.B(n_618),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_L g1496 ( 
.A(n_923),
.B(n_357),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_703),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_779),
.B(n_618),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_739),
.B(n_469),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_739),
.A2(n_601),
.B1(n_567),
.B2(n_568),
.Y(n_1500)
);

INVx8_ASAP7_75t_L g1501 ( 
.A(n_930),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_779),
.B(n_618),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_691),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_779),
.B(n_618),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_739),
.B(n_279),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_736),
.Y(n_1506)
);

AO221x1_ASAP7_75t_L g1507 ( 
.A1(n_1021),
.A2(n_361),
.B1(n_784),
.B2(n_459),
.C(n_372),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_739),
.B(n_469),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_691),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_779),
.B(n_618),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_739),
.A2(n_601),
.B1(n_567),
.B2(n_568),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_739),
.B(n_279),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_739),
.A2(n_601),
.B1(n_567),
.B2(n_568),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_714),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_779),
.B(n_618),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_714),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_779),
.B(n_618),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_990),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_691),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_691),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_779),
.B(n_618),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_736),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_799),
.A2(n_485),
.B1(n_490),
.B2(n_382),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1142),
.B(n_1209),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1061),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1368),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1142),
.A2(n_1042),
.B1(n_1209),
.B2(n_1207),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1084),
.A2(n_1269),
.B1(n_1037),
.B2(n_1348),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1418),
.A2(n_1435),
.B1(n_1478),
.B2(n_1462),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1111),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1121),
.B(n_1274),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1121),
.B(n_1221),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1269),
.A2(n_1348),
.B1(n_1106),
.B2(n_1122),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1257),
.A2(n_1441),
.B(n_1428),
.C(n_1429),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1221),
.B(n_1154),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1315),
.B(n_1327),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1080),
.B(n_1198),
.Y(n_1539)
);

O2A1O1Ixp5_ASAP7_75t_L g1540 ( 
.A1(n_1458),
.A2(n_1152),
.B(n_1234),
.C(n_1060),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1315),
.B(n_1327),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1348),
.A2(n_1124),
.B1(n_1125),
.B2(n_1105),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1418),
.A2(n_1523),
.B1(n_1507),
.B2(n_1071),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1154),
.B(n_1102),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1061),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1452),
.A2(n_1496),
.B(n_1486),
.Y(n_1546)
);

CKINVDCx8_ASAP7_75t_R g1547 ( 
.A(n_1057),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1399),
.B(n_1353),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1218),
.B(n_1128),
.Y(n_1549)
);

NOR2x2_ASAP7_75t_L g1550 ( 
.A(n_1200),
.B(n_1172),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1229),
.A2(n_1108),
.B1(n_1164),
.B2(n_1272),
.Y(n_1551)
);

NOR3xp33_ASAP7_75t_L g1552 ( 
.A(n_1146),
.B(n_1449),
.C(n_1443),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1426),
.A2(n_1434),
.B(n_1450),
.C(n_1440),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1043),
.Y(n_1554)
);

INVx5_ASAP7_75t_L g1555 ( 
.A(n_1392),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1196),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1134),
.B(n_1137),
.Y(n_1557)
);

AND2x6_ASAP7_75t_SL g1558 ( 
.A(n_1163),
.B(n_1160),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1061),
.B(n_1282),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1043),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1046),
.Y(n_1561)
);

NOR2x2_ASAP7_75t_L g1562 ( 
.A(n_1200),
.B(n_1183),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1139),
.B(n_1150),
.Y(n_1563)
);

O2A1O1Ixp5_ASAP7_75t_L g1564 ( 
.A1(n_1072),
.A2(n_1097),
.B(n_1157),
.C(n_1036),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1392),
.Y(n_1565)
);

OAI22x1_ASAP7_75t_L g1566 ( 
.A1(n_1308),
.A2(n_1418),
.B1(n_1345),
.B2(n_1437),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1282),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1162),
.B(n_1184),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_SL g1569 ( 
.A1(n_1418),
.A2(n_1507),
.B1(n_1071),
.B2(n_1107),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1399),
.B(n_1353),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1368),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1069),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1196),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1368),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1453),
.B(n_1474),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1186),
.B(n_1190),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1518),
.Y(n_1577)
);

NOR2xp67_ASAP7_75t_SL g1578 ( 
.A(n_1310),
.B(n_1177),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1046),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1305),
.B(n_1338),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1392),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1067),
.Y(n_1582)
);

INVx5_ASAP7_75t_L g1583 ( 
.A(n_1392),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_SL g1584 ( 
.A(n_1437),
.B(n_1500),
.C(n_1470),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1107),
.A2(n_1185),
.B1(n_1153),
.B2(n_1273),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1202),
.B(n_1203),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1392),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1470),
.B(n_1500),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1067),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1415),
.A2(n_1055),
.B(n_1347),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1371),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1211),
.B(n_1213),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1252),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1100),
.B(n_1083),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1227),
.B(n_1148),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1045),
.B(n_1305),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1252),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1148),
.B(n_1149),
.Y(n_1598)
);

NAND2x1p5_ASAP7_75t_L g1599 ( 
.A(n_1387),
.B(n_1388),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1149),
.B(n_1167),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1513),
.B(n_1464),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1069),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1074),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1338),
.B(n_1074),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1371),
.Y(n_1605)
);

NAND2x1p5_ASAP7_75t_L g1606 ( 
.A(n_1387),
.B(n_1388),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1475),
.B(n_1479),
.Y(n_1607)
);

AO22x1_ASAP7_75t_L g1608 ( 
.A1(n_1492),
.A2(n_1254),
.B1(n_1294),
.B2(n_1235),
.Y(n_1608)
);

INVx6_ASAP7_75t_L g1609 ( 
.A(n_1168),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1107),
.A2(n_1153),
.B1(n_1073),
.B2(n_1214),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1167),
.B(n_1176),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1088),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1513),
.B(n_1511),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1489),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1176),
.B(n_1178),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1482),
.A2(n_1491),
.B1(n_1495),
.B2(n_1493),
.C(n_1487),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1498),
.B(n_1502),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1178),
.B(n_1182),
.Y(n_1618)
);

AND2x6_ASAP7_75t_SL g1619 ( 
.A(n_1460),
.B(n_1465),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1504),
.B(n_1510),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1247),
.A2(n_1517),
.B1(n_1521),
.B2(n_1515),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1371),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1518),
.B(n_1179),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1088),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1098),
.B(n_1035),
.Y(n_1625)
);

OAI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1308),
.A2(n_1246),
.B1(n_1126),
.B2(n_1260),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1182),
.B(n_1194),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1356),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1356),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1466),
.A2(n_1505),
.B1(n_1512),
.B2(n_1476),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1092),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1107),
.A2(n_1153),
.B1(n_1220),
.B2(n_1253),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1204),
.B(n_1050),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1194),
.B(n_1205),
.Y(n_1634)
);

NAND2x1p5_ASAP7_75t_L g1635 ( 
.A(n_1389),
.B(n_1093),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1282),
.B(n_1171),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1205),
.B(n_1208),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1115),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1208),
.B(n_1231),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1231),
.B(n_1233),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1233),
.B(n_1243),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1243),
.B(n_1245),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1092),
.B(n_1112),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1112),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1153),
.A2(n_1045),
.B1(n_1225),
.B2(n_1201),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1232),
.A2(n_1236),
.B1(n_1296),
.B2(n_1289),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1123),
.B(n_1131),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1444),
.B(n_1469),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1123),
.B(n_1131),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1245),
.B(n_1248),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1138),
.B(n_1141),
.Y(n_1651)
);

AO22x1_ASAP7_75t_L g1652 ( 
.A1(n_1294),
.A2(n_1235),
.B1(n_1270),
.B2(n_1217),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1473),
.B(n_1079),
.Y(n_1653)
);

AOI22x1_ASAP7_75t_L g1654 ( 
.A1(n_1311),
.A2(n_1332),
.B1(n_1346),
.B2(n_1331),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1151),
.A2(n_1258),
.B(n_1239),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1115),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1115),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1248),
.B(n_1250),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1250),
.B(n_1266),
.Y(n_1659)
);

NOR3xp33_ASAP7_75t_L g1660 ( 
.A(n_1052),
.B(n_1039),
.C(n_1448),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1044),
.A2(n_1038),
.B1(n_1040),
.B2(n_1101),
.Y(n_1661)
);

AND2x6_ASAP7_75t_L g1662 ( 
.A(n_1395),
.B(n_1345),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_SL g1663 ( 
.A1(n_1116),
.A2(n_1159),
.B1(n_1446),
.B2(n_1120),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1489),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1138),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1141),
.B(n_1143),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1252),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1170),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1062),
.B(n_1066),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1158),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1423),
.B(n_1051),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1473),
.B(n_1079),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1117),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1266),
.B(n_1268),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1075),
.A2(n_1193),
.B1(n_1286),
.B2(n_1104),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1143),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1117),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1268),
.B(n_1289),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1431),
.B(n_1432),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1454),
.A2(n_1461),
.B(n_1471),
.C(n_1457),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1431),
.B(n_1432),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1117),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1439),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1051),
.B(n_1070),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1170),
.Y(n_1685)
);

INVx4_ASAP7_75t_L g1686 ( 
.A(n_1116),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1439),
.B(n_1442),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1051),
.A2(n_1433),
.B1(n_1459),
.B2(n_1070),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1442),
.B(n_1451),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1451),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1477),
.B(n_1485),
.Y(n_1691)
);

INVx8_ASAP7_75t_L g1692 ( 
.A(n_1116),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1488),
.B(n_1497),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1488),
.B(n_1497),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1477),
.B(n_1485),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1490),
.B(n_1503),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1490),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1353),
.B(n_1445),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_SL g1699 ( 
.A1(n_1256),
.A2(n_1262),
.B(n_1173),
.C(n_1259),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1127),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1503),
.B(n_1509),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1353),
.B(n_1445),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1216),
.B(n_1303),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1353),
.B(n_1445),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1230),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1051),
.A2(n_1433),
.B1(n_1459),
.B2(n_1070),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1509),
.B(n_1519),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1519),
.B(n_1520),
.Y(n_1708)
);

BUFx12f_ASAP7_75t_L g1709 ( 
.A(n_1230),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1070),
.A2(n_1433),
.B1(n_1481),
.B2(n_1459),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1171),
.B(n_1064),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1520),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1171),
.B(n_1064),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1177),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1316),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1252),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1064),
.B(n_1433),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1337),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1447),
.B(n_1456),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_SL g1720 ( 
.A(n_1287),
.B(n_1508),
.C(n_1499),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1217),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1316),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1459),
.A2(n_1481),
.B1(n_1219),
.B2(n_1264),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1041),
.A2(n_1251),
.B1(n_1212),
.B2(n_1210),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1171),
.B(n_1064),
.Y(n_1725)
);

OAI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1219),
.A2(n_1174),
.B1(n_1463),
.B2(n_1047),
.C(n_1228),
.Y(n_1726)
);

AND2x6_ASAP7_75t_L g1727 ( 
.A(n_1395),
.B(n_1389),
.Y(n_1727)
);

OAI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1126),
.A2(n_1120),
.B1(n_1159),
.B2(n_1116),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1328),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1127),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1328),
.Y(n_1731)
);

OR2x6_ASAP7_75t_L g1732 ( 
.A(n_1216),
.B(n_1303),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1158),
.B(n_1483),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1300),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1481),
.A2(n_1309),
.B1(n_1288),
.B2(n_1290),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1216),
.B(n_1303),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1481),
.B(n_1235),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1300),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1283),
.A2(n_1292),
.B1(n_1237),
.B2(n_1216),
.Y(n_1739)
);

NAND2x1p5_ASAP7_75t_L g1740 ( 
.A(n_1093),
.B(n_1168),
.Y(n_1740)
);

INVx2_ASAP7_75t_SL g1741 ( 
.A(n_1337),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1304),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1297),
.Y(n_1743)
);

NOR2x1p5_ASAP7_75t_L g1744 ( 
.A(n_1048),
.B(n_1516),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1304),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1216),
.A2(n_1303),
.B1(n_1094),
.B2(n_1212),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1337),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1127),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1235),
.B(n_1421),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1235),
.B(n_1421),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1048),
.B(n_1516),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1132),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1132),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1235),
.B(n_1472),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1353),
.B(n_1445),
.Y(n_1755)
);

AND2x2_ASAP7_75t_SL g1756 ( 
.A(n_1412),
.B(n_1413),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1095),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1095),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1158),
.Y(n_1759)
);

NAND3xp33_ASAP7_75t_SL g1760 ( 
.A(n_1103),
.B(n_1078),
.C(n_1077),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1158),
.B(n_1483),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1235),
.B(n_1472),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1303),
.A2(n_1210),
.B1(n_1516),
.B2(n_1048),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1483),
.B(n_1168),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1472),
.B(n_1436),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1132),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1472),
.B(n_1329),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1087),
.A2(n_1126),
.B1(n_1199),
.B2(n_1353),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1126),
.A2(n_1353),
.B1(n_1445),
.B2(n_1217),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1445),
.B(n_1275),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1336),
.B(n_1331),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1445),
.B(n_1280),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_SL g1773 ( 
.A1(n_1116),
.A2(n_1159),
.B1(n_1446),
.B2(n_1120),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1126),
.A2(n_1445),
.B1(n_1217),
.B2(n_1238),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1136),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1168),
.B(n_1483),
.Y(n_1776)
);

NAND2x1p5_ASAP7_75t_L g1777 ( 
.A(n_1169),
.B(n_1244),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1331),
.B(n_1346),
.Y(n_1778)
);

O2A1O1Ixp5_ASAP7_75t_L g1779 ( 
.A1(n_1344),
.A2(n_1398),
.B(n_1376),
.C(n_1375),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1170),
.Y(n_1780)
);

CKINVDCx6p67_ASAP7_75t_R g1781 ( 
.A(n_1058),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1346),
.B(n_1362),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1362),
.B(n_1522),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1372),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1175),
.B(n_1333),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1362),
.B(n_1522),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1522),
.B(n_1136),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1095),
.Y(n_1788)
);

NAND2xp33_ASAP7_75t_L g1789 ( 
.A(n_1311),
.B(n_1332),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1136),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1224),
.A2(n_1277),
.B1(n_1053),
.B2(n_1065),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1436),
.B(n_1455),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1140),
.B(n_1144),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1140),
.B(n_1144),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1140),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1144),
.B(n_1145),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1145),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1455),
.B(n_1468),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1145),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1147),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1468),
.A2(n_1514),
.B1(n_1285),
.B2(n_1241),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1295),
.A2(n_1365),
.B(n_1110),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1147),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1147),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1514),
.B(n_1057),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1155),
.B(n_1506),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1155),
.B(n_1506),
.Y(n_1807)
);

NOR3xp33_ASAP7_75t_L g1808 ( 
.A(n_1082),
.B(n_1089),
.C(n_1086),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1155),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1318),
.B(n_1322),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1120),
.A2(n_1159),
.B1(n_1501),
.B2(n_1446),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1467),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1129),
.B(n_1130),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1206),
.B(n_1302),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1165),
.B(n_1166),
.Y(n_1815)
);

OR2x2_ASAP7_75t_SL g1816 ( 
.A(n_1397),
.B(n_1081),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1166),
.B(n_1187),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1187),
.B(n_1189),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1187),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1189),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1189),
.B(n_1192),
.Y(n_1821)
);

AND2x2_ASAP7_75t_SL g1822 ( 
.A(n_1351),
.B(n_1361),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1049),
.B(n_1113),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1192),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1192),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1195),
.B(n_1222),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1378),
.B(n_1382),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1056),
.A2(n_1424),
.B1(n_1494),
.B2(n_1480),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1206),
.B(n_1161),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1195),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1222),
.Y(n_1831)
);

NOR3xp33_ASAP7_75t_L g1832 ( 
.A(n_1090),
.B(n_1099),
.C(n_1096),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1255),
.Y(n_1833)
);

INVx4_ASAP7_75t_L g1834 ( 
.A(n_1120),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1351),
.B(n_1361),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1467),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1255),
.B(n_1278),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1114),
.B(n_1118),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1119),
.A2(n_1242),
.B(n_1249),
.C(n_1181),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1161),
.B(n_1180),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1281),
.A2(n_1215),
.B1(n_1446),
.B2(n_1159),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1378),
.B(n_1382),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1279),
.B(n_1299),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1279),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1056),
.A2(n_1430),
.B1(n_1480),
.B2(n_1091),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1299),
.Y(n_1847)
);

OAI22x1_ASAP7_75t_SL g1848 ( 
.A1(n_1325),
.A2(n_1109),
.B1(n_1484),
.B2(n_1058),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1299),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1063),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1063),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1076),
.B(n_1223),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1417),
.B(n_1386),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1076),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1427),
.B(n_1430),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1427),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1058),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1446),
.A2(n_1501),
.B1(n_1109),
.B2(n_1263),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1438),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1438),
.B(n_1383),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_1467),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1383),
.B(n_1501),
.Y(n_1862)
);

AND2x4_ASAP7_75t_SL g1863 ( 
.A(n_1351),
.B(n_1361),
.Y(n_1863)
);

AOI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1501),
.A2(n_1265),
.B1(n_1261),
.B2(n_1059),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1501),
.B(n_1334),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1307),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1291),
.B(n_1170),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1334),
.B(n_1341),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1341),
.B(n_1342),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1170),
.B(n_1226),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1081),
.Y(n_1871)
);

A2O1A1Ixp33_ASAP7_75t_L g1872 ( 
.A1(n_1271),
.A2(n_1313),
.B(n_1055),
.C(n_1408),
.Y(n_1872)
);

INVx3_ASAP7_75t_L g1873 ( 
.A(n_1226),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1342),
.B(n_1352),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1226),
.B(n_1317),
.Y(n_1875)
);

BUFx2_ASAP7_75t_L g1876 ( 
.A(n_1372),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1312),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1352),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1354),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1354),
.B(n_1359),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1359),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1363),
.B(n_1366),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1054),
.B(n_1363),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1372),
.B(n_1393),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_1381),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1366),
.B(n_1384),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1226),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1393),
.Y(n_1888)
);

OAI221xp5_ASAP7_75t_L g1889 ( 
.A1(n_1240),
.A2(n_1355),
.B1(n_1325),
.B2(n_1364),
.C(n_1349),
.Y(n_1889)
);

AND2x6_ASAP7_75t_SL g1890 ( 
.A(n_1133),
.B(n_1156),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1377),
.A2(n_1306),
.B1(n_1484),
.B2(n_1133),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1226),
.B(n_1317),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1339),
.B(n_1343),
.Y(n_1893)
);

AO22x1_ASAP7_75t_L g1894 ( 
.A1(n_1405),
.A2(n_1420),
.B1(n_1351),
.B2(n_1361),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1350),
.B(n_1357),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1394),
.B(n_1374),
.Y(n_1896)
);

BUFx4f_ASAP7_75t_L g1897 ( 
.A(n_1422),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1393),
.Y(n_1898)
);

INVx2_ASAP7_75t_SL g1899 ( 
.A(n_1317),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1133),
.A2(n_1484),
.B1(n_1156),
.B2(n_1411),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1156),
.A2(n_1197),
.B1(n_1191),
.B2(n_1180),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1420),
.A2(n_1326),
.B1(n_1324),
.B2(n_1191),
.Y(n_1902)
);

BUFx4f_ASAP7_75t_L g1903 ( 
.A(n_1422),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1319),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1374),
.B(n_1367),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1374),
.B(n_1370),
.Y(n_1906)
);

INVx4_ASAP7_75t_L g1907 ( 
.A(n_1422),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1370),
.B(n_1407),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1197),
.A2(n_1081),
.B1(n_1321),
.B2(n_1293),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1404),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1385),
.A2(n_1335),
.B1(n_1330),
.B2(n_1373),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1370),
.B(n_1404),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1404),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1407),
.B(n_1396),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1370),
.B(n_1407),
.Y(n_1915)
);

NAND3xp33_ASAP7_75t_SL g1916 ( 
.A(n_1409),
.B(n_1403),
.C(n_1401),
.Y(n_1916)
);

OAI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1402),
.A2(n_1379),
.B1(n_1380),
.B2(n_1301),
.C(n_1284),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1081),
.A2(n_1323),
.B1(n_1320),
.B2(n_1314),
.Y(n_1918)
);

NAND2xp33_ASAP7_75t_L g1919 ( 
.A(n_1317),
.B(n_1373),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1267),
.A2(n_1298),
.B1(n_1276),
.B2(n_1340),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1317),
.B(n_1425),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1373),
.B(n_1425),
.Y(n_1922)
);

INVx5_ASAP7_75t_L g1923 ( 
.A(n_1422),
.Y(n_1923)
);

OAI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1410),
.A2(n_1188),
.B1(n_1422),
.B2(n_1068),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1373),
.Y(n_1925)
);

INVxp33_ASAP7_75t_L g1926 ( 
.A(n_1169),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1360),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_SL g1928 ( 
.A(n_1360),
.B(n_1244),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1373),
.A2(n_1425),
.B1(n_1068),
.B2(n_1406),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1390),
.A2(n_1391),
.B(n_1400),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_SL g1931 ( 
.A(n_1188),
.B(n_1419),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1425),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1358),
.A2(n_1369),
.B(n_1425),
.Y(n_1933)
);

OAI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1410),
.A2(n_1419),
.B(n_1414),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1416),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1368),
.Y(n_1936)
);

INVx3_ASAP7_75t_L g1937 ( 
.A(n_1392),
.Y(n_1937)
);

NAND2x1p5_ASAP7_75t_L g1938 ( 
.A(n_1348),
.B(n_1387),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1142),
.B(n_739),
.Y(n_1940)
);

AND3x1_ASAP7_75t_L g1941 ( 
.A(n_1042),
.B(n_1142),
.C(n_1164),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1121),
.B(n_1135),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1368),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1142),
.B(n_739),
.Y(n_1944)
);

INVx1_ASAP7_75t_SL g1945 ( 
.A(n_1518),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1368),
.Y(n_1946)
);

HB1xp67_ASAP7_75t_L g1947 ( 
.A(n_1135),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1368),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1368),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1348),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1142),
.B(n_739),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1954)
);

BUFx12f_ASAP7_75t_L g1955 ( 
.A(n_1230),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1142),
.A2(n_1209),
.B1(n_1084),
.B2(n_868),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1196),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1043),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1043),
.Y(n_1960)
);

AND2x6_ASAP7_75t_SL g1961 ( 
.A(n_1164),
.B(n_1163),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1142),
.B(n_739),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1121),
.B(n_1085),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1043),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1348),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1142),
.B(n_1209),
.Y(n_1970)
);

AOI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_SL g1972 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1142),
.B(n_1209),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1043),
.Y(n_1974)
);

AOI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1142),
.A2(n_1042),
.B1(n_519),
.B2(n_1209),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1142),
.B(n_1209),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1142),
.A2(n_1209),
.B1(n_1084),
.B2(n_868),
.Y(n_1978)
);

AO22x1_ASAP7_75t_L g1979 ( 
.A1(n_1042),
.A2(n_810),
.B1(n_1415),
.B2(n_822),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1142),
.A2(n_1042),
.B1(n_519),
.B2(n_1209),
.Y(n_1980)
);

NAND3xp33_ASAP7_75t_L g1981 ( 
.A(n_1042),
.B(n_1142),
.C(n_1257),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1982)
);

INVx8_ASAP7_75t_L g1983 ( 
.A(n_1116),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1368),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1142),
.B(n_1209),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1043),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1368),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1142),
.B(n_1209),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1043),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1172),
.Y(n_1993)
);

INVx2_ASAP7_75t_SL g1994 ( 
.A(n_1196),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1043),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1043),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1998)
);

NOR2xp67_ASAP7_75t_L g1999 ( 
.A(n_1370),
.B(n_1397),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1368),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1142),
.B(n_739),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1043),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1121),
.B(n_1085),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_L g2006 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1368),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2008)
);

AO22x1_ASAP7_75t_L g2009 ( 
.A1(n_1042),
.A2(n_810),
.B1(n_1415),
.B2(n_822),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1043),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1348),
.Y(n_2011)
);

AOI22xp5_ASAP7_75t_L g2012 ( 
.A1(n_1142),
.A2(n_1042),
.B1(n_519),
.B2(n_1209),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1043),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1142),
.B(n_739),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1142),
.B(n_739),
.Y(n_2015)
);

AND2x4_ASAP7_75t_L g2016 ( 
.A(n_1315),
.B(n_1061),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1142),
.B(n_739),
.Y(n_2018)
);

BUFx3_ASAP7_75t_L g2019 ( 
.A(n_1061),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2022)
);

A2O1A1Ixp33_ASAP7_75t_L g2023 ( 
.A1(n_1142),
.A2(n_1209),
.B(n_1042),
.C(n_1257),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1043),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1368),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2035)
);

INVxp67_ASAP7_75t_L g2036 ( 
.A(n_1079),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_SL g2039 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2039)
);

NOR2x2_ASAP7_75t_L g2040 ( 
.A(n_1200),
.B(n_368),
.Y(n_2040)
);

OR2x6_ASAP7_75t_L g2041 ( 
.A(n_1392),
.B(n_1216),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1043),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1142),
.A2(n_1209),
.B1(n_1084),
.B2(n_868),
.Y(n_2043)
);

INVx2_ASAP7_75t_SL g2044 ( 
.A(n_1196),
.Y(n_2044)
);

AO22x1_ASAP7_75t_L g2045 ( 
.A1(n_1042),
.A2(n_810),
.B1(n_1415),
.B2(n_822),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1368),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2047)
);

AND2x6_ASAP7_75t_SL g2048 ( 
.A(n_1164),
.B(n_1163),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1142),
.A2(n_1042),
.B1(n_519),
.B2(n_1209),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2050)
);

NAND3xp33_ASAP7_75t_SL g2051 ( 
.A(n_1142),
.B(n_1042),
.C(n_1209),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1043),
.Y(n_2053)
);

INVx8_ASAP7_75t_L g2054 ( 
.A(n_1116),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1142),
.B(n_739),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1368),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_SL g2057 ( 
.A(n_1348),
.B(n_1116),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1043),
.Y(n_2058)
);

AND2x6_ASAP7_75t_L g2059 ( 
.A(n_1415),
.B(n_1327),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1348),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1142),
.B(n_739),
.Y(n_2062)
);

NOR3xp33_ASAP7_75t_L g2063 ( 
.A(n_1042),
.B(n_1441),
.C(n_1108),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1368),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1368),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2070)
);

NAND2x1p5_ASAP7_75t_L g2071 ( 
.A(n_1348),
.B(n_1387),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1142),
.B(n_739),
.Y(n_2073)
);

O2A1O1Ixp33_ASAP7_75t_L g2074 ( 
.A1(n_1042),
.A2(n_913),
.B(n_906),
.C(n_923),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_L g2075 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1142),
.B(n_739),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1142),
.B(n_739),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1043),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1368),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1142),
.B(n_739),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2083)
);

INVx8_ASAP7_75t_L g2084 ( 
.A(n_1116),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1043),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1043),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1043),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1121),
.B(n_1135),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1043),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2090)
);

BUFx3_ASAP7_75t_L g2091 ( 
.A(n_1061),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2092)
);

AOI22xp33_ASAP7_75t_L g2093 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2093)
);

AOI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_1142),
.A2(n_1042),
.B1(n_519),
.B2(n_1209),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1368),
.Y(n_2095)
);

NAND2x1p5_ASAP7_75t_L g2096 ( 
.A(n_1348),
.B(n_1387),
.Y(n_2096)
);

AOI21xp33_ASAP7_75t_L g2097 ( 
.A1(n_1418),
.A2(n_1142),
.B(n_1209),
.Y(n_2097)
);

AOI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2098)
);

NOR2x2_ASAP7_75t_L g2099 ( 
.A(n_1200),
.B(n_368),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1043),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1142),
.B(n_739),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_1061),
.Y(n_2102)
);

HB1xp67_ASAP7_75t_L g2103 ( 
.A(n_1135),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1043),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_1142),
.B(n_739),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_1142),
.B(n_739),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_1348),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1142),
.B(n_739),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1368),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_L g2113 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_1135),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1043),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_1142),
.B(n_739),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2120)
);

INVx5_ASAP7_75t_L g2121 ( 
.A(n_1392),
.Y(n_2121)
);

NAND2x1p5_ASAP7_75t_L g2122 ( 
.A(n_1348),
.B(n_1387),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1043),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1368),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_1142),
.B(n_739),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1368),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1142),
.B(n_739),
.Y(n_2131)
);

INVxp67_ASAP7_75t_L g2132 ( 
.A(n_1079),
.Y(n_2132)
);

BUFx3_ASAP7_75t_L g2133 ( 
.A(n_1061),
.Y(n_2133)
);

AOI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_1142),
.A2(n_1042),
.B1(n_519),
.B2(n_1209),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2135)
);

NAND3xp33_ASAP7_75t_L g2136 ( 
.A(n_1042),
.B(n_1142),
.C(n_1257),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2137)
);

OAI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1142),
.A2(n_1209),
.B1(n_1084),
.B2(n_868),
.Y(n_2138)
);

HB1xp67_ASAP7_75t_L g2139 ( 
.A(n_1135),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1043),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1142),
.B(n_739),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1172),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1043),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_1142),
.B(n_739),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2146)
);

INVx2_ASAP7_75t_SL g2147 ( 
.A(n_1196),
.Y(n_2147)
);

AOI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_1142),
.A2(n_1042),
.B1(n_519),
.B2(n_1209),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1368),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2153)
);

INVx1_ASAP7_75t_SL g2154 ( 
.A(n_1518),
.Y(n_2154)
);

OAI22xp5_ASAP7_75t_L g2155 ( 
.A1(n_1142),
.A2(n_1209),
.B1(n_1084),
.B2(n_868),
.Y(n_2155)
);

CKINVDCx11_ASAP7_75t_R g2156 ( 
.A(n_1177),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1043),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_1142),
.B(n_739),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1043),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_SL g2163 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_1142),
.A2(n_1042),
.B1(n_519),
.B2(n_1209),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1368),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_1142),
.B(n_739),
.Y(n_2168)
);

AOI22xp33_ASAP7_75t_L g2169 ( 
.A1(n_1418),
.A2(n_382),
.B1(n_490),
.B2(n_485),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2170)
);

O2A1O1Ixp33_ASAP7_75t_L g2171 ( 
.A1(n_1042),
.A2(n_913),
.B(n_906),
.C(n_923),
.Y(n_2171)
);

AND2x6_ASAP7_75t_SL g2172 ( 
.A(n_1164),
.B(n_1163),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1043),
.Y(n_2173)
);

INVx5_ASAP7_75t_L g2174 ( 
.A(n_1392),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1368),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1085),
.B(n_1135),
.Y(n_2178)
);

OAI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_1142),
.A2(n_1209),
.B1(n_1084),
.B2(n_868),
.Y(n_2179)
);

AND2x4_ASAP7_75t_L g2180 ( 
.A(n_1315),
.B(n_1061),
.Y(n_2180)
);

NOR2xp67_ASAP7_75t_L g2181 ( 
.A(n_1370),
.B(n_1397),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1142),
.B(n_1209),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1368),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1526),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_1942),
.B(n_2088),
.Y(n_2186)
);

HB1xp67_ASAP7_75t_L g2187 ( 
.A(n_1556),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1557),
.B(n_1563),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1557),
.B(n_1563),
.Y(n_2189)
);

OR2x6_ASAP7_75t_L g2190 ( 
.A(n_1732),
.B(n_2041),
.Y(n_2190)
);

NOR3xp33_ASAP7_75t_SL g2191 ( 
.A(n_1993),
.B(n_2143),
.C(n_1705),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_1668),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1568),
.B(n_1576),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_2041),
.B(n_1555),
.Y(n_2194)
);

BUFx6f_ASAP7_75t_L g2195 ( 
.A(n_1668),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_1941),
.B(n_1528),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1942),
.B(n_2088),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_1947),
.B(n_2103),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1628),
.Y(n_2199)
);

INVx5_ASAP7_75t_L g2200 ( 
.A(n_2041),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1526),
.Y(n_2201)
);

INVxp67_ASAP7_75t_L g2202 ( 
.A(n_1693),
.Y(n_2202)
);

BUFx2_ASAP7_75t_L g2203 ( 
.A(n_1556),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1526),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_2041),
.B(n_1555),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1942),
.B(n_2088),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1568),
.B(n_1576),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1571),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1628),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_2041),
.B(n_1555),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_1534),
.B(n_1604),
.Y(n_2211)
);

BUFx3_ASAP7_75t_L g2212 ( 
.A(n_1816),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_1940),
.A2(n_1962),
.B1(n_2003),
.B2(n_1953),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_1941),
.B(n_1528),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_1981),
.B(n_2136),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_1534),
.B(n_1604),
.Y(n_2216)
);

NOR2xp67_ASAP7_75t_L g2217 ( 
.A(n_1556),
.B(n_1573),
.Y(n_2217)
);

BUFx2_ASAP7_75t_L g2218 ( 
.A(n_1573),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1571),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_SL g2220 ( 
.A(n_1981),
.B(n_2136),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_L g2221 ( 
.A1(n_1972),
.A2(n_2039),
.B1(n_1971),
.B2(n_1976),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1628),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1629),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1571),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1586),
.B(n_1592),
.Y(n_2225)
);

AND3x1_ASAP7_75t_SL g2226 ( 
.A(n_1616),
.B(n_1619),
.C(n_1630),
.Y(n_2226)
);

NAND2x1p5_ASAP7_75t_L g2227 ( 
.A(n_1698),
.B(n_1702),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1574),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1574),
.Y(n_2229)
);

OAI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_1551),
.A2(n_2148),
.B1(n_2164),
.B2(n_2012),
.Y(n_2230)
);

BUFx2_ASAP7_75t_SL g2231 ( 
.A(n_1573),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1586),
.B(n_1592),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_1940),
.B(n_1953),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1629),
.Y(n_2234)
);

BUFx3_ASAP7_75t_L g2235 ( 
.A(n_1816),
.Y(n_2235)
);

BUFx6f_ASAP7_75t_L g2236 ( 
.A(n_1668),
.Y(n_2236)
);

INVx3_ASAP7_75t_SL g2237 ( 
.A(n_1562),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_1958),
.Y(n_2238)
);

BUFx6f_ASAP7_75t_L g2239 ( 
.A(n_1668),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1544),
.B(n_1549),
.Y(n_2240)
);

BUFx2_ASAP7_75t_L g2241 ( 
.A(n_1958),
.Y(n_2241)
);

NOR2x1p5_ASAP7_75t_L g2242 ( 
.A(n_1781),
.B(n_2051),
.Y(n_2242)
);

OAI22xp5_ASAP7_75t_SL g2243 ( 
.A1(n_1630),
.A2(n_1975),
.B1(n_2012),
.B2(n_1980),
.Y(n_2243)
);

BUFx6f_ASAP7_75t_L g2244 ( 
.A(n_1668),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_1534),
.B(n_1604),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_1572),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_L g2247 ( 
.A(n_1962),
.B(n_2003),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1629),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_2014),
.B(n_2015),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1574),
.Y(n_2250)
);

NOR3xp33_ASAP7_75t_SL g2251 ( 
.A(n_1616),
.B(n_1720),
.C(n_1614),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_1668),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1591),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1591),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1544),
.B(n_1549),
.Y(n_2255)
);

HB1xp67_ASAP7_75t_L g2256 ( 
.A(n_1958),
.Y(n_2256)
);

INVx2_ASAP7_75t_SL g2257 ( 
.A(n_1994),
.Y(n_2257)
);

BUFx2_ASAP7_75t_L g2258 ( 
.A(n_1994),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1591),
.Y(n_2259)
);

INVxp67_ASAP7_75t_SL g2260 ( 
.A(n_1531),
.Y(n_2260)
);

BUFx6f_ASAP7_75t_SL g2261 ( 
.A(n_1952),
.Y(n_2261)
);

BUFx3_ASAP7_75t_L g2262 ( 
.A(n_1816),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2014),
.B(n_2015),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1605),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1605),
.Y(n_2265)
);

INVx2_ASAP7_75t_SL g2266 ( 
.A(n_1994),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_1537),
.B(n_1947),
.Y(n_2267)
);

BUFx6f_ASAP7_75t_L g2268 ( 
.A(n_1685),
.Y(n_2268)
);

BUFx6f_ASAP7_75t_L g2269 ( 
.A(n_1685),
.Y(n_2269)
);

BUFx2_ASAP7_75t_L g2270 ( 
.A(n_2044),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1537),
.B(n_2103),
.Y(n_2271)
);

BUFx2_ASAP7_75t_L g2272 ( 
.A(n_2044),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1605),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1622),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2041),
.B(n_1555),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_1555),
.B(n_1583),
.Y(n_2276)
);

NOR3xp33_ASAP7_75t_SL g2277 ( 
.A(n_1720),
.B(n_1664),
.C(n_1602),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1622),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_1904),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_2156),
.Y(n_2280)
);

BUFx4f_ASAP7_75t_L g2281 ( 
.A(n_1777),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2115),
.B(n_2139),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1622),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_2018),
.B(n_2055),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1936),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1936),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_2018),
.B(n_2055),
.Y(n_2287)
);

BUFx12f_ASAP7_75t_L g2288 ( 
.A(n_1890),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_1555),
.B(n_1583),
.Y(n_2289)
);

AND2x4_ASAP7_75t_L g2290 ( 
.A(n_1555),
.B(n_1583),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_2108),
.B(n_2128),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2115),
.B(n_2139),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1533),
.B(n_1531),
.Y(n_2293)
);

NOR3xp33_ASAP7_75t_SL g2294 ( 
.A(n_2051),
.B(n_1714),
.C(n_1648),
.Y(n_2294)
);

OAI22xp33_ASAP7_75t_L g2295 ( 
.A1(n_1551),
.A2(n_1980),
.B1(n_2094),
.B2(n_1975),
.Y(n_2295)
);

INVx4_ASAP7_75t_L g2296 ( 
.A(n_1555),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1936),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1533),
.B(n_1595),
.Y(n_2298)
);

INVx1_ASAP7_75t_SL g2299 ( 
.A(n_1577),
.Y(n_2299)
);

NAND3xp33_ASAP7_75t_SL g2300 ( 
.A(n_2049),
.B(n_2134),
.C(n_2094),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1943),
.Y(n_2301)
);

A2O1A1Ixp33_ASAP7_75t_L g2302 ( 
.A1(n_2108),
.A2(n_2128),
.B(n_2160),
.C(n_2145),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1943),
.Y(n_2303)
);

CKINVDCx20_ASAP7_75t_R g2304 ( 
.A(n_1547),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_1943),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1946),
.Y(n_2306)
);

HB1xp67_ASAP7_75t_L g2307 ( 
.A(n_2044),
.Y(n_2307)
);

INVxp67_ASAP7_75t_L g2308 ( 
.A(n_1693),
.Y(n_2308)
);

CKINVDCx20_ASAP7_75t_R g2309 ( 
.A(n_1547),
.Y(n_2309)
);

AND2x6_ASAP7_75t_L g2310 ( 
.A(n_1952),
.B(n_1969),
.Y(n_2310)
);

OR2x6_ASAP7_75t_L g2311 ( 
.A(n_1732),
.B(n_1524),
.Y(n_2311)
);

INVx4_ASAP7_75t_L g2312 ( 
.A(n_1583),
.Y(n_2312)
);

AOI22xp5_ASAP7_75t_L g2313 ( 
.A1(n_2145),
.A2(n_2168),
.B1(n_2160),
.B2(n_1970),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_1946),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2168),
.B(n_2049),
.Y(n_2315)
);

A2O1A1Ixp33_ASAP7_75t_L g2316 ( 
.A1(n_2023),
.A2(n_1970),
.B(n_1973),
.C(n_1524),
.Y(n_2316)
);

AND2x4_ASAP7_75t_L g2317 ( 
.A(n_1583),
.B(n_2121),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1946),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_1580),
.B(n_1538),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1533),
.B(n_1595),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_1583),
.B(n_2121),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1594),
.B(n_1643),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_1949),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1949),
.Y(n_2324)
);

OR2x2_ASAP7_75t_L g2325 ( 
.A(n_1973),
.B(n_1977),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_2134),
.B(n_2148),
.Y(n_2326)
);

AOI22xp33_ASAP7_75t_L g2327 ( 
.A1(n_1972),
.A2(n_2039),
.B1(n_1967),
.B2(n_1976),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_1949),
.Y(n_2328)
);

INVx4_ASAP7_75t_L g2329 ( 
.A(n_1583),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1951),
.Y(n_2330)
);

INVx2_ASAP7_75t_SL g2331 ( 
.A(n_2147),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_1594),
.B(n_1643),
.Y(n_2332)
);

HB1xp67_ASAP7_75t_L g2333 ( 
.A(n_2147),
.Y(n_2333)
);

INVx5_ASAP7_75t_L g2334 ( 
.A(n_1952),
.Y(n_2334)
);

NOR3xp33_ASAP7_75t_SL g2335 ( 
.A(n_1584),
.B(n_2171),
.C(n_2074),
.Y(n_2335)
);

OAI21xp5_ASAP7_75t_L g2336 ( 
.A1(n_1977),
.A2(n_2182),
.B(n_1991),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_1685),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_2164),
.B(n_1619),
.Y(n_2338)
);

BUFx2_ASAP7_75t_L g2339 ( 
.A(n_2147),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_1583),
.B(n_2121),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_1709),
.Y(n_2341)
);

OR2x6_ASAP7_75t_SL g2342 ( 
.A(n_1956),
.B(n_1978),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_1580),
.B(n_1538),
.Y(n_2343)
);

CKINVDCx5p33_ASAP7_75t_R g2344 ( 
.A(n_1709),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1643),
.B(n_1647),
.Y(n_2345)
);

AND2x2_ASAP7_75t_SL g2346 ( 
.A(n_1610),
.B(n_1543),
.Y(n_2346)
);

HB1xp67_ASAP7_75t_L g2347 ( 
.A(n_1910),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_1647),
.B(n_1649),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_1621),
.B(n_1539),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1984),
.Y(n_2350)
);

OR2x6_ASAP7_75t_L g2351 ( 
.A(n_1732),
.B(n_1985),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1984),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1989),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1647),
.B(n_1649),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_1649),
.B(n_1651),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_1989),
.Y(n_2356)
);

INVx4_ASAP7_75t_L g2357 ( 
.A(n_2121),
.Y(n_2357)
);

INVx8_ASAP7_75t_L g2358 ( 
.A(n_1692),
.Y(n_2358)
);

AND2x4_ASAP7_75t_L g2359 ( 
.A(n_2121),
.B(n_2174),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1989),
.Y(n_2360)
);

BUFx6f_ASAP7_75t_L g2361 ( 
.A(n_1685),
.Y(n_2361)
);

BUFx8_ASAP7_75t_SL g2362 ( 
.A(n_1709),
.Y(n_2362)
);

AOI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_1985),
.A2(n_2000),
.B1(n_2022),
.B2(n_1991),
.Y(n_2363)
);

INVx5_ASAP7_75t_L g2364 ( 
.A(n_1952),
.Y(n_2364)
);

INVxp67_ASAP7_75t_L g2365 ( 
.A(n_1694),
.Y(n_2365)
);

BUFx10_ASAP7_75t_L g2366 ( 
.A(n_1890),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_1542),
.B(n_1535),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_1651),
.B(n_1666),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_1651),
.B(n_1666),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_SL g2370 ( 
.A(n_1928),
.B(n_2057),
.Y(n_2370)
);

BUFx8_ASAP7_75t_L g2371 ( 
.A(n_1952),
.Y(n_2371)
);

A2O1A1Ixp33_ASAP7_75t_L g2372 ( 
.A1(n_2182),
.A2(n_2183),
.B(n_2022),
.C(n_2024),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_1955),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2002),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_SL g2375 ( 
.A(n_1928),
.B(n_2057),
.Y(n_2375)
);

NOR3xp33_ASAP7_75t_SL g2376 ( 
.A(n_1584),
.B(n_2171),
.C(n_2074),
.Y(n_2376)
);

INVx2_ASAP7_75t_SL g2377 ( 
.A(n_1685),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_R g2378 ( 
.A(n_1721),
.B(n_1822),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_1780),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2002),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_1967),
.A2(n_1971),
.B1(n_2025),
.B2(n_2006),
.Y(n_2381)
);

BUFx6f_ASAP7_75t_L g2382 ( 
.A(n_1780),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2002),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2007),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_1542),
.B(n_1535),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2007),
.Y(n_2386)
);

AND2x6_ASAP7_75t_L g2387 ( 
.A(n_1952),
.B(n_1969),
.Y(n_2387)
);

HB1xp67_ASAP7_75t_L g2388 ( 
.A(n_1910),
.Y(n_2388)
);

BUFx4_ASAP7_75t_SL g2389 ( 
.A(n_1558),
.Y(n_2389)
);

BUFx3_ASAP7_75t_L g2390 ( 
.A(n_1662),
.Y(n_2390)
);

BUFx2_ASAP7_75t_L g2391 ( 
.A(n_1670),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_1666),
.B(n_1527),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_1527),
.B(n_1532),
.Y(n_2393)
);

OAI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2000),
.A2(n_2029),
.B1(n_2033),
.B2(n_2024),
.Y(n_2394)
);

BUFx3_ASAP7_75t_L g2395 ( 
.A(n_1662),
.Y(n_2395)
);

INVx2_ASAP7_75t_SL g2396 ( 
.A(n_1780),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2034),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_1532),
.B(n_1939),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_SL g2399 ( 
.A(n_1621),
.B(n_1529),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2034),
.Y(n_2400)
);

INVx3_ASAP7_75t_L g2401 ( 
.A(n_1780),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2034),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_L g2403 ( 
.A(n_1539),
.B(n_1944),
.Y(n_2403)
);

BUFx3_ASAP7_75t_L g2404 ( 
.A(n_1662),
.Y(n_2404)
);

OR2x6_ASAP7_75t_L g2405 ( 
.A(n_1732),
.B(n_2029),
.Y(n_2405)
);

AO22x1_ASAP7_75t_L g2406 ( 
.A1(n_1662),
.A2(n_2063),
.B1(n_1978),
.B2(n_2043),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2046),
.Y(n_2407)
);

BUFx6f_ASAP7_75t_L g2408 ( 
.A(n_1780),
.Y(n_2408)
);

AOI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2033),
.A2(n_2038),
.B1(n_2163),
.B2(n_2157),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_1939),
.B(n_1948),
.Y(n_2410)
);

AND2x4_ASAP7_75t_L g2411 ( 
.A(n_2121),
.B(n_2174),
.Y(n_2411)
);

INVx8_ASAP7_75t_L g2412 ( 
.A(n_1692),
.Y(n_2412)
);

INVx3_ASAP7_75t_L g2413 ( 
.A(n_1932),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2046),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2056),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_L g2416 ( 
.A(n_1952),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_2121),
.B(n_2174),
.Y(n_2417)
);

INVxp67_ASAP7_75t_L g2418 ( 
.A(n_1694),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2121),
.B(n_2174),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_1948),
.B(n_1950),
.Y(n_2420)
);

NOR2x1p5_ASAP7_75t_L g2421 ( 
.A(n_1781),
.B(n_1737),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2056),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_SL g2423 ( 
.A(n_1529),
.B(n_2038),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_1950),
.B(n_1954),
.Y(n_2424)
);

BUFx2_ASAP7_75t_SL g2425 ( 
.A(n_2174),
.Y(n_2425)
);

INVx1_ASAP7_75t_SL g2426 ( 
.A(n_1577),
.Y(n_2426)
);

HB1xp67_ASAP7_75t_L g2427 ( 
.A(n_1670),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_2174),
.B(n_1732),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_1954),
.B(n_1957),
.Y(n_2429)
);

INVx3_ASAP7_75t_SL g2430 ( 
.A(n_1857),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_1969),
.Y(n_2431)
);

NAND2xp33_ASAP7_75t_L g2432 ( 
.A(n_1777),
.B(n_1552),
.Y(n_2432)
);

OR2x4_ASAP7_75t_L g2433 ( 
.A(n_1760),
.B(n_1963),
.Y(n_2433)
);

BUFx4f_ASAP7_75t_L g2434 ( 
.A(n_1777),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_1969),
.Y(n_2435)
);

BUFx10_ASAP7_75t_L g2436 ( 
.A(n_1805),
.Y(n_2436)
);

NAND2xp33_ASAP7_75t_SL g2437 ( 
.A(n_2175),
.B(n_2176),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_1957),
.B(n_1965),
.Y(n_2438)
);

AND3x1_ASAP7_75t_SL g2439 ( 
.A(n_1552),
.B(n_1550),
.C(n_1961),
.Y(n_2439)
);

NAND3xp33_ASAP7_75t_SL g2440 ( 
.A(n_2063),
.B(n_1536),
.C(n_1553),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2064),
.Y(n_2441)
);

BUFx4f_ASAP7_75t_L g2442 ( 
.A(n_1777),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_SL g2443 ( 
.A(n_2097),
.B(n_1686),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2064),
.Y(n_2444)
);

BUFx4f_ASAP7_75t_L g2445 ( 
.A(n_1969),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_1965),
.B(n_1966),
.Y(n_2446)
);

BUFx3_ASAP7_75t_L g2447 ( 
.A(n_1662),
.Y(n_2447)
);

BUFx6f_ASAP7_75t_L g2448 ( 
.A(n_1969),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_SL g2449 ( 
.A(n_2175),
.B(n_2176),
.Y(n_2449)
);

BUFx2_ASAP7_75t_L g2450 ( 
.A(n_1759),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_1580),
.B(n_1538),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2064),
.Y(n_2452)
);

OAI22xp5_ASAP7_75t_L g2453 ( 
.A1(n_2183),
.A2(n_1956),
.B1(n_2138),
.B2(n_2043),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2069),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2069),
.Y(n_2455)
);

BUFx3_ASAP7_75t_L g2456 ( 
.A(n_1662),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_1969),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2079),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_1963),
.B(n_2005),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2079),
.Y(n_2460)
);

BUFx2_ASAP7_75t_L g2461 ( 
.A(n_1759),
.Y(n_2461)
);

BUFx3_ASAP7_75t_L g2462 ( 
.A(n_1662),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2079),
.Y(n_2463)
);

AOI22xp33_ASAP7_75t_L g2464 ( 
.A1(n_2006),
.A2(n_2025),
.B1(n_2047),
.B2(n_2030),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_1955),
.Y(n_2465)
);

BUFx2_ASAP7_75t_L g2466 ( 
.A(n_1590),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_R g2467 ( 
.A(n_1822),
.B(n_1789),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_1966),
.B(n_1968),
.Y(n_2468)
);

INVx2_ASAP7_75t_SL g2469 ( 
.A(n_1609),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_1932),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2095),
.Y(n_2471)
);

OR2x6_ASAP7_75t_L g2472 ( 
.A(n_1732),
.B(n_1703),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2095),
.Y(n_2473)
);

BUFx6f_ASAP7_75t_L g2474 ( 
.A(n_2011),
.Y(n_2474)
);

HB1xp67_ASAP7_75t_L g2475 ( 
.A(n_1784),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_SL g2476 ( 
.A(n_1553),
.B(n_2138),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_1541),
.B(n_1963),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2095),
.Y(n_2478)
);

BUFx8_ASAP7_75t_L g2479 ( 
.A(n_2011),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2112),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_1968),
.B(n_1982),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_1982),
.B(n_1986),
.Y(n_2482)
);

INVx1_ASAP7_75t_SL g2483 ( 
.A(n_1945),
.Y(n_2483)
);

INVxp67_ASAP7_75t_L g2484 ( 
.A(n_1726),
.Y(n_2484)
);

BUFx3_ASAP7_75t_L g2485 ( 
.A(n_1662),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2112),
.Y(n_2486)
);

XNOR2xp5_ASAP7_75t_L g2487 ( 
.A(n_2030),
.B(n_2047),
.Y(n_2487)
);

NOR2xp33_ASAP7_75t_L g2488 ( 
.A(n_2062),
.B(n_2073),
.Y(n_2488)
);

INVx4_ASAP7_75t_L g2489 ( 
.A(n_2174),
.Y(n_2489)
);

BUFx3_ASAP7_75t_L g2490 ( 
.A(n_1662),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2125),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2125),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_R g2493 ( 
.A(n_1822),
.B(n_1547),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_1541),
.B(n_2005),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2125),
.Y(n_2495)
);

INVx1_ASAP7_75t_SL g2496 ( 
.A(n_1945),
.Y(n_2496)
);

BUFx4f_ASAP7_75t_SL g2497 ( 
.A(n_1955),
.Y(n_2497)
);

OR2x6_ASAP7_75t_L g2498 ( 
.A(n_1703),
.B(n_1736),
.Y(n_2498)
);

CKINVDCx5p33_ASAP7_75t_R g2499 ( 
.A(n_1558),
.Y(n_2499)
);

OR2x6_ASAP7_75t_L g2500 ( 
.A(n_1703),
.B(n_1736),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2011),
.Y(n_2501)
);

AND2x4_ASAP7_75t_SL g2502 ( 
.A(n_2011),
.B(n_2060),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_SL g2503 ( 
.A(n_2155),
.B(n_2179),
.Y(n_2503)
);

OR2x6_ASAP7_75t_L g2504 ( 
.A(n_1736),
.B(n_1652),
.Y(n_2504)
);

CKINVDCx20_ASAP7_75t_R g2505 ( 
.A(n_1781),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_1986),
.B(n_1987),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2129),
.Y(n_2507)
);

INVx1_ASAP7_75t_SL g2508 ( 
.A(n_2154),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2129),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_1541),
.B(n_2005),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2129),
.Y(n_2511)
);

BUFx3_ASAP7_75t_L g2512 ( 
.A(n_1662),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_1987),
.B(n_1990),
.Y(n_2513)
);

NOR2xp33_ASAP7_75t_R g2514 ( 
.A(n_1822),
.B(n_2011),
.Y(n_2514)
);

BUFx2_ASAP7_75t_L g2515 ( 
.A(n_1590),
.Y(n_2515)
);

INVx3_ASAP7_75t_L g2516 ( 
.A(n_1932),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2150),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_1961),
.Y(n_2518)
);

INVx1_ASAP7_75t_SL g2519 ( 
.A(n_2154),
.Y(n_2519)
);

BUFx3_ASAP7_75t_L g2520 ( 
.A(n_2059),
.Y(n_2520)
);

CKINVDCx16_ASAP7_75t_R g2521 ( 
.A(n_1661),
.Y(n_2521)
);

HB1xp67_ASAP7_75t_L g2522 ( 
.A(n_1784),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_1990),
.B(n_1995),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2150),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2165),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_1995),
.B(n_1998),
.Y(n_2526)
);

INVx3_ASAP7_75t_L g2527 ( 
.A(n_1873),
.Y(n_2527)
);

AND2x4_ASAP7_75t_L g2528 ( 
.A(n_2174),
.B(n_1733),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2165),
.Y(n_2529)
);

AOI22xp33_ASAP7_75t_L g2530 ( 
.A1(n_2075),
.A2(n_2083),
.B1(n_2098),
.B2(n_2093),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2165),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_1998),
.B(n_2001),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2001),
.B(n_2008),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2008),
.B(n_2017),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2177),
.Y(n_2535)
);

BUFx2_ASAP7_75t_L g2536 ( 
.A(n_1599),
.Y(n_2536)
);

AND2x4_ASAP7_75t_L g2537 ( 
.A(n_1733),
.B(n_1761),
.Y(n_2537)
);

BUFx2_ASAP7_75t_L g2538 ( 
.A(n_1599),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2177),
.Y(n_2539)
);

BUFx2_ASAP7_75t_L g2540 ( 
.A(n_1599),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2177),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2184),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_SL g2543 ( 
.A(n_2155),
.B(n_2179),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2017),
.B(n_2020),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_2048),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2184),
.Y(n_2546)
);

AND2x6_ASAP7_75t_SL g2547 ( 
.A(n_1805),
.B(n_1575),
.Y(n_2547)
);

INVx3_ASAP7_75t_L g2548 ( 
.A(n_1873),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2020),
.B(n_2021),
.Y(n_2549)
);

AND2x4_ASAP7_75t_L g2550 ( 
.A(n_1733),
.B(n_1761),
.Y(n_2550)
);

AOI22xp5_ASAP7_75t_L g2551 ( 
.A1(n_2075),
.A2(n_2093),
.B1(n_2098),
.B2(n_2083),
.Y(n_2551)
);

INVx3_ASAP7_75t_L g2552 ( 
.A(n_1873),
.Y(n_2552)
);

HB1xp67_ASAP7_75t_L g2553 ( 
.A(n_1876),
.Y(n_2553)
);

NOR2xp33_ASAP7_75t_L g2554 ( 
.A(n_2076),
.B(n_2077),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2184),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2021),
.B(n_2027),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2027),
.B(n_2028),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2028),
.B(n_2031),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_2048),
.Y(n_2559)
);

AND2x4_ASAP7_75t_L g2560 ( 
.A(n_1761),
.B(n_1776),
.Y(n_2560)
);

BUFx6f_ASAP7_75t_L g2561 ( 
.A(n_2060),
.Y(n_2561)
);

BUFx6f_ASAP7_75t_L g2562 ( 
.A(n_2060),
.Y(n_2562)
);

BUFx6f_ASAP7_75t_L g2563 ( 
.A(n_2060),
.Y(n_2563)
);

OR2x6_ASAP7_75t_L g2564 ( 
.A(n_1652),
.B(n_1894),
.Y(n_2564)
);

BUFx6f_ASAP7_75t_L g2565 ( 
.A(n_2060),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_1884),
.B(n_2031),
.Y(n_2566)
);

BUFx8_ASAP7_75t_L g2567 ( 
.A(n_2060),
.Y(n_2567)
);

AOI22xp5_ASAP7_75t_L g2568 ( 
.A1(n_2104),
.A2(n_2123),
.B1(n_2149),
.B2(n_2113),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2032),
.B(n_2035),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2032),
.B(n_2035),
.Y(n_2570)
);

AND2x2_ASAP7_75t_L g2571 ( 
.A(n_1884),
.B(n_2037),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2080),
.B(n_2101),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_1715),
.Y(n_2573)
);

AOI22xp33_ASAP7_75t_L g2574 ( 
.A1(n_2104),
.A2(n_2113),
.B1(n_2149),
.B2(n_2123),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_1715),
.Y(n_2575)
);

BUFx6f_ASAP7_75t_L g2576 ( 
.A(n_2060),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_1638),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_1638),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_1722),
.Y(n_2579)
);

BUFx12f_ASAP7_75t_L g2580 ( 
.A(n_1686),
.Y(n_2580)
);

INVx3_ASAP7_75t_L g2581 ( 
.A(n_1873),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_2172),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_L g2583 ( 
.A(n_2106),
.B(n_2111),
.Y(n_2583)
);

AND2x4_ASAP7_75t_L g2584 ( 
.A(n_1776),
.B(n_1937),
.Y(n_2584)
);

NOR3xp33_ASAP7_75t_SL g2585 ( 
.A(n_1575),
.B(n_1617),
.C(n_1607),
.Y(n_2585)
);

OR2x6_ASAP7_75t_L g2586 ( 
.A(n_1894),
.B(n_1608),
.Y(n_2586)
);

AND2x4_ASAP7_75t_L g2587 ( 
.A(n_1776),
.B(n_1937),
.Y(n_2587)
);

INVx3_ASAP7_75t_L g2588 ( 
.A(n_1873),
.Y(n_2588)
);

AOI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2169),
.A2(n_1530),
.B1(n_2097),
.B2(n_1543),
.Y(n_2589)
);

OR2x2_ASAP7_75t_SL g2590 ( 
.A(n_1737),
.B(n_2037),
.Y(n_2590)
);

BUFx6f_ASAP7_75t_L g2591 ( 
.A(n_2110),
.Y(n_2591)
);

BUFx6f_ASAP7_75t_SL g2592 ( 
.A(n_2110),
.Y(n_2592)
);

BUFx4f_ASAP7_75t_L g2593 ( 
.A(n_2110),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_1722),
.Y(n_2594)
);

OR2x4_ASAP7_75t_L g2595 ( 
.A(n_1760),
.B(n_1883),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2050),
.B(n_2052),
.Y(n_2596)
);

INVx4_ASAP7_75t_L g2597 ( 
.A(n_2110),
.Y(n_2597)
);

BUFx6f_ASAP7_75t_L g2598 ( 
.A(n_2110),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2050),
.B(n_2052),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_SL g2600 ( 
.A(n_1675),
.B(n_1801),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_1884),
.B(n_2061),
.Y(n_2601)
);

AND2x2_ASAP7_75t_SL g2602 ( 
.A(n_1610),
.B(n_1632),
.Y(n_2602)
);

AOI22xp33_ASAP7_75t_L g2603 ( 
.A1(n_2169),
.A2(n_1530),
.B1(n_1585),
.B2(n_1569),
.Y(n_2603)
);

BUFx6f_ASAP7_75t_L g2604 ( 
.A(n_2110),
.Y(n_2604)
);

AND2x6_ASAP7_75t_L g2605 ( 
.A(n_1565),
.B(n_1937),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_R g2606 ( 
.A(n_1897),
.B(n_1903),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_1656),
.Y(n_2607)
);

AND2x2_ASAP7_75t_SL g2608 ( 
.A(n_1632),
.B(n_1769),
.Y(n_2608)
);

XNOR2xp5_ASAP7_75t_L g2609 ( 
.A(n_1566),
.B(n_1585),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_1729),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_1657),
.Y(n_2611)
);

BUFx6f_ASAP7_75t_L g2612 ( 
.A(n_1565),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_1729),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_1657),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_1731),
.Y(n_2615)
);

HB1xp67_ASAP7_75t_L g2616 ( 
.A(n_1876),
.Y(n_2616)
);

NAND2x1p5_ASAP7_75t_L g2617 ( 
.A(n_1698),
.B(n_1702),
.Y(n_2617)
);

BUFx4_ASAP7_75t_SL g2618 ( 
.A(n_2172),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2119),
.A2(n_2142),
.B1(n_2131),
.B2(n_1617),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_L g2620 ( 
.A(n_1588),
.B(n_1633),
.Y(n_2620)
);

BUFx10_ASAP7_75t_L g2621 ( 
.A(n_1765),
.Y(n_2621)
);

HB1xp67_ASAP7_75t_L g2622 ( 
.A(n_1914),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_1657),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_1776),
.B(n_1937),
.Y(n_2624)
);

HAxp5_ASAP7_75t_L g2625 ( 
.A(n_1536),
.B(n_1607),
.CON(n_2625),
.SN(n_2625)
);

AOI22xp33_ASAP7_75t_L g2626 ( 
.A1(n_1569),
.A2(n_1566),
.B1(n_1613),
.B2(n_1601),
.Y(n_2626)
);

NAND2xp33_ASAP7_75t_SL g2627 ( 
.A(n_1767),
.B(n_1754),
.Y(n_2627)
);

OR2x2_ASAP7_75t_L g2628 ( 
.A(n_2061),
.B(n_2065),
.Y(n_2628)
);

AND2x4_ASAP7_75t_L g2629 ( 
.A(n_1776),
.B(n_1937),
.Y(n_2629)
);

CKINVDCx20_ASAP7_75t_R g2630 ( 
.A(n_1661),
.Y(n_2630)
);

A2O1A1Ixp33_ASAP7_75t_L g2631 ( 
.A1(n_1546),
.A2(n_1540),
.B(n_1675),
.C(n_1564),
.Y(n_2631)
);

A2O1A1Ixp33_ASAP7_75t_L g2632 ( 
.A1(n_1546),
.A2(n_1540),
.B(n_1564),
.C(n_1646),
.Y(n_2632)
);

BUFx5_ASAP7_75t_L g2633 ( 
.A(n_1727),
.Y(n_2633)
);

BUFx2_ASAP7_75t_L g2634 ( 
.A(n_1599),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_1625),
.B(n_1623),
.Y(n_2635)
);

HB1xp67_ASAP7_75t_L g2636 ( 
.A(n_1914),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_1673),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_1731),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_1554),
.Y(n_2639)
);

BUFx2_ASAP7_75t_L g2640 ( 
.A(n_1606),
.Y(n_2640)
);

INVx1_ASAP7_75t_SL g2641 ( 
.A(n_1896),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2065),
.B(n_2066),
.Y(n_2642)
);

OR2x6_ASAP7_75t_L g2643 ( 
.A(n_1608),
.B(n_1566),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_1673),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_1554),
.Y(n_2645)
);

BUFx3_ASAP7_75t_L g2646 ( 
.A(n_2059),
.Y(n_2646)
);

BUFx6f_ASAP7_75t_L g2647 ( 
.A(n_1565),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_1560),
.Y(n_2648)
);

AND2x6_ASAP7_75t_SL g2649 ( 
.A(n_1813),
.B(n_1839),
.Y(n_2649)
);

INVx1_ASAP7_75t_SL g2650 ( 
.A(n_1896),
.Y(n_2650)
);

CKINVDCx11_ASAP7_75t_R g2651 ( 
.A(n_1927),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_R g2652 ( 
.A(n_1897),
.B(n_1903),
.Y(n_2652)
);

INVx5_ASAP7_75t_L g2653 ( 
.A(n_1565),
.Y(n_2653)
);

HB1xp67_ASAP7_75t_L g2654 ( 
.A(n_1914),
.Y(n_2654)
);

NOR2xp67_ASAP7_75t_L g2655 ( 
.A(n_1655),
.B(n_1802),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_1677),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_1560),
.Y(n_2657)
);

OR2x6_ASAP7_75t_L g2658 ( 
.A(n_1979),
.B(n_2009),
.Y(n_2658)
);

AND2x4_ASAP7_75t_L g2659 ( 
.A(n_1597),
.B(n_1835),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_R g2660 ( 
.A(n_1897),
.B(n_1903),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_1677),
.Y(n_2661)
);

AOI22xp5_ASAP7_75t_L g2662 ( 
.A1(n_1626),
.A2(n_1646),
.B1(n_1620),
.B2(n_1653),
.Y(n_2662)
);

HB1xp67_ASAP7_75t_L g2663 ( 
.A(n_1898),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_1561),
.Y(n_2664)
);

AOI22xp5_ASAP7_75t_L g2665 ( 
.A1(n_1626),
.A2(n_1672),
.B1(n_1653),
.B2(n_1735),
.Y(n_2665)
);

INVx3_ASAP7_75t_L g2666 ( 
.A(n_1887),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2066),
.B(n_2067),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2067),
.B(n_2068),
.Y(n_2668)
);

AND2x4_ASAP7_75t_L g2669 ( 
.A(n_1597),
.B(n_1835),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2068),
.B(n_2070),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2070),
.B(n_2072),
.Y(n_2671)
);

INVxp67_ASAP7_75t_SL g2672 ( 
.A(n_1902),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_1898),
.Y(n_2673)
);

BUFx3_ASAP7_75t_L g2674 ( 
.A(n_2059),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_1677),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2072),
.B(n_2081),
.Y(n_2676)
);

INVx2_ASAP7_75t_SL g2677 ( 
.A(n_1609),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_1561),
.Y(n_2678)
);

CKINVDCx6p67_ASAP7_75t_R g2679 ( 
.A(n_1923),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2081),
.B(n_2082),
.Y(n_2680)
);

CKINVDCx5p33_ASAP7_75t_R g2681 ( 
.A(n_1848),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2082),
.B(n_2090),
.Y(n_2682)
);

AND2x4_ASAP7_75t_L g2683 ( 
.A(n_1597),
.B(n_1835),
.Y(n_2683)
);

NAND3xp33_ASAP7_75t_L g2684 ( 
.A(n_1660),
.B(n_1699),
.C(n_2045),
.Y(n_2684)
);

BUFx2_ASAP7_75t_L g2685 ( 
.A(n_1606),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_1579),
.Y(n_2686)
);

OR2x6_ASAP7_75t_L g2687 ( 
.A(n_2045),
.B(n_1692),
.Y(n_2687)
);

BUFx2_ASAP7_75t_L g2688 ( 
.A(n_1606),
.Y(n_2688)
);

AND2x4_ASAP7_75t_L g2689 ( 
.A(n_1597),
.B(n_1835),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2090),
.B(n_2092),
.Y(n_2690)
);

HB1xp67_ASAP7_75t_L g2691 ( 
.A(n_1898),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2092),
.B(n_2107),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2107),
.B(n_2109),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_1579),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_1582),
.Y(n_2695)
);

BUFx6f_ASAP7_75t_L g2696 ( 
.A(n_1565),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_1848),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_1582),
.Y(n_2698)
);

NOR3xp33_ASAP7_75t_SL g2699 ( 
.A(n_1813),
.B(n_1680),
.C(n_1889),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_L g2700 ( 
.A(n_1672),
.B(n_2036),
.Y(n_2700)
);

INVx4_ASAP7_75t_L g2701 ( 
.A(n_1923),
.Y(n_2701)
);

INVx5_ASAP7_75t_L g2702 ( 
.A(n_1565),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_L g2703 ( 
.A(n_2036),
.B(n_2132),
.Y(n_2703)
);

NAND2xp33_ASAP7_75t_R g2704 ( 
.A(n_1655),
.B(n_1762),
.Y(n_2704)
);

AOI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_1735),
.A2(n_1671),
.B1(n_2114),
.B2(n_2109),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_1589),
.Y(n_2706)
);

INVxp67_ASAP7_75t_SL g2707 ( 
.A(n_1902),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2114),
.B(n_2117),
.Y(n_2708)
);

BUFx3_ASAP7_75t_L g2709 ( 
.A(n_2059),
.Y(n_2709)
);

INVx3_ASAP7_75t_L g2710 ( 
.A(n_1887),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_1719),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_1589),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2117),
.B(n_2118),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2118),
.B(n_2120),
.Y(n_2714)
);

AOI22xp33_ASAP7_75t_L g2715 ( 
.A1(n_1645),
.A2(n_2120),
.B1(n_2127),
.B2(n_2126),
.Y(n_2715)
);

HB1xp67_ASAP7_75t_L g2716 ( 
.A(n_1913),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_1603),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2126),
.B(n_2127),
.Y(n_2718)
);

NOR3xp33_ASAP7_75t_SL g2719 ( 
.A(n_1680),
.B(n_1889),
.C(n_1840),
.Y(n_2719)
);

NOR2xp33_ASAP7_75t_L g2720 ( 
.A(n_2132),
.B(n_1717),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2130),
.B(n_2135),
.Y(n_2721)
);

BUFx6f_ASAP7_75t_L g2722 ( 
.A(n_1565),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_1603),
.Y(n_2723)
);

INVx1_ASAP7_75t_SL g2724 ( 
.A(n_1743),
.Y(n_2724)
);

AOI22xp5_ASAP7_75t_L g2725 ( 
.A1(n_2130),
.A2(n_2137),
.B1(n_2140),
.B2(n_2135),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2137),
.B(n_2140),
.Y(n_2726)
);

BUFx2_ASAP7_75t_L g2727 ( 
.A(n_1606),
.Y(n_2727)
);

INVxp67_ASAP7_75t_L g2728 ( 
.A(n_1883),
.Y(n_2728)
);

CKINVDCx20_ASAP7_75t_R g2729 ( 
.A(n_1927),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2146),
.B(n_2151),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_1682),
.Y(n_2731)
);

AND2x4_ASAP7_75t_L g2732 ( 
.A(n_1597),
.B(n_1835),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_1612),
.Y(n_2733)
);

BUFx2_ASAP7_75t_L g2734 ( 
.A(n_1756),
.Y(n_2734)
);

INVxp67_ASAP7_75t_L g2735 ( 
.A(n_1905),
.Y(n_2735)
);

BUFx6f_ASAP7_75t_L g2736 ( 
.A(n_1704),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_1612),
.Y(n_2737)
);

BUFx6f_ASAP7_75t_L g2738 ( 
.A(n_1704),
.Y(n_2738)
);

INVx3_ASAP7_75t_L g2739 ( 
.A(n_1887),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2146),
.B(n_2151),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_1624),
.Y(n_2741)
);

NOR2xp33_ASAP7_75t_L g2742 ( 
.A(n_1717),
.B(n_1810),
.Y(n_2742)
);

OR2x2_ASAP7_75t_SL g2743 ( 
.A(n_2152),
.B(n_2153),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_1624),
.Y(n_2744)
);

OR2x6_ASAP7_75t_L g2745 ( 
.A(n_1692),
.B(n_1983),
.Y(n_2745)
);

NAND2x1p5_ASAP7_75t_L g2746 ( 
.A(n_1755),
.B(n_1785),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_1631),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_1700),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_1631),
.Y(n_2749)
);

AO22x1_ASAP7_75t_L g2750 ( 
.A1(n_2059),
.A2(n_1727),
.B1(n_1811),
.B2(n_1926),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_1684),
.B(n_1801),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2152),
.B(n_2153),
.Y(n_2752)
);

BUFx4f_ASAP7_75t_L g2753 ( 
.A(n_1983),
.Y(n_2753)
);

HB1xp67_ASAP7_75t_L g2754 ( 
.A(n_1913),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2158),
.B(n_2161),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_1700),
.Y(n_2756)
);

NOR3xp33_ASAP7_75t_SL g2757 ( 
.A(n_1840),
.B(n_1823),
.C(n_1839),
.Y(n_2757)
);

AOI211xp5_ASAP7_75t_L g2758 ( 
.A1(n_1699),
.A2(n_1660),
.B(n_1823),
.C(n_1832),
.Y(n_2758)
);

OR2x6_ASAP7_75t_SL g2759 ( 
.A(n_1764),
.B(n_1811),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_1913),
.Y(n_2760)
);

BUFx3_ASAP7_75t_L g2761 ( 
.A(n_2059),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2158),
.B(n_2161),
.Y(n_2762)
);

INVxp67_ASAP7_75t_L g2763 ( 
.A(n_1905),
.Y(n_2763)
);

AND3x1_ASAP7_75t_SL g2764 ( 
.A(n_1744),
.B(n_2099),
.C(n_2040),
.Y(n_2764)
);

AO21x2_ASAP7_75t_L g2765 ( 
.A1(n_1785),
.A2(n_1930),
.B(n_1772),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_1644),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2166),
.B(n_2167),
.Y(n_2767)
);

BUFx3_ASAP7_75t_L g2768 ( 
.A(n_2059),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2166),
.B(n_2167),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2170),
.B(n_2178),
.Y(n_2770)
);

AND2x4_ASAP7_75t_SL g2771 ( 
.A(n_1686),
.B(n_1834),
.Y(n_2771)
);

INVx4_ASAP7_75t_L g2772 ( 
.A(n_1923),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_1719),
.Y(n_2773)
);

INVx1_ASAP7_75t_SL g2774 ( 
.A(n_1743),
.Y(n_2774)
);

HB1xp67_ASAP7_75t_L g2775 ( 
.A(n_1888),
.Y(n_2775)
);

AND2x4_ASAP7_75t_L g2776 ( 
.A(n_1887),
.B(n_1999),
.Y(n_2776)
);

NOR2xp33_ASAP7_75t_R g2777 ( 
.A(n_1897),
.B(n_1903),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_1645),
.A2(n_2170),
.B1(n_2178),
.B2(n_1746),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_1598),
.B(n_1600),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_1700),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_1644),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_1669),
.B(n_1872),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_1598),
.B(n_1600),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_1665),
.Y(n_2784)
);

AND2x4_ASAP7_75t_L g2785 ( 
.A(n_1999),
.B(n_2181),
.Y(n_2785)
);

BUFx3_ASAP7_75t_L g2786 ( 
.A(n_2059),
.Y(n_2786)
);

AOI21x1_ASAP7_75t_L g2787 ( 
.A1(n_1802),
.A2(n_1867),
.B(n_1853),
.Y(n_2787)
);

NOR3xp33_ASAP7_75t_SL g2788 ( 
.A(n_1765),
.B(n_1867),
.C(n_1762),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_1881),
.B(n_1665),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_1611),
.B(n_1615),
.Y(n_2790)
);

INVx4_ASAP7_75t_L g2791 ( 
.A(n_1923),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_1730),
.Y(n_2792)
);

BUFx4f_ASAP7_75t_L g2793 ( 
.A(n_1983),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_1611),
.B(n_1615),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_1730),
.Y(n_2795)
);

AND2x4_ASAP7_75t_L g2796 ( 
.A(n_2181),
.B(n_1581),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_1752),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_1676),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_1618),
.B(n_1627),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_1676),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_1683),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_1881),
.B(n_1683),
.Y(n_2802)
);

NOR2xp33_ASAP7_75t_R g2803 ( 
.A(n_1897),
.B(n_1903),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_R g2804 ( 
.A(n_1983),
.B(n_2054),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_1690),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_1618),
.B(n_1627),
.Y(n_2806)
);

INVx4_ASAP7_75t_L g2807 ( 
.A(n_1923),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_SL g2808 ( 
.A(n_1911),
.B(n_1924),
.Y(n_2808)
);

BUFx12f_ASAP7_75t_L g2809 ( 
.A(n_1686),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_1690),
.Y(n_2810)
);

NOR3xp33_ASAP7_75t_SL g2811 ( 
.A(n_1917),
.B(n_1895),
.C(n_1893),
.Y(n_2811)
);

NOR3xp33_ASAP7_75t_SL g2812 ( 
.A(n_1917),
.B(n_1895),
.C(n_1893),
.Y(n_2812)
);

BUFx3_ASAP7_75t_L g2813 ( 
.A(n_2059),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_1634),
.B(n_1637),
.Y(n_2814)
);

INVx2_ASAP7_75t_SL g2815 ( 
.A(n_1609),
.Y(n_2815)
);

BUFx4f_ASAP7_75t_L g2816 ( 
.A(n_1983),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_1697),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_1634),
.B(n_1637),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_1797),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_1797),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_1799),
.Y(n_2821)
);

AND2x4_ASAP7_75t_L g2822 ( 
.A(n_1581),
.B(n_1587),
.Y(n_2822)
);

NOR2xp33_ASAP7_75t_R g2823 ( 
.A(n_1983),
.B(n_2054),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_1697),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_1639),
.B(n_1640),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_1799),
.Y(n_2826)
);

NOR3xp33_ASAP7_75t_SL g2827 ( 
.A(n_1853),
.B(n_1906),
.C(n_1841),
.Y(n_2827)
);

NOR2xp67_ASAP7_75t_L g2828 ( 
.A(n_1923),
.B(n_1916),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_1639),
.B(n_1640),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_1712),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_1712),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_1911),
.B(n_1924),
.Y(n_2832)
);

BUFx2_ASAP7_75t_L g2833 ( 
.A(n_1756),
.Y(n_2833)
);

INVxp67_ASAP7_75t_SL g2834 ( 
.A(n_1679),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_1959),
.Y(n_2835)
);

INVx3_ASAP7_75t_L g2836 ( 
.A(n_1907),
.Y(n_2836)
);

BUFx6f_ASAP7_75t_L g2837 ( 
.A(n_1755),
.Y(n_2837)
);

NAND2x1p5_ASAP7_75t_L g2838 ( 
.A(n_1548),
.B(n_1570),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_1799),
.Y(n_2839)
);

BUFx6f_ASAP7_75t_L g2840 ( 
.A(n_1938),
.Y(n_2840)
);

AOI22xp33_ASAP7_75t_L g2841 ( 
.A1(n_2221),
.A2(n_2059),
.B1(n_1739),
.B2(n_1596),
.Y(n_2841)
);

CKINVDCx16_ASAP7_75t_R g2842 ( 
.A(n_2378),
.Y(n_2842)
);

AOI21xp5_ASAP7_75t_L g2843 ( 
.A1(n_2302),
.A2(n_1919),
.B(n_1772),
.Y(n_2843)
);

AOI21xp5_ASAP7_75t_L g2844 ( 
.A1(n_2302),
.A2(n_1770),
.B(n_1870),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_2362),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_SL g2846 ( 
.A(n_2213),
.B(n_1724),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2645),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_SL g2848 ( 
.A(n_2213),
.B(n_2313),
.Y(n_2848)
);

AOI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2630),
.A2(n_1723),
.B1(n_1746),
.B2(n_1724),
.Y(n_2849)
);

NOR2xp33_ASAP7_75t_L g2850 ( 
.A(n_2247),
.B(n_1858),
.Y(n_2850)
);

AOI21xp5_ASAP7_75t_L g2851 ( 
.A1(n_2367),
.A2(n_1892),
.B(n_1875),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_SL g2852 ( 
.A(n_2313),
.B(n_1901),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2645),
.Y(n_2853)
);

BUFx2_ASAP7_75t_L g2854 ( 
.A(n_2759),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2233),
.B(n_1959),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2233),
.B(n_1960),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2247),
.B(n_1960),
.Y(n_2857)
);

AOI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2385),
.A2(n_1570),
.B(n_1921),
.Y(n_2858)
);

INVx4_ASAP7_75t_L g2859 ( 
.A(n_2281),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2645),
.Y(n_2860)
);

BUFx2_ASAP7_75t_L g2861 ( 
.A(n_2759),
.Y(n_2861)
);

NAND2x2_ASAP7_75t_L g2862 ( 
.A(n_2242),
.B(n_1744),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2192),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2291),
.A2(n_1706),
.B1(n_1710),
.B2(n_1688),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2291),
.B(n_1858),
.Y(n_2865)
);

NOR2xp33_ASAP7_75t_L g2866 ( 
.A(n_2349),
.B(n_1871),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2249),
.B(n_1964),
.Y(n_2867)
);

NOR2xp33_ASAP7_75t_R g2868 ( 
.A(n_2280),
.B(n_1871),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2249),
.B(n_1964),
.Y(n_2869)
);

A2O1A1Ixp33_ASAP7_75t_L g2870 ( 
.A1(n_2349),
.A2(n_1578),
.B(n_1864),
.C(n_1763),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2648),
.Y(n_2871)
);

AOI21xp5_ASAP7_75t_L g2872 ( 
.A1(n_2215),
.A2(n_1922),
.B(n_1921),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2211),
.B(n_1974),
.Y(n_2873)
);

A2O1A1Ixp33_ASAP7_75t_L g2874 ( 
.A1(n_2338),
.A2(n_1578),
.B(n_1864),
.C(n_1763),
.Y(n_2874)
);

BUFx12f_ASAP7_75t_L g2875 ( 
.A(n_2280),
.Y(n_2875)
);

HB1xp67_ASAP7_75t_L g2876 ( 
.A(n_2475),
.Y(n_2876)
);

O2A1O1Ixp33_ASAP7_75t_L g2877 ( 
.A1(n_2196),
.A2(n_1832),
.B(n_1808),
.C(n_1814),
.Y(n_2877)
);

INVx4_ASAP7_75t_L g2878 ( 
.A(n_2281),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2263),
.B(n_1974),
.Y(n_2879)
);

AOI21xp5_ASAP7_75t_L g2880 ( 
.A1(n_2215),
.A2(n_1922),
.B(n_1771),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2199),
.Y(n_2881)
);

OAI21xp33_ASAP7_75t_L g2882 ( 
.A1(n_2335),
.A2(n_1642),
.B(n_1641),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2263),
.B(n_1988),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2648),
.Y(n_2884)
);

AOI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2220),
.A2(n_1771),
.B(n_1642),
.Y(n_2885)
);

OR2x2_ASAP7_75t_L g2886 ( 
.A(n_2622),
.B(n_1596),
.Y(n_2886)
);

A2O1A1Ixp33_ASAP7_75t_L g2887 ( 
.A1(n_2338),
.A2(n_1774),
.B(n_1792),
.C(n_1751),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2648),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2706),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_SL g2890 ( 
.A(n_2370),
.B(n_1686),
.Y(n_2890)
);

INVx3_ASAP7_75t_L g2891 ( 
.A(n_2192),
.Y(n_2891)
);

NOR2xp33_ASAP7_75t_L g2892 ( 
.A(n_2711),
.B(n_2773),
.Y(n_2892)
);

CKINVDCx16_ASAP7_75t_R g2893 ( 
.A(n_2378),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2706),
.Y(n_2894)
);

AOI22xp33_ASAP7_75t_L g2895 ( 
.A1(n_2221),
.A2(n_1739),
.B1(n_1596),
.B2(n_1723),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2199),
.Y(n_2896)
);

OAI22xp5_ASAP7_75t_SL g2897 ( 
.A1(n_2243),
.A2(n_1688),
.B1(n_1710),
.B2(n_1706),
.Y(n_2897)
);

AOI21xp5_ASAP7_75t_L g2898 ( 
.A1(n_2220),
.A2(n_1650),
.B(n_1641),
.Y(n_2898)
);

NOR3xp33_ASAP7_75t_L g2899 ( 
.A(n_2440),
.B(n_1808),
.C(n_1829),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2284),
.B(n_1988),
.Y(n_2900)
);

AOI21xp5_ASAP7_75t_L g2901 ( 
.A1(n_2631),
.A2(n_1658),
.B(n_1650),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2199),
.Y(n_2902)
);

AOI22xp33_ASAP7_75t_L g2903 ( 
.A1(n_2327),
.A2(n_1791),
.B1(n_1559),
.B2(n_1525),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2706),
.Y(n_2904)
);

BUFx12f_ASAP7_75t_L g2905 ( 
.A(n_2366),
.Y(n_2905)
);

HB1xp67_ASAP7_75t_L g2906 ( 
.A(n_2475),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2284),
.B(n_1992),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2712),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_L g2909 ( 
.A(n_2711),
.B(n_1871),
.Y(n_2909)
);

INVxp67_ASAP7_75t_L g2910 ( 
.A(n_2773),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2199),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2631),
.A2(n_1659),
.B(n_1658),
.Y(n_2912)
);

AO22x1_ASAP7_75t_L g2913 ( 
.A1(n_2672),
.A2(n_1727),
.B1(n_1559),
.B2(n_1545),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2287),
.B(n_1992),
.Y(n_2914)
);

INVx4_ASAP7_75t_L g2915 ( 
.A(n_2281),
.Y(n_2915)
);

INVxp67_ASAP7_75t_L g2916 ( 
.A(n_2635),
.Y(n_2916)
);

AND2x2_ASAP7_75t_SL g2917 ( 
.A(n_2521),
.B(n_1769),
.Y(n_2917)
);

OAI22xp5_ASAP7_75t_L g2918 ( 
.A1(n_2287),
.A2(n_1791),
.B1(n_1774),
.B2(n_1674),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2712),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2712),
.Y(n_2920)
);

A2O1A1Ixp33_ASAP7_75t_SL g2921 ( 
.A1(n_2758),
.A2(n_1918),
.B(n_1909),
.C(n_1920),
.Y(n_2921)
);

AOI22xp33_ASAP7_75t_L g2922 ( 
.A1(n_2327),
.A2(n_1559),
.B1(n_1545),
.B2(n_1525),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2209),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2209),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_2834),
.B(n_1996),
.Y(n_2925)
);

AOI21xp5_ASAP7_75t_L g2926 ( 
.A1(n_2503),
.A2(n_1674),
.B(n_1659),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2390),
.B(n_1636),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2834),
.B(n_2641),
.Y(n_2928)
);

AOI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2503),
.A2(n_2543),
.B(n_2476),
.Y(n_2929)
);

CKINVDCx20_ASAP7_75t_R g2930 ( 
.A(n_2304),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2403),
.B(n_1711),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2543),
.A2(n_1929),
.B(n_1681),
.Y(n_2932)
);

AOI21xp5_ASAP7_75t_L g2933 ( 
.A1(n_2476),
.A2(n_1929),
.B(n_1681),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2641),
.B(n_1996),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2650),
.B(n_1997),
.Y(n_2935)
);

NOR2xp33_ASAP7_75t_L g2936 ( 
.A(n_2403),
.B(n_1711),
.Y(n_2936)
);

NOR3xp33_ASAP7_75t_SL g2937 ( 
.A(n_2440),
.B(n_1906),
.C(n_1869),
.Y(n_2937)
);

NOR2xp67_ASAP7_75t_SL g2938 ( 
.A(n_2399),
.B(n_1907),
.Y(n_2938)
);

NOR2xp33_ASAP7_75t_L g2939 ( 
.A(n_2518),
.B(n_2545),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2650),
.B(n_1997),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2211),
.B(n_2004),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2735),
.B(n_2004),
.Y(n_2942)
);

O2A1O1Ixp33_ASAP7_75t_L g2943 ( 
.A1(n_2196),
.A2(n_1798),
.B(n_1865),
.C(n_1885),
.Y(n_2943)
);

OAI21x1_ASAP7_75t_L g2944 ( 
.A1(n_2787),
.A2(n_1933),
.B(n_1930),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2741),
.Y(n_2945)
);

AOI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2453),
.A2(n_1687),
.B(n_1679),
.Y(n_2946)
);

AOI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2453),
.A2(n_1689),
.B(n_1687),
.Y(n_2947)
);

AOI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_2214),
.A2(n_1691),
.B(n_1689),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2735),
.B(n_2010),
.Y(n_2949)
);

OAI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2316),
.A2(n_2376),
.B(n_2335),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_2518),
.B(n_1711),
.Y(n_2951)
);

O2A1O1Ixp33_ASAP7_75t_L g2952 ( 
.A1(n_2214),
.A2(n_1865),
.B(n_1885),
.C(n_1779),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2763),
.B(n_2010),
.Y(n_2953)
);

OAI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2342),
.A2(n_1750),
.B1(n_1749),
.B2(n_1900),
.Y(n_2954)
);

INVx1_ASAP7_75t_SL g2955 ( 
.A(n_2724),
.Y(n_2955)
);

NOR2xp33_ASAP7_75t_L g2956 ( 
.A(n_2545),
.B(n_1711),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2209),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_SL g2958 ( 
.A(n_2370),
.B(n_1834),
.Y(n_2958)
);

AND2x4_ASAP7_75t_L g2959 ( 
.A(n_2390),
.B(n_1636),
.Y(n_2959)
);

BUFx6f_ASAP7_75t_L g2960 ( 
.A(n_2192),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2209),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2619),
.B(n_1891),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2744),
.Y(n_2963)
);

AOI21xp5_ASAP7_75t_L g2964 ( 
.A1(n_2406),
.A2(n_2315),
.B(n_2632),
.Y(n_2964)
);

A2O1A1Ixp33_ASAP7_75t_L g2965 ( 
.A1(n_2399),
.A2(n_1792),
.B(n_1751),
.C(n_1891),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2744),
.Y(n_2966)
);

NOR2xp67_ASAP7_75t_L g2967 ( 
.A(n_2684),
.B(n_1916),
.Y(n_2967)
);

OR2x6_ASAP7_75t_L g2968 ( 
.A(n_2586),
.B(n_2054),
.Y(n_2968)
);

AOI22xp5_ASAP7_75t_L g2969 ( 
.A1(n_2630),
.A2(n_1842),
.B1(n_1768),
.B2(n_1725),
.Y(n_2969)
);

O2A1O1Ixp5_ASAP7_75t_L g2970 ( 
.A1(n_2406),
.A2(n_1779),
.B(n_1934),
.C(n_1935),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2763),
.B(n_2013),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_SL g2972 ( 
.A(n_2619),
.B(n_1918),
.Y(n_2972)
);

OAI22xp5_ASAP7_75t_L g2973 ( 
.A1(n_2342),
.A2(n_1750),
.B1(n_1749),
.B2(n_1900),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2744),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_SL g2975 ( 
.A(n_2585),
.B(n_1654),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2293),
.B(n_2013),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2293),
.B(n_2026),
.Y(n_2977)
);

BUFx6f_ASAP7_75t_L g2978 ( 
.A(n_2192),
.Y(n_2978)
);

A2O1A1Ixp33_ASAP7_75t_L g2979 ( 
.A1(n_2811),
.A2(n_1842),
.B(n_1768),
.C(n_1862),
.Y(n_2979)
);

BUFx6f_ASAP7_75t_L g2980 ( 
.A(n_2192),
.Y(n_2980)
);

AOI21xp5_ASAP7_75t_L g2981 ( 
.A1(n_2406),
.A2(n_1695),
.B(n_1691),
.Y(n_2981)
);

AOI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_2315),
.A2(n_1696),
.B(n_1695),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_SL g2983 ( 
.A(n_2375),
.B(n_2672),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2766),
.Y(n_2984)
);

NOR3xp33_ASAP7_75t_SL g2985 ( 
.A(n_2559),
.B(n_2582),
.C(n_2344),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2222),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2222),
.Y(n_2987)
);

OAI21xp5_ASAP7_75t_L g2988 ( 
.A1(n_2316),
.A2(n_1654),
.B(n_1920),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2632),
.A2(n_1701),
.B(n_1696),
.Y(n_2989)
);

OAI21xp33_ASAP7_75t_SL g2990 ( 
.A1(n_2326),
.A2(n_1707),
.B(n_1701),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2240),
.B(n_2026),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2766),
.Y(n_2992)
);

AOI21xp5_ASAP7_75t_L g2993 ( 
.A1(n_2281),
.A2(n_1708),
.B(n_1707),
.Y(n_2993)
);

BUFx6f_ASAP7_75t_L g2994 ( 
.A(n_2192),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2830),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_SL g2996 ( 
.A(n_2585),
.B(n_1909),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2240),
.B(n_2042),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2830),
.Y(n_2998)
);

AND2x4_ASAP7_75t_L g2999 ( 
.A(n_2390),
.B(n_1636),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2830),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2255),
.B(n_2042),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2831),
.Y(n_3002)
);

BUFx6f_ASAP7_75t_L g3003 ( 
.A(n_2192),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_SL g3004 ( 
.A(n_2559),
.B(n_1636),
.Y(n_3004)
);

AOI21xp5_ASAP7_75t_L g3005 ( 
.A1(n_2281),
.A2(n_1708),
.B(n_1718),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2831),
.Y(n_3006)
);

NOR2xp33_ASAP7_75t_L g3007 ( 
.A(n_2582),
.B(n_1711),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2831),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2499),
.B(n_1713),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2255),
.B(n_2053),
.Y(n_3010)
);

AND2x2_ASAP7_75t_L g3011 ( 
.A(n_2211),
.B(n_2053),
.Y(n_3011)
);

OR2x2_ASAP7_75t_L g3012 ( 
.A(n_2622),
.B(n_2058),
.Y(n_3012)
);

AND2x4_ASAP7_75t_L g3013 ( 
.A(n_2390),
.B(n_1636),
.Y(n_3013)
);

OAI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2342),
.A2(n_2144),
.B1(n_2105),
.B2(n_2173),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2222),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2188),
.B(n_2058),
.Y(n_3016)
);

BUFx2_ASAP7_75t_L g3017 ( 
.A(n_2759),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2188),
.B(n_2078),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2499),
.B(n_1713),
.Y(n_3019)
);

AOI21xp5_ASAP7_75t_L g3020 ( 
.A1(n_2434),
.A2(n_1741),
.B(n_1718),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2547),
.B(n_2246),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2835),
.Y(n_3022)
);

INVx5_ASAP7_75t_L g3023 ( 
.A(n_2586),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2222),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2835),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2189),
.B(n_2078),
.Y(n_3026)
);

NOR2xp33_ASAP7_75t_L g3027 ( 
.A(n_2547),
.B(n_1713),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_SL g3028 ( 
.A(n_2294),
.B(n_1931),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2216),
.B(n_2085),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2189),
.B(n_2085),
.Y(n_3030)
);

NOR2xp33_ASAP7_75t_L g3031 ( 
.A(n_2246),
.B(n_1713),
.Y(n_3031)
);

OAI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2363),
.A2(n_2409),
.B1(n_2243),
.B2(n_2372),
.Y(n_3032)
);

AND2x4_ASAP7_75t_L g3033 ( 
.A(n_2395),
.B(n_2016),
.Y(n_3033)
);

AOI21xp5_ASAP7_75t_L g3034 ( 
.A1(n_2434),
.A2(n_1741),
.B(n_1718),
.Y(n_3034)
);

BUFx3_ASAP7_75t_L g3035 ( 
.A(n_2520),
.Y(n_3035)
);

NOR2xp33_ASAP7_75t_L g3036 ( 
.A(n_2202),
.B(n_1713),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2193),
.B(n_2086),
.Y(n_3037)
);

INVx1_ASAP7_75t_SL g3038 ( 
.A(n_2724),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_L g3039 ( 
.A(n_2202),
.B(n_1725),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2193),
.B(n_2086),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2207),
.B(n_2087),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2207),
.B(n_2087),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2835),
.Y(n_3043)
);

O2A1O1Ixp5_ASAP7_75t_L g3044 ( 
.A1(n_2600),
.A2(n_1907),
.B(n_1925),
.C(n_1915),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2223),
.Y(n_3045)
);

AO32x1_ASAP7_75t_L g3046 ( 
.A1(n_2230),
.A2(n_1888),
.A3(n_2173),
.B1(n_2162),
.B2(n_2089),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2225),
.B(n_2089),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2223),
.Y(n_3048)
);

BUFx6f_ASAP7_75t_L g3049 ( 
.A(n_2192),
.Y(n_3049)
);

BUFx3_ASAP7_75t_L g3050 ( 
.A(n_2520),
.Y(n_3050)
);

CKINVDCx11_ASAP7_75t_R g3051 ( 
.A(n_2237),
.Y(n_3051)
);

NOR2xp67_ASAP7_75t_L g3052 ( 
.A(n_2684),
.B(n_1899),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2573),
.Y(n_3053)
);

A2O1A1Ixp33_ASAP7_75t_L g3054 ( 
.A1(n_2811),
.A2(n_2812),
.B(n_2251),
.C(n_2707),
.Y(n_3054)
);

AOI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2434),
.A2(n_1741),
.B(n_1747),
.Y(n_3055)
);

O2A1O1Ixp33_ASAP7_75t_SL g3056 ( 
.A1(n_2326),
.A2(n_1880),
.B(n_1882),
.C(n_1874),
.Y(n_3056)
);

NOR2xp33_ASAP7_75t_L g3057 ( 
.A(n_2308),
.B(n_1725),
.Y(n_3057)
);

O2A1O1Ixp33_ASAP7_75t_L g3058 ( 
.A1(n_2625),
.A2(n_2376),
.B(n_2230),
.C(n_2295),
.Y(n_3058)
);

AOI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_2434),
.A2(n_1747),
.B(n_1728),
.Y(n_3059)
);

CKINVDCx5p33_ASAP7_75t_R g3060 ( 
.A(n_2362),
.Y(n_3060)
);

AOI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_2434),
.A2(n_1747),
.B(n_1728),
.Y(n_3061)
);

OAI22x1_ASAP7_75t_L g3062 ( 
.A1(n_2707),
.A2(n_2105),
.B1(n_2100),
.B2(n_2162),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2225),
.B(n_2100),
.Y(n_3063)
);

INVx4_ASAP7_75t_L g3064 ( 
.A(n_2442),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_2308),
.B(n_1725),
.Y(n_3065)
);

OR2x4_ASAP7_75t_L g3066 ( 
.A(n_2300),
.B(n_1764),
.Y(n_3066)
);

O2A1O1Ixp33_ASAP7_75t_L g3067 ( 
.A1(n_2625),
.A2(n_1869),
.B(n_1868),
.C(n_1882),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2232),
.B(n_2116),
.Y(n_3068)
);

AND2x4_ASAP7_75t_L g3069 ( 
.A(n_2395),
.B(n_2016),
.Y(n_3069)
);

NOR3xp33_ASAP7_75t_L g3070 ( 
.A(n_2782),
.B(n_2116),
.C(n_2159),
.Y(n_3070)
);

HB1xp67_ASAP7_75t_L g3071 ( 
.A(n_2522),
.Y(n_3071)
);

O2A1O1Ixp33_ASAP7_75t_L g3072 ( 
.A1(n_2625),
.A2(n_1868),
.B(n_1886),
.C(n_2124),
.Y(n_3072)
);

OAI22xp5_ASAP7_75t_SL g3073 ( 
.A1(n_2226),
.A2(n_1773),
.B1(n_1663),
.B2(n_1725),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2232),
.B(n_2124),
.Y(n_3074)
);

AOI21xp5_ASAP7_75t_L g3075 ( 
.A1(n_2442),
.A2(n_1678),
.B(n_1899),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2442),
.A2(n_1678),
.B(n_1899),
.Y(n_3076)
);

OAI21xp5_ASAP7_75t_L g3077 ( 
.A1(n_2372),
.A2(n_1908),
.B(n_1912),
.Y(n_3077)
);

AOI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2442),
.A2(n_1915),
.B(n_1908),
.Y(n_3078)
);

AOI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_2442),
.A2(n_2423),
.B(n_2437),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2251),
.B(n_1593),
.Y(n_3080)
);

AOI21xp5_ASAP7_75t_L g3081 ( 
.A1(n_2423),
.A2(n_2437),
.B(n_2260),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2573),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2260),
.A2(n_1912),
.B(n_1782),
.Y(n_3083)
);

O2A1O1Ixp5_ASAP7_75t_L g3084 ( 
.A1(n_2295),
.A2(n_1907),
.B(n_1881),
.C(n_1778),
.Y(n_3084)
);

OAI21xp33_ASAP7_75t_L g3085 ( 
.A1(n_2719),
.A2(n_1879),
.B(n_1878),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2298),
.B(n_2141),
.Y(n_3086)
);

INVx2_ASAP7_75t_L g3087 ( 
.A(n_2223),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_L g3088 ( 
.A(n_2365),
.B(n_2418),
.Y(n_3088)
);

BUFx3_ASAP7_75t_L g3089 ( 
.A(n_2520),
.Y(n_3089)
);

AOI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2432),
.A2(n_1782),
.B(n_1778),
.Y(n_3090)
);

NOR2xp33_ASAP7_75t_L g3091 ( 
.A(n_2365),
.B(n_2141),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_2223),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2298),
.B(n_2144),
.Y(n_3093)
);

AND2x4_ASAP7_75t_L g3094 ( 
.A(n_2395),
.B(n_2016),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2575),
.Y(n_3095)
);

OAI22xp5_ASAP7_75t_L g3096 ( 
.A1(n_2363),
.A2(n_2159),
.B1(n_1663),
.B2(n_1773),
.Y(n_3096)
);

NOR2xp33_ASAP7_75t_SL g3097 ( 
.A(n_2375),
.B(n_1834),
.Y(n_3097)
);

CKINVDCx5p33_ASAP7_75t_R g3098 ( 
.A(n_2279),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2234),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2234),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_SL g3101 ( 
.A(n_2827),
.B(n_1593),
.Y(n_3101)
);

OAI21xp33_ASAP7_75t_L g3102 ( 
.A1(n_2719),
.A2(n_2699),
.B(n_2488),
.Y(n_3102)
);

NOR2xp33_ASAP7_75t_L g3103 ( 
.A(n_2418),
.B(n_1593),
.Y(n_3103)
);

AOI21xp5_ASAP7_75t_L g3104 ( 
.A1(n_2394),
.A2(n_1587),
.B(n_1861),
.Y(n_3104)
);

O2A1O1Ixp33_ASAP7_75t_L g3105 ( 
.A1(n_2782),
.A2(n_1886),
.B(n_1862),
.C(n_1764),
.Y(n_3105)
);

NOR2xp33_ASAP7_75t_L g3106 ( 
.A(n_2728),
.B(n_1667),
.Y(n_3106)
);

NOR2xp33_ASAP7_75t_L g3107 ( 
.A(n_2728),
.B(n_1667),
.Y(n_3107)
);

BUFx12f_ASAP7_75t_L g3108 ( 
.A(n_2366),
.Y(n_3108)
);

BUFx2_ASAP7_75t_L g3109 ( 
.A(n_2391),
.Y(n_3109)
);

INVx1_ASAP7_75t_SL g3110 ( 
.A(n_2774),
.Y(n_3110)
);

OAI321xp33_ASAP7_75t_L g3111 ( 
.A1(n_2626),
.A2(n_1635),
.A3(n_2122),
.B1(n_2096),
.B2(n_1938),
.C(n_2071),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2320),
.B(n_1734),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2320),
.B(n_1734),
.Y(n_3113)
);

A2O1A1Ixp33_ASAP7_75t_L g3114 ( 
.A1(n_2812),
.A2(n_1863),
.B(n_2133),
.C(n_1567),
.Y(n_3114)
);

OAI21x1_ASAP7_75t_L g3115 ( 
.A1(n_2787),
.A2(n_1635),
.B(n_2122),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_SL g3116 ( 
.A(n_2827),
.B(n_1667),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_SL g3117 ( 
.A(n_2699),
.B(n_1716),
.Y(n_3117)
);

OAI21x1_ASAP7_75t_L g3118 ( 
.A1(n_2787),
.A2(n_1635),
.B(n_2122),
.Y(n_3118)
);

BUFx2_ASAP7_75t_L g3119 ( 
.A(n_2391),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2575),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_L g3121 ( 
.A(n_2649),
.B(n_1716),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2636),
.B(n_1738),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2234),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_SL g3124 ( 
.A(n_2757),
.B(n_1716),
.Y(n_3124)
);

NAND3xp33_ASAP7_75t_SL g3125 ( 
.A(n_2226),
.B(n_1635),
.C(n_2122),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2636),
.B(n_1738),
.Y(n_3126)
);

AOI22xp33_ASAP7_75t_L g3127 ( 
.A1(n_2487),
.A2(n_1559),
.B1(n_1545),
.B2(n_1567),
.Y(n_3127)
);

AND2x4_ASAP7_75t_L g3128 ( 
.A(n_2395),
.B(n_2016),
.Y(n_3128)
);

AND2x4_ASAP7_75t_L g3129 ( 
.A(n_2404),
.B(n_2016),
.Y(n_3129)
);

O2A1O1Ixp5_ASAP7_75t_SL g3130 ( 
.A1(n_2484),
.A2(n_1745),
.B(n_1742),
.C(n_1775),
.Y(n_3130)
);

BUFx2_ASAP7_75t_L g3131 ( 
.A(n_2391),
.Y(n_3131)
);

AOI21x1_ASAP7_75t_L g3132 ( 
.A1(n_2655),
.A2(n_1786),
.B(n_1783),
.Y(n_3132)
);

OAI22xp5_ASAP7_75t_L g3133 ( 
.A1(n_2409),
.A2(n_1834),
.B1(n_1756),
.B2(n_2054),
.Y(n_3133)
);

BUFx6f_ASAP7_75t_L g3134 ( 
.A(n_2195),
.Y(n_3134)
);

AND2x4_ASAP7_75t_L g3135 ( 
.A(n_2404),
.B(n_2180),
.Y(n_3135)
);

INVx3_ASAP7_75t_L g3136 ( 
.A(n_2195),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2579),
.Y(n_3137)
);

BUFx2_ASAP7_75t_SL g3138 ( 
.A(n_2633),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2234),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2654),
.B(n_1742),
.Y(n_3140)
);

AND2x4_ASAP7_75t_L g3141 ( 
.A(n_2404),
.B(n_2180),
.Y(n_3141)
);

INVx2_ASAP7_75t_SL g3142 ( 
.A(n_2347),
.Y(n_3142)
);

OAI22xp5_ASAP7_75t_L g3143 ( 
.A1(n_2381),
.A2(n_2464),
.B1(n_2574),
.B2(n_2530),
.Y(n_3143)
);

CKINVDCx20_ASAP7_75t_R g3144 ( 
.A(n_2304),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_2216),
.B(n_2180),
.Y(n_3145)
);

AOI21x1_ASAP7_75t_L g3146 ( 
.A1(n_2828),
.A2(n_1783),
.B(n_1745),
.Y(n_3146)
);

CKINVDCx20_ASAP7_75t_R g3147 ( 
.A(n_2309),
.Y(n_3147)
);

A2O1A1Ixp33_ASAP7_75t_L g3148 ( 
.A1(n_2551),
.A2(n_1863),
.B(n_2133),
.C(n_2102),
.Y(n_3148)
);

A2O1A1Ixp33_ASAP7_75t_L g3149 ( 
.A1(n_2551),
.A2(n_1863),
.B(n_2133),
.C(n_2102),
.Y(n_3149)
);

AOI21xp5_ASAP7_75t_L g3150 ( 
.A1(n_2808),
.A2(n_1758),
.B(n_1756),
.Y(n_3150)
);

AOI22xp5_ASAP7_75t_L g3151 ( 
.A1(n_2626),
.A2(n_2180),
.B1(n_1727),
.B2(n_1559),
.Y(n_3151)
);

HB1xp67_ASAP7_75t_L g3152 ( 
.A(n_2522),
.Y(n_3152)
);

CKINVDCx20_ASAP7_75t_R g3153 ( 
.A(n_2309),
.Y(n_3153)
);

A2O1A1Ixp33_ASAP7_75t_L g3154 ( 
.A1(n_2568),
.A2(n_2300),
.B(n_2665),
.C(n_2751),
.Y(n_3154)
);

BUFx6f_ASAP7_75t_L g3155 ( 
.A(n_2195),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2579),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2594),
.Y(n_3157)
);

AOI21xp33_ASAP7_75t_L g3158 ( 
.A1(n_2484),
.A2(n_1843),
.B(n_1827),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2654),
.B(n_1827),
.Y(n_3159)
);

A2O1A1Ixp33_ASAP7_75t_L g3160 ( 
.A1(n_2568),
.A2(n_2019),
.B(n_2102),
.C(n_2091),
.Y(n_3160)
);

NAND2xp33_ASAP7_75t_L g3161 ( 
.A(n_2467),
.B(n_2277),
.Y(n_3161)
);

AOI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_2627),
.A2(n_2832),
.B(n_2449),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_R g3163 ( 
.A(n_2237),
.B(n_2019),
.Y(n_3163)
);

HB1xp67_ASAP7_75t_L g3164 ( 
.A(n_2553),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2757),
.B(n_2180),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2322),
.B(n_1843),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_2216),
.B(n_2091),
.Y(n_3167)
);

BUFx6f_ASAP7_75t_L g3168 ( 
.A(n_2195),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2824),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_SL g3170 ( 
.A(n_2467),
.B(n_2091),
.Y(n_3170)
);

AOI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_2487),
.A2(n_1866),
.B1(n_1877),
.B2(n_1727),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2248),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2824),
.Y(n_3173)
);

NOR2xp33_ASAP7_75t_L g3174 ( 
.A(n_2649),
.B(n_1609),
.Y(n_3174)
);

BUFx6f_ASAP7_75t_L g3175 ( 
.A(n_2195),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2248),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2594),
.Y(n_3177)
);

BUFx3_ASAP7_75t_L g3178 ( 
.A(n_2520),
.Y(n_3178)
);

A2O1A1Ixp33_ASAP7_75t_L g3179 ( 
.A1(n_2665),
.A2(n_2084),
.B(n_2054),
.C(n_1860),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2729),
.B(n_1609),
.Y(n_3180)
);

OAI22x1_ASAP7_75t_L g3181 ( 
.A1(n_2487),
.A2(n_1740),
.B1(n_1847),
.B2(n_1775),
.Y(n_3181)
);

AND2x4_ASAP7_75t_L g3182 ( 
.A(n_2404),
.B(n_1727),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_SL g3183 ( 
.A(n_2620),
.B(n_1812),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2322),
.B(n_1866),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2610),
.Y(n_3185)
);

CKINVDCx16_ASAP7_75t_R g3186 ( 
.A(n_2505),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2332),
.B(n_2779),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2332),
.B(n_1866),
.Y(n_3188)
);

NOR2xp67_ASAP7_75t_L g3189 ( 
.A(n_2200),
.B(n_1836),
.Y(n_3189)
);

BUFx3_ASAP7_75t_L g3190 ( 
.A(n_2646),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2610),
.Y(n_3191)
);

BUFx10_ASAP7_75t_L g3192 ( 
.A(n_2242),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2613),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_SL g3194 ( 
.A(n_2620),
.B(n_2662),
.Y(n_3194)
);

INVxp67_ASAP7_75t_L g3195 ( 
.A(n_2635),
.Y(n_3195)
);

NOR2x1_ASAP7_75t_R g3196 ( 
.A(n_2288),
.B(n_1609),
.Y(n_3196)
);

OR2x6_ASAP7_75t_L g3197 ( 
.A(n_2586),
.B(n_2084),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2779),
.B(n_1877),
.Y(n_3198)
);

AO21x1_ASAP7_75t_L g3199 ( 
.A1(n_2336),
.A2(n_1847),
.B(n_1795),
.Y(n_3199)
);

INVx1_ASAP7_75t_SL g3200 ( 
.A(n_2774),
.Y(n_3200)
);

BUFx6f_ASAP7_75t_L g3201 ( 
.A(n_2195),
.Y(n_3201)
);

O2A1O1Ixp5_ASAP7_75t_SL g3202 ( 
.A1(n_2187),
.A2(n_1790),
.B(n_1833),
.C(n_1748),
.Y(n_3202)
);

BUFx6f_ASAP7_75t_L g3203 ( 
.A(n_2195),
.Y(n_3203)
);

AND2x4_ASAP7_75t_L g3204 ( 
.A(n_2447),
.B(n_1727),
.Y(n_3204)
);

A2O1A1Ixp33_ASAP7_75t_L g3205 ( 
.A1(n_2751),
.A2(n_1877),
.B(n_1836),
.C(n_1788),
.Y(n_3205)
);

BUFx6f_ASAP7_75t_L g3206 ( 
.A(n_2195),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2783),
.B(n_1825),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2613),
.Y(n_3208)
);

O2A1O1Ixp33_ASAP7_75t_SL g3209 ( 
.A1(n_2554),
.A2(n_1757),
.B(n_1825),
.C(n_1748),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_SL g3210 ( 
.A(n_2572),
.B(n_1757),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2783),
.B(n_1795),
.Y(n_3211)
);

BUFx2_ASAP7_75t_L g3212 ( 
.A(n_2450),
.Y(n_3212)
);

AOI21xp5_ASAP7_75t_L g3213 ( 
.A1(n_2572),
.A2(n_2583),
.B(n_2586),
.Y(n_3213)
);

BUFx6f_ASAP7_75t_L g3214 ( 
.A(n_2236),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_2493),
.B(n_1740),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_L g3216 ( 
.A(n_2729),
.B(n_1740),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_2586),
.A2(n_1818),
.B(n_1844),
.Y(n_3217)
);

INVx1_ASAP7_75t_SL g3218 ( 
.A(n_2299),
.Y(n_3218)
);

BUFx2_ASAP7_75t_L g3219 ( 
.A(n_2450),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2248),
.Y(n_3220)
);

INVx2_ASAP7_75t_SL g3221 ( 
.A(n_2388),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_2586),
.A2(n_1817),
.B(n_1838),
.Y(n_3222)
);

BUFx6f_ASAP7_75t_L g3223 ( 
.A(n_2236),
.Y(n_3223)
);

OAI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_2466),
.A2(n_2515),
.B(n_2325),
.Y(n_3224)
);

CKINVDCx5p33_ASAP7_75t_R g3225 ( 
.A(n_2191),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_2245),
.B(n_1820),
.Y(n_3226)
);

AND2x4_ASAP7_75t_L g3227 ( 
.A(n_2447),
.B(n_2456),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_SL g3228 ( 
.A(n_2493),
.B(n_1859),
.Y(n_3228)
);

AO22x1_ASAP7_75t_L g3229 ( 
.A1(n_2681),
.A2(n_1727),
.B1(n_1859),
.B2(n_1850),
.Y(n_3229)
);

AOI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_2586),
.A2(n_1826),
.B(n_1837),
.Y(n_3230)
);

BUFx10_ASAP7_75t_L g3231 ( 
.A(n_2771),
.Y(n_3231)
);

AOI21xp5_ASAP7_75t_L g3232 ( 
.A1(n_2658),
.A2(n_1826),
.B(n_1837),
.Y(n_3232)
);

BUFx8_ASAP7_75t_L g3233 ( 
.A(n_2261),
.Y(n_3233)
);

OR2x6_ASAP7_75t_SL g3234 ( 
.A(n_2681),
.B(n_1845),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_2790),
.B(n_1833),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2248),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2790),
.B(n_2794),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2615),
.Y(n_3238)
);

HB1xp67_ASAP7_75t_L g3239 ( 
.A(n_2553),
.Y(n_3239)
);

BUFx6f_ASAP7_75t_L g3240 ( 
.A(n_2236),
.Y(n_3240)
);

INVx3_ASAP7_75t_L g3241 ( 
.A(n_2236),
.Y(n_3241)
);

A2O1A1Ixp33_ASAP7_75t_SL g3242 ( 
.A1(n_2703),
.A2(n_1803),
.B(n_1753),
.C(n_1766),
.Y(n_3242)
);

AOI22xp5_ASAP7_75t_L g3243 ( 
.A1(n_2464),
.A2(n_2530),
.B1(n_2574),
.B2(n_2346),
.Y(n_3243)
);

NOR2xp33_ASAP7_75t_L g3244 ( 
.A(n_2651),
.B(n_1727),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_2259),
.Y(n_3245)
);

CKINVDCx5p33_ASAP7_75t_R g3246 ( 
.A(n_2191),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2794),
.B(n_1845),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_2259),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2615),
.Y(n_3249)
);

CKINVDCx5p33_ASAP7_75t_R g3250 ( 
.A(n_2341),
.Y(n_3250)
);

A2O1A1Ixp33_ASAP7_75t_SL g3251 ( 
.A1(n_2703),
.A2(n_1800),
.B(n_1753),
.C(n_1766),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2638),
.Y(n_3252)
);

A2O1A1Ixp33_ASAP7_75t_L g3253 ( 
.A1(n_2603),
.A2(n_1790),
.B(n_1803),
.C(n_1800),
.Y(n_3253)
);

A2O1A1Ixp33_ASAP7_75t_L g3254 ( 
.A1(n_2603),
.A2(n_1854),
.B(n_1850),
.C(n_1793),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2799),
.B(n_1820),
.Y(n_3255)
);

CKINVDCx20_ASAP7_75t_R g3256 ( 
.A(n_2237),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_2259),
.Y(n_3257)
);

O2A1O1Ixp5_ASAP7_75t_L g3258 ( 
.A1(n_2750),
.A2(n_2325),
.B(n_2593),
.C(n_2445),
.Y(n_3258)
);

BUFx3_ASAP7_75t_L g3259 ( 
.A(n_2646),
.Y(n_3259)
);

A2O1A1Ixp33_ASAP7_75t_L g3260 ( 
.A1(n_2589),
.A2(n_1854),
.B(n_1787),
.C(n_1793),
.Y(n_3260)
);

BUFx2_ASAP7_75t_L g3261 ( 
.A(n_2450),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_2436),
.B(n_1856),
.Y(n_3262)
);

NOR2xp33_ASAP7_75t_L g3263 ( 
.A(n_2651),
.B(n_1727),
.Y(n_3263)
);

HB1xp67_ASAP7_75t_L g3264 ( 
.A(n_2616),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2259),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_2278),
.Y(n_3266)
);

O2A1O1Ixp33_ASAP7_75t_L g3267 ( 
.A1(n_2325),
.A2(n_1852),
.B(n_1855),
.C(n_1796),
.Y(n_3267)
);

INVx1_ASAP7_75t_SL g3268 ( 
.A(n_2299),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2799),
.B(n_1820),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_2278),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_2806),
.B(n_1849),
.Y(n_3271)
);

BUFx3_ASAP7_75t_L g3272 ( 
.A(n_2646),
.Y(n_3272)
);

A2O1A1Ixp33_ASAP7_75t_L g3273 ( 
.A1(n_2589),
.A2(n_1787),
.B(n_1794),
.C(n_1796),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_2806),
.B(n_1824),
.Y(n_3274)
);

AOI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_2658),
.A2(n_1806),
.B(n_1807),
.Y(n_3275)
);

HB1xp67_ASAP7_75t_L g3276 ( 
.A(n_2616),
.Y(n_3276)
);

NOR2xp33_ASAP7_75t_SL g3277 ( 
.A(n_2288),
.B(n_2447),
.Y(n_3277)
);

BUFx10_ASAP7_75t_L g3278 ( 
.A(n_2771),
.Y(n_3278)
);

AOI22xp33_ASAP7_75t_L g3279 ( 
.A1(n_2346),
.A2(n_1856),
.B1(n_1851),
.B2(n_1828),
.Y(n_3279)
);

AND2x4_ASAP7_75t_L g3280 ( 
.A(n_2447),
.B(n_1804),
.Y(n_3280)
);

OR2x2_ASAP7_75t_L g3281 ( 
.A(n_2743),
.B(n_2388),
.Y(n_3281)
);

NOR2xp33_ASAP7_75t_L g3282 ( 
.A(n_2430),
.B(n_1815),
.Y(n_3282)
);

BUFx12f_ASAP7_75t_L g3283 ( 
.A(n_2366),
.Y(n_3283)
);

OAI21xp33_ASAP7_75t_L g3284 ( 
.A1(n_2788),
.A2(n_2277),
.B(n_2705),
.Y(n_3284)
);

BUFx2_ASAP7_75t_L g3285 ( 
.A(n_2461),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2638),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_2814),
.B(n_1804),
.Y(n_3287)
);

O2A1O1Ixp5_ASAP7_75t_L g3288 ( 
.A1(n_2750),
.A2(n_1821),
.B(n_1815),
.C(n_1809),
.Y(n_3288)
);

NOR3xp33_ASAP7_75t_SL g3289 ( 
.A(n_2341),
.B(n_1855),
.C(n_1852),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2814),
.B(n_1804),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_2278),
.Y(n_3291)
);

OR2x6_ASAP7_75t_L g3292 ( 
.A(n_2564),
.B(n_1809),
.Y(n_3292)
);

NOR2xp33_ASAP7_75t_L g3293 ( 
.A(n_2430),
.B(n_1821),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_2236),
.A2(n_1809),
.B(n_1819),
.Y(n_3294)
);

CKINVDCx20_ASAP7_75t_R g3295 ( 
.A(n_2237),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2818),
.B(n_1819),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2639),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_SL g3298 ( 
.A(n_2436),
.B(n_1851),
.Y(n_3298)
);

BUFx3_ASAP7_75t_L g3299 ( 
.A(n_2646),
.Y(n_3299)
);

NOR2xp33_ASAP7_75t_L g3300 ( 
.A(n_2430),
.B(n_1824),
.Y(n_3300)
);

BUFx6f_ASAP7_75t_L g3301 ( 
.A(n_2236),
.Y(n_3301)
);

CKINVDCx8_ASAP7_75t_R g3302 ( 
.A(n_2697),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2639),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2657),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_2278),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2818),
.B(n_1830),
.Y(n_3306)
);

AO32x1_ASAP7_75t_L g3307 ( 
.A1(n_2257),
.A2(n_1830),
.A3(n_1831),
.B1(n_1849),
.B2(n_1851),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_2305),
.Y(n_3308)
);

AND2x4_ASAP7_75t_L g3309 ( 
.A(n_2456),
.B(n_1831),
.Y(n_3309)
);

BUFx3_ASAP7_75t_L g3310 ( 
.A(n_2674),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_2825),
.B(n_1831),
.Y(n_3311)
);

CKINVDCx5p33_ASAP7_75t_R g3312 ( 
.A(n_2344),
.Y(n_3312)
);

NOR3xp33_ASAP7_75t_L g3313 ( 
.A(n_2515),
.B(n_2700),
.C(n_2266),
.Y(n_3313)
);

OR2x2_ASAP7_75t_L g3314 ( 
.A(n_2743),
.B(n_1828),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_2825),
.B(n_1846),
.Y(n_3315)
);

HB1xp67_ASAP7_75t_L g3316 ( 
.A(n_2461),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_2305),
.Y(n_3317)
);

A2O1A1Ixp33_ASAP7_75t_L g3318 ( 
.A1(n_2456),
.A2(n_2462),
.B(n_2490),
.C(n_2485),
.Y(n_3318)
);

OAI22xp5_ASAP7_75t_L g3319 ( 
.A1(n_2725),
.A2(n_2715),
.B1(n_2459),
.B2(n_2743),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_SL g3320 ( 
.A(n_2436),
.B(n_2785),
.Y(n_3320)
);

BUFx3_ASAP7_75t_L g3321 ( 
.A(n_2674),
.Y(n_3321)
);

BUFx3_ASAP7_75t_L g3322 ( 
.A(n_2674),
.Y(n_3322)
);

BUFx2_ASAP7_75t_L g3323 ( 
.A(n_2564),
.Y(n_3323)
);

O2A1O1Ixp33_ASAP7_75t_L g3324 ( 
.A1(n_2439),
.A2(n_2788),
.B(n_2187),
.C(n_2256),
.Y(n_3324)
);

AOI221xp5_ASAP7_75t_L g3325 ( 
.A1(n_2715),
.A2(n_2770),
.B1(n_2778),
.B2(n_2700),
.C(n_2393),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_2829),
.B(n_2267),
.Y(n_3326)
);

AOI22xp33_ASAP7_75t_L g3327 ( 
.A1(n_2346),
.A2(n_2602),
.B1(n_2608),
.B2(n_2609),
.Y(n_3327)
);

O2A1O1Ixp33_ASAP7_75t_L g3328 ( 
.A1(n_2439),
.A2(n_2256),
.B(n_2307),
.C(n_2238),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_2305),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_SL g3330 ( 
.A(n_2436),
.B(n_2785),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2829),
.B(n_2267),
.Y(n_3331)
);

BUFx12f_ASAP7_75t_L g3332 ( 
.A(n_2366),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2271),
.B(n_2566),
.Y(n_3333)
);

INVx3_ASAP7_75t_L g3334 ( 
.A(n_2236),
.Y(n_3334)
);

INVx3_ASAP7_75t_L g3335 ( 
.A(n_2239),
.Y(n_3335)
);

CKINVDCx5p33_ASAP7_75t_R g3336 ( 
.A(n_2373),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_L g3337 ( 
.A(n_2770),
.B(n_2186),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_2186),
.B(n_2197),
.Y(n_3338)
);

INVx3_ASAP7_75t_L g3339 ( 
.A(n_2239),
.Y(n_3339)
);

O2A1O1Ixp5_ASAP7_75t_L g3340 ( 
.A1(n_2750),
.A2(n_2445),
.B(n_2593),
.C(n_2785),
.Y(n_3340)
);

O2A1O1Ixp5_ASAP7_75t_SL g3341 ( 
.A1(n_2238),
.A2(n_2333),
.B(n_2307),
.C(n_2775),
.Y(n_3341)
);

O2A1O1Ixp33_ASAP7_75t_L g3342 ( 
.A1(n_2333),
.A2(n_2618),
.B(n_2266),
.C(n_2331),
.Y(n_3342)
);

AOI22xp33_ASAP7_75t_L g3343 ( 
.A1(n_2346),
.A2(n_2602),
.B1(n_2608),
.B2(n_2609),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_2186),
.B(n_2197),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_R g3345 ( 
.A(n_2505),
.B(n_2373),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_2245),
.B(n_2319),
.Y(n_3346)
);

O2A1O1Ixp33_ASAP7_75t_L g3347 ( 
.A1(n_2257),
.A2(n_2331),
.B(n_2266),
.C(n_2742),
.Y(n_3347)
);

O2A1O1Ixp33_ASAP7_75t_L g3348 ( 
.A1(n_2257),
.A2(n_2331),
.B(n_2742),
.C(n_2483),
.Y(n_3348)
);

INVx5_ASAP7_75t_L g3349 ( 
.A(n_2564),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_2271),
.B(n_2566),
.Y(n_3350)
);

BUFx2_ASAP7_75t_L g3351 ( 
.A(n_2564),
.Y(n_3351)
);

BUFx3_ASAP7_75t_L g3352 ( 
.A(n_2674),
.Y(n_3352)
);

OAI22x1_ASAP7_75t_L g3353 ( 
.A1(n_2609),
.A2(n_2697),
.B1(n_2725),
.B2(n_2203),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_2566),
.B(n_2571),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_2571),
.B(n_2601),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_2245),
.B(n_2319),
.Y(n_3356)
);

NOR2xp33_ASAP7_75t_R g3357 ( 
.A(n_2465),
.B(n_2497),
.Y(n_3357)
);

O2A1O1Ixp33_ASAP7_75t_L g3358 ( 
.A1(n_2426),
.A2(n_2483),
.B(n_2508),
.C(n_2496),
.Y(n_3358)
);

NOR2x1_ASAP7_75t_L g3359 ( 
.A(n_2421),
.B(n_2765),
.Y(n_3359)
);

INVx5_ASAP7_75t_L g3360 ( 
.A(n_2564),
.Y(n_3360)
);

BUFx4f_ASAP7_75t_L g3361 ( 
.A(n_2679),
.Y(n_3361)
);

INVx6_ASAP7_75t_L g3362 ( 
.A(n_2371),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_2571),
.B(n_2601),
.Y(n_3363)
);

CKINVDCx8_ASAP7_75t_R g3364 ( 
.A(n_2231),
.Y(n_3364)
);

BUFx4f_ASAP7_75t_L g3365 ( 
.A(n_2679),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_2601),
.B(n_2282),
.Y(n_3366)
);

OAI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_2459),
.A2(n_2628),
.B1(n_2778),
.B2(n_2398),
.Y(n_3367)
);

INVx2_ASAP7_75t_L g3368 ( 
.A(n_2305),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_2282),
.B(n_2292),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_2657),
.Y(n_3370)
);

INVx1_ASAP7_75t_SL g3371 ( 
.A(n_2426),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_2314),
.Y(n_3372)
);

INVx2_ASAP7_75t_SL g3373 ( 
.A(n_2421),
.Y(n_3373)
);

AOI21x1_ASAP7_75t_L g3374 ( 
.A1(n_2785),
.A2(n_2217),
.B(n_2203),
.Y(n_3374)
);

BUFx6f_ASAP7_75t_L g3375 ( 
.A(n_2239),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_SL g3376 ( 
.A(n_2785),
.B(n_2621),
.Y(n_3376)
);

BUFx12f_ASAP7_75t_L g3377 ( 
.A(n_2366),
.Y(n_3377)
);

OAI22xp5_ASAP7_75t_L g3378 ( 
.A1(n_2459),
.A2(n_2628),
.B1(n_2398),
.B2(n_2410),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_SL g3379 ( 
.A(n_2785),
.B(n_2621),
.Y(n_3379)
);

AND2x4_ASAP7_75t_L g3380 ( 
.A(n_2456),
.B(n_2462),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_2292),
.B(n_2789),
.Y(n_3381)
);

HB1xp67_ASAP7_75t_L g3382 ( 
.A(n_2427),
.Y(n_3382)
);

AOI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_2753),
.A2(n_2816),
.B(n_2793),
.Y(n_3383)
);

NAND3xp33_ASAP7_75t_SL g3384 ( 
.A(n_2465),
.B(n_2389),
.C(n_2496),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_2664),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_2664),
.Y(n_3386)
);

INVx3_ASAP7_75t_SL g3387 ( 
.A(n_2679),
.Y(n_3387)
);

OAI22xp5_ASAP7_75t_L g3388 ( 
.A1(n_2628),
.A2(n_2410),
.B1(n_2420),
.B2(n_2393),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_SL g3389 ( 
.A(n_2621),
.B(n_2217),
.Y(n_3389)
);

BUFx2_ASAP7_75t_L g3390 ( 
.A(n_2564),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_SL g3391 ( 
.A(n_2621),
.B(n_2796),
.Y(n_3391)
);

INVx1_ASAP7_75t_SL g3392 ( 
.A(n_2508),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_2789),
.B(n_2802),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_2789),
.B(n_2802),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_2802),
.B(n_2392),
.Y(n_3395)
);

BUFx6f_ASAP7_75t_L g3396 ( 
.A(n_2239),
.Y(n_3396)
);

OR2x6_ASAP7_75t_L g3397 ( 
.A(n_2564),
.B(n_2462),
.Y(n_3397)
);

OAI21x1_ASAP7_75t_L g3398 ( 
.A1(n_2746),
.A2(n_2617),
.B(n_2227),
.Y(n_3398)
);

NAND3xp33_ASAP7_75t_SL g3399 ( 
.A(n_2389),
.B(n_2519),
.C(n_2720),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2678),
.Y(n_3400)
);

A2O1A1Ixp33_ASAP7_75t_SL g3401 ( 
.A1(n_2413),
.A2(n_2516),
.B(n_2470),
.C(n_2527),
.Y(n_3401)
);

NOR2xp33_ASAP7_75t_L g3402 ( 
.A(n_2197),
.B(n_2206),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_2314),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_L g3404 ( 
.A(n_2206),
.B(n_2420),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_2392),
.B(n_2198),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_2198),
.B(n_2670),
.Y(n_3406)
);

BUFx3_ASAP7_75t_L g3407 ( 
.A(n_2709),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_2198),
.B(n_2670),
.Y(n_3408)
);

OAI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_2424),
.A2(n_2438),
.B1(n_2446),
.B2(n_2429),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_2319),
.B(n_2343),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_2670),
.B(n_2682),
.Y(n_3411)
);

BUFx6f_ASAP7_75t_L g3412 ( 
.A(n_2239),
.Y(n_3412)
);

OAI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_2424),
.A2(n_2438),
.B1(n_2446),
.B2(n_2429),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_2206),
.B(n_2468),
.Y(n_3414)
);

OAI22xp5_ASAP7_75t_L g3415 ( 
.A1(n_2468),
.A2(n_2481),
.B1(n_2506),
.B2(n_2482),
.Y(n_3415)
);

A2O1A1Ixp33_ASAP7_75t_L g3416 ( 
.A1(n_2462),
.A2(n_2490),
.B(n_2512),
.C(n_2485),
.Y(n_3416)
);

CKINVDCx5p33_ASAP7_75t_R g3417 ( 
.A(n_2497),
.Y(n_3417)
);

BUFx2_ASAP7_75t_L g3418 ( 
.A(n_2239),
.Y(n_3418)
);

A2O1A1Ixp33_ASAP7_75t_L g3419 ( 
.A1(n_2485),
.A2(n_2512),
.B(n_2490),
.C(n_2212),
.Y(n_3419)
);

OAI22xp5_ASAP7_75t_L g3420 ( 
.A1(n_2481),
.A2(n_2506),
.B1(n_2513),
.B2(n_2482),
.Y(n_3420)
);

AOI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_2602),
.A2(n_2608),
.B1(n_2720),
.B2(n_2764),
.Y(n_3421)
);

OAI22xp5_ASAP7_75t_L g3422 ( 
.A1(n_2513),
.A2(n_2526),
.B1(n_2532),
.B2(n_2523),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_2682),
.B(n_2692),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_2621),
.B(n_2796),
.Y(n_3424)
);

O2A1O1Ixp33_ASAP7_75t_L g3425 ( 
.A1(n_2519),
.A2(n_2218),
.B(n_2241),
.C(n_2203),
.Y(n_3425)
);

BUFx10_ASAP7_75t_L g3426 ( 
.A(n_2771),
.Y(n_3426)
);

AOI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_2765),
.A2(n_2445),
.B(n_2595),
.Y(n_3427)
);

OAI22xp5_ASAP7_75t_L g3428 ( 
.A1(n_2523),
.A2(n_2532),
.B1(n_2533),
.B2(n_2526),
.Y(n_3428)
);

HB1xp67_ASAP7_75t_L g3429 ( 
.A(n_2427),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_2682),
.B(n_2692),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_SL g3431 ( 
.A(n_2288),
.B(n_2485),
.Y(n_3431)
);

AOI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_2595),
.A2(n_2677),
.B(n_2469),
.Y(n_3432)
);

AOI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_2595),
.A2(n_2677),
.B(n_2469),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_L g3434 ( 
.A(n_2692),
.B(n_2721),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_SL g3435 ( 
.A(n_2796),
.B(n_2212),
.Y(n_3435)
);

BUFx6f_ASAP7_75t_L g3436 ( 
.A(n_2239),
.Y(n_3436)
);

AOI22xp33_ASAP7_75t_L g3437 ( 
.A1(n_2602),
.A2(n_2608),
.B1(n_2643),
.B2(n_2212),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_2678),
.Y(n_3438)
);

INVx3_ASAP7_75t_L g3439 ( 
.A(n_2244),
.Y(n_3439)
);

INVx1_ASAP7_75t_SL g3440 ( 
.A(n_2231),
.Y(n_3440)
);

OAI22xp5_ASAP7_75t_L g3441 ( 
.A1(n_2533),
.A2(n_2544),
.B1(n_2549),
.B2(n_2534),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_2244),
.A2(n_2268),
.B(n_2252),
.Y(n_3442)
);

HB1xp67_ASAP7_75t_L g3443 ( 
.A(n_2876),
.Y(n_3443)
);

A2O1A1Ixp33_ASAP7_75t_L g3444 ( 
.A1(n_3058),
.A2(n_2512),
.B(n_2490),
.C(n_2212),
.Y(n_3444)
);

AOI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_2848),
.A2(n_2595),
.B(n_2512),
.Y(n_3445)
);

OAI21x1_ASAP7_75t_L g3446 ( 
.A1(n_2944),
.A2(n_2617),
.B(n_2227),
.Y(n_3446)
);

OAI21x1_ASAP7_75t_L g3447 ( 
.A1(n_3202),
.A2(n_2838),
.B(n_2836),
.Y(n_3447)
);

INVx3_ASAP7_75t_L g3448 ( 
.A(n_3436),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_2855),
.B(n_2775),
.Y(n_3449)
);

OAI21x1_ASAP7_75t_L g3450 ( 
.A1(n_3132),
.A2(n_3130),
.B(n_3427),
.Y(n_3450)
);

O2A1O1Ixp33_ASAP7_75t_SL g3451 ( 
.A1(n_3102),
.A2(n_2544),
.B(n_2549),
.C(n_2534),
.Y(n_3451)
);

INVx4_ASAP7_75t_L g3452 ( 
.A(n_3361),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2855),
.B(n_2686),
.Y(n_3453)
);

OAI22x1_ASAP7_75t_L g3454 ( 
.A1(n_3421),
.A2(n_2833),
.B1(n_2734),
.B2(n_2218),
.Y(n_3454)
);

INVxp67_ASAP7_75t_L g3455 ( 
.A(n_2892),
.Y(n_3455)
);

A2O1A1Ixp33_ASAP7_75t_L g3456 ( 
.A1(n_3154),
.A2(n_2235),
.B(n_2262),
.C(n_2709),
.Y(n_3456)
);

INVx1_ASAP7_75t_SL g3457 ( 
.A(n_3218),
.Y(n_3457)
);

OAI21x1_ASAP7_75t_L g3458 ( 
.A1(n_3132),
.A2(n_2838),
.B(n_2836),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_3346),
.B(n_2537),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_2856),
.B(n_2686),
.Y(n_3460)
);

INVx2_ASAP7_75t_SL g3461 ( 
.A(n_3382),
.Y(n_3461)
);

INVx1_ASAP7_75t_SL g3462 ( 
.A(n_3218),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_2847),
.Y(n_3463)
);

OAI21xp5_ASAP7_75t_L g3464 ( 
.A1(n_2950),
.A2(n_2241),
.B(n_2218),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_2847),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_2856),
.B(n_2694),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_2857),
.B(n_2694),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_2857),
.B(n_2695),
.Y(n_3468)
);

OAI21xp5_ASAP7_75t_L g3469 ( 
.A1(n_2950),
.A2(n_2258),
.B(n_2241),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_2988),
.A2(n_2252),
.B(n_2244),
.Y(n_3470)
);

OAI21x1_ASAP7_75t_L g3471 ( 
.A1(n_3130),
.A2(n_2838),
.B(n_2836),
.Y(n_3471)
);

NAND3xp33_ASAP7_75t_SL g3472 ( 
.A(n_3102),
.B(n_2652),
.C(n_2606),
.Y(n_3472)
);

AND2x4_ASAP7_75t_L g3473 ( 
.A(n_3182),
.B(n_2709),
.Y(n_3473)
);

NOR2xp67_ASAP7_75t_L g3474 ( 
.A(n_3349),
.B(n_2288),
.Y(n_3474)
);

OAI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_3032),
.A2(n_2270),
.B(n_2258),
.Y(n_3475)
);

CKINVDCx5p33_ASAP7_75t_R g3476 ( 
.A(n_2875),
.Y(n_3476)
);

OA21x2_ASAP7_75t_L g3477 ( 
.A1(n_3288),
.A2(n_2270),
.B(n_2258),
.Y(n_3477)
);

INVx2_ASAP7_75t_SL g3478 ( 
.A(n_3429),
.Y(n_3478)
);

OAI21xp5_ASAP7_75t_L g3479 ( 
.A1(n_3032),
.A2(n_2272),
.B(n_2270),
.Y(n_3479)
);

BUFx2_ASAP7_75t_L g3480 ( 
.A(n_2854),
.Y(n_3480)
);

BUFx6f_ASAP7_75t_L g3481 ( 
.A(n_2960),
.Y(n_3481)
);

BUFx6f_ASAP7_75t_L g3482 ( 
.A(n_2960),
.Y(n_3482)
);

BUFx8_ASAP7_75t_L g3483 ( 
.A(n_2875),
.Y(n_3483)
);

BUFx3_ASAP7_75t_L g3484 ( 
.A(n_2905),
.Y(n_3484)
);

OA22x2_ASAP7_75t_L g3485 ( 
.A1(n_3421),
.A2(n_2643),
.B1(n_2311),
.B2(n_2405),
.Y(n_3485)
);

OAI22xp5_ASAP7_75t_L g3486 ( 
.A1(n_3243),
.A2(n_3343),
.B1(n_3327),
.B2(n_2846),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3237),
.B(n_2695),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_SL g3488 ( 
.A(n_2842),
.B(n_2235),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3237),
.B(n_2698),
.Y(n_3489)
);

NAND3x1_ASAP7_75t_L g3490 ( 
.A(n_2964),
.B(n_2451),
.C(n_2343),
.Y(n_3490)
);

A2O1A1Ixp33_ASAP7_75t_L g3491 ( 
.A1(n_3054),
.A2(n_2262),
.B(n_2235),
.C(n_2709),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3326),
.B(n_2698),
.Y(n_3492)
);

BUFx3_ASAP7_75t_L g3493 ( 
.A(n_2905),
.Y(n_3493)
);

AO31x2_ASAP7_75t_L g3494 ( 
.A1(n_3199),
.A2(n_2833),
.A3(n_2734),
.B(n_2318),
.Y(n_3494)
);

OAI21xp33_ASAP7_75t_L g3495 ( 
.A1(n_2990),
.A2(n_2262),
.B(n_2235),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_2853),
.Y(n_3496)
);

OAI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_2967),
.A2(n_2339),
.B(n_2272),
.Y(n_3497)
);

AO21x2_ASAP7_75t_L g3498 ( 
.A1(n_3199),
.A2(n_2204),
.B(n_2201),
.Y(n_3498)
);

NAND2x1p5_ASAP7_75t_L g3499 ( 
.A(n_3361),
.B(n_2200),
.Y(n_3499)
);

CKINVDCx5p33_ASAP7_75t_R g3500 ( 
.A(n_2875),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_2853),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3326),
.B(n_2717),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3331),
.B(n_3378),
.Y(n_3503)
);

AOI211x1_ASAP7_75t_L g3504 ( 
.A1(n_3284),
.A2(n_2996),
.B(n_3194),
.C(n_2929),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_3245),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3331),
.B(n_2717),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3245),
.Y(n_3507)
);

NAND2x1_ASAP7_75t_L g3508 ( 
.A(n_2938),
.B(n_2413),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3378),
.B(n_2723),
.Y(n_3509)
);

BUFx2_ASAP7_75t_L g3510 ( 
.A(n_2854),
.Y(n_3510)
);

A2O1A1Ixp33_ASAP7_75t_L g3511 ( 
.A1(n_3284),
.A2(n_2262),
.B(n_2768),
.C(n_2761),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3346),
.B(n_2537),
.Y(n_3512)
);

INVx3_ASAP7_75t_L g3513 ( 
.A(n_2960),
.Y(n_3513)
);

OAI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_2967),
.A2(n_2339),
.B(n_2272),
.Y(n_3514)
);

BUFx6f_ASAP7_75t_L g3515 ( 
.A(n_2960),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_2860),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_3243),
.A2(n_3143),
.B1(n_2972),
.B2(n_2850),
.Y(n_3517)
);

A2O1A1Ixp33_ASAP7_75t_L g3518 ( 
.A1(n_2870),
.A2(n_2761),
.B(n_2786),
.C(n_2768),
.Y(n_3518)
);

AOI221xp5_ASAP7_75t_SL g3519 ( 
.A1(n_3014),
.A2(n_2339),
.B1(n_2590),
.B2(n_2556),
.C(n_2558),
.Y(n_3519)
);

OAI22xp5_ASAP7_75t_L g3520 ( 
.A1(n_3143),
.A2(n_2865),
.B1(n_2897),
.B2(n_3325),
.Y(n_3520)
);

AOI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_2946),
.A2(n_2252),
.B(n_2244),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3388),
.B(n_2723),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_L g3523 ( 
.A(n_3186),
.B(n_2556),
.Y(n_3523)
);

O2A1O1Ixp5_ASAP7_75t_L g3524 ( 
.A1(n_2975),
.A2(n_2962),
.B(n_2852),
.C(n_3096),
.Y(n_3524)
);

BUFx2_ASAP7_75t_L g3525 ( 
.A(n_2861),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_2860),
.Y(n_3526)
);

AO21x2_ASAP7_75t_L g3527 ( 
.A1(n_3242),
.A2(n_2204),
.B(n_2201),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_SL g3528 ( 
.A(n_2842),
.B(n_2633),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_2871),
.Y(n_3529)
);

NAND2x1_ASAP7_75t_L g3530 ( 
.A(n_2938),
.B(n_2413),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_2947),
.A2(n_2252),
.B(n_2244),
.Y(n_3531)
);

AOI21xp5_ASAP7_75t_L g3532 ( 
.A1(n_3081),
.A2(n_2268),
.B(n_2252),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3046),
.A2(n_2269),
.B(n_2268),
.Y(n_3533)
);

OAI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_3162),
.A2(n_2443),
.B(n_2734),
.Y(n_3534)
);

OAI21x1_ASAP7_75t_SL g3535 ( 
.A1(n_3324),
.A2(n_3374),
.B(n_3328),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_2871),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_2884),
.Y(n_3537)
);

BUFx6f_ASAP7_75t_L g3538 ( 
.A(n_2960),
.Y(n_3538)
);

OAI22x1_ASAP7_75t_L g3539 ( 
.A1(n_3151),
.A2(n_2833),
.B1(n_2737),
.B2(n_2747),
.Y(n_3539)
);

AO21x2_ASAP7_75t_L g3540 ( 
.A1(n_3251),
.A2(n_2219),
.B(n_2208),
.Y(n_3540)
);

AO21x1_ASAP7_75t_L g3541 ( 
.A1(n_3096),
.A2(n_2737),
.B(n_2733),
.Y(n_3541)
);

INVxp67_ASAP7_75t_SL g3542 ( 
.A(n_3358),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_2893),
.B(n_2633),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_2884),
.Y(n_3544)
);

OR2x2_ASAP7_75t_L g3545 ( 
.A(n_3366),
.B(n_2590),
.Y(n_3545)
);

O2A1O1Ixp5_ASAP7_75t_L g3546 ( 
.A1(n_3028),
.A2(n_2776),
.B(n_2470),
.C(n_2516),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3046),
.A2(n_3162),
.B(n_3209),
.Y(n_3547)
);

AOI221x1_ASAP7_75t_L g3548 ( 
.A1(n_2899),
.A2(n_2231),
.B1(n_2516),
.B2(n_2470),
.C(n_2413),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3388),
.B(n_2733),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_2888),
.Y(n_3550)
);

NOR3xp33_ASAP7_75t_SL g3551 ( 
.A(n_3225),
.B(n_2704),
.C(n_2348),
.Y(n_3551)
);

A2O1A1Ixp33_ASAP7_75t_L g3552 ( 
.A1(n_2874),
.A2(n_2761),
.B(n_2786),
.C(n_2768),
.Y(n_3552)
);

AOI22xp5_ASAP7_75t_L g3553 ( 
.A1(n_2897),
.A2(n_2764),
.B1(n_2311),
.B2(n_2405),
.Y(n_3553)
);

OR2x2_ASAP7_75t_L g3554 ( 
.A(n_3366),
.B(n_2590),
.Y(n_3554)
);

AOI21x1_ASAP7_75t_L g3555 ( 
.A1(n_3146),
.A2(n_2796),
.B(n_2776),
.Y(n_3555)
);

BUFx2_ASAP7_75t_L g3556 ( 
.A(n_2861),
.Y(n_3556)
);

INVx1_ASAP7_75t_SL g3557 ( 
.A(n_3268),
.Y(n_3557)
);

NAND3xp33_ASAP7_75t_SL g3558 ( 
.A(n_2921),
.B(n_2652),
.C(n_2606),
.Y(n_3558)
);

AOI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_3046),
.A2(n_2269),
.B(n_2268),
.Y(n_3559)
);

NAND3x1_ASAP7_75t_L g3560 ( 
.A(n_3213),
.B(n_2451),
.C(n_2343),
.Y(n_3560)
);

AOI22xp5_ASAP7_75t_L g3561 ( 
.A1(n_2864),
.A2(n_2311),
.B1(n_2405),
.B2(n_2351),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_3046),
.A2(n_2269),
.B(n_2268),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_SL g3563 ( 
.A(n_2893),
.B(n_2633),
.Y(n_3563)
);

AO31x2_ASAP7_75t_L g3564 ( 
.A1(n_3062),
.A2(n_2318),
.A3(n_2323),
.B(n_2314),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_SL g3565 ( 
.A1(n_3114),
.A2(n_2768),
.B(n_2761),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_SL g3566 ( 
.A(n_3163),
.B(n_2633),
.Y(n_3566)
);

OAI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_2933),
.A2(n_2443),
.B(n_2351),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3187),
.B(n_2747),
.Y(n_3568)
);

AO32x2_ASAP7_75t_L g3569 ( 
.A1(n_3319),
.A2(n_2396),
.A3(n_2377),
.B1(n_2677),
.B2(n_2469),
.Y(n_3569)
);

NAND2x1p5_ASAP7_75t_L g3570 ( 
.A(n_3361),
.B(n_2200),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3187),
.B(n_2749),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3369),
.B(n_2749),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_2888),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3245),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3369),
.B(n_2781),
.Y(n_3575)
);

INVx4_ASAP7_75t_L g3576 ( 
.A(n_3361),
.Y(n_3576)
);

INVx3_ASAP7_75t_L g3577 ( 
.A(n_3436),
.Y(n_3577)
);

AOI21x1_ASAP7_75t_SL g3578 ( 
.A1(n_2867),
.A2(n_2776),
.B(n_2822),
.Y(n_3578)
);

OA21x2_ASAP7_75t_L g3579 ( 
.A1(n_3084),
.A2(n_2384),
.B(n_2185),
.Y(n_3579)
);

OA22x2_ASAP7_75t_L g3580 ( 
.A1(n_3151),
.A2(n_2643),
.B1(n_2311),
.B2(n_2405),
.Y(n_3580)
);

AOI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_3046),
.A2(n_2269),
.B(n_2268),
.Y(n_3581)
);

OAI21xp5_ASAP7_75t_L g3582 ( 
.A1(n_2932),
.A2(n_2351),
.B(n_2311),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_2889),
.Y(n_3583)
);

AO21x2_ASAP7_75t_L g3584 ( 
.A1(n_3294),
.A2(n_2219),
.B(n_2208),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_SL g3585 ( 
.A1(n_3179),
.A2(n_2813),
.B(n_2786),
.Y(n_3585)
);

INVx1_ASAP7_75t_SL g3586 ( 
.A(n_3268),
.Y(n_3586)
);

NOR2xp67_ASAP7_75t_SL g3587 ( 
.A(n_3364),
.B(n_2425),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_2889),
.Y(n_3588)
);

INVx1_ASAP7_75t_SL g3589 ( 
.A(n_3371),
.Y(n_3589)
);

OAI21xp5_ASAP7_75t_SL g3590 ( 
.A1(n_3014),
.A2(n_2494),
.B(n_2477),
.Y(n_3590)
);

BUFx8_ASAP7_75t_L g3591 ( 
.A(n_2905),
.Y(n_3591)
);

INVx1_ASAP7_75t_SL g3592 ( 
.A(n_3371),
.Y(n_3592)
);

AOI221xp5_ASAP7_75t_SL g3593 ( 
.A1(n_3085),
.A2(n_2569),
.B1(n_2570),
.B2(n_2558),
.C(n_2557),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_2894),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3409),
.B(n_2781),
.Y(n_3595)
);

AO31x2_ASAP7_75t_L g3596 ( 
.A1(n_3062),
.A2(n_2318),
.A3(n_2323),
.B(n_2314),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_SL g3597 ( 
.A(n_3313),
.B(n_3174),
.Y(n_3597)
);

AOI21xp5_ASAP7_75t_L g3598 ( 
.A1(n_2913),
.A2(n_2433),
.B(n_2687),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_2913),
.A2(n_2433),
.B(n_2687),
.Y(n_3599)
);

AO21x2_ASAP7_75t_L g3600 ( 
.A1(n_3217),
.A2(n_2228),
.B(n_2224),
.Y(n_3600)
);

NOR2xp33_ASAP7_75t_L g3601 ( 
.A(n_3186),
.B(n_2569),
.Y(n_3601)
);

AOI21xp5_ASAP7_75t_L g3602 ( 
.A1(n_2983),
.A2(n_2433),
.B(n_2687),
.Y(n_3602)
);

AOI211x1_ASAP7_75t_L g3603 ( 
.A1(n_3117),
.A2(n_2596),
.B(n_2599),
.C(n_2570),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3409),
.B(n_2784),
.Y(n_3604)
);

OAI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_2901),
.A2(n_2351),
.B(n_2311),
.Y(n_3605)
);

OAI22xp5_ASAP7_75t_L g3606 ( 
.A1(n_3325),
.A2(n_2596),
.B1(n_2642),
.B2(n_2599),
.Y(n_3606)
);

OR2x2_ASAP7_75t_L g3607 ( 
.A(n_3333),
.B(n_2345),
.Y(n_3607)
);

AND3x4_ASAP7_75t_L g3608 ( 
.A(n_3070),
.B(n_2813),
.C(n_2587),
.Y(n_3608)
);

NAND2xp33_ASAP7_75t_R g3609 ( 
.A(n_2845),
.B(n_2514),
.Y(n_3609)
);

NOR2xp33_ASAP7_75t_SL g3610 ( 
.A(n_2890),
.B(n_2633),
.Y(n_3610)
);

OAI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_2912),
.A2(n_2351),
.B(n_2311),
.Y(n_3611)
);

OAI22xp5_ASAP7_75t_L g3612 ( 
.A1(n_2849),
.A2(n_2642),
.B1(n_2668),
.B2(n_2667),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3413),
.B(n_2784),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_2894),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3413),
.B(n_2798),
.Y(n_3615)
);

OAI22xp5_ASAP7_75t_L g3616 ( 
.A1(n_2849),
.A2(n_2667),
.B1(n_2671),
.B2(n_2668),
.Y(n_3616)
);

NOR2x1_ASAP7_75t_SL g3617 ( 
.A(n_3374),
.B(n_2687),
.Y(n_3617)
);

AOI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_3056),
.A2(n_2433),
.B(n_2687),
.Y(n_3618)
);

OA21x2_ASAP7_75t_L g3619 ( 
.A1(n_3044),
.A2(n_2384),
.B(n_2185),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3415),
.B(n_2798),
.Y(n_3620)
);

AOI21xp33_ASAP7_75t_L g3621 ( 
.A1(n_3085),
.A2(n_2704),
.B(n_2643),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3415),
.B(n_2800),
.Y(n_3622)
);

AOI22xp5_ASAP7_75t_L g3623 ( 
.A1(n_2864),
.A2(n_2351),
.B1(n_2405),
.B2(n_2643),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_2904),
.Y(n_3624)
);

NAND3x1_ASAP7_75t_L g3625 ( 
.A(n_3359),
.B(n_2451),
.C(n_2477),
.Y(n_3625)
);

AO21x1_ASAP7_75t_L g3626 ( 
.A1(n_3319),
.A2(n_2801),
.B(n_2800),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3248),
.Y(n_3627)
);

AOI21x1_ASAP7_75t_L g3628 ( 
.A1(n_3052),
.A2(n_2776),
.B(n_2822),
.Y(n_3628)
);

AOI21xp5_ASAP7_75t_L g3629 ( 
.A1(n_3046),
.A2(n_2269),
.B(n_2268),
.Y(n_3629)
);

OA21x2_ASAP7_75t_L g3630 ( 
.A1(n_2970),
.A2(n_2384),
.B(n_2185),
.Y(n_3630)
);

AND2x4_ASAP7_75t_L g3631 ( 
.A(n_3182),
.B(n_2813),
.Y(n_3631)
);

NAND3xp33_ASAP7_75t_SL g3632 ( 
.A(n_2877),
.B(n_2777),
.C(n_2660),
.Y(n_3632)
);

AND2x2_ASAP7_75t_L g3633 ( 
.A(n_3356),
.B(n_2537),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3356),
.B(n_2537),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3420),
.B(n_2801),
.Y(n_3635)
);

OAI21x1_ASAP7_75t_L g3636 ( 
.A1(n_3442),
.A2(n_3118),
.B(n_3115),
.Y(n_3636)
);

INVx2_ASAP7_75t_L g3637 ( 
.A(n_3248),
.Y(n_3637)
);

OA22x2_ASAP7_75t_L g3638 ( 
.A1(n_3353),
.A2(n_2643),
.B1(n_2405),
.B2(n_2351),
.Y(n_3638)
);

AOI21x1_ASAP7_75t_L g3639 ( 
.A1(n_3052),
.A2(n_2776),
.B(n_2822),
.Y(n_3639)
);

NOR2xp33_ASAP7_75t_L g3640 ( 
.A(n_2910),
.B(n_2671),
.Y(n_3640)
);

INVx1_ASAP7_75t_SL g3641 ( 
.A(n_3392),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3248),
.Y(n_3642)
);

OAI21x1_ASAP7_75t_SL g3643 ( 
.A1(n_3079),
.A2(n_2680),
.B(n_2676),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3420),
.B(n_2805),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3257),
.Y(n_3645)
);

INVx4_ASAP7_75t_L g3646 ( 
.A(n_3365),
.Y(n_3646)
);

AND3x4_ASAP7_75t_L g3647 ( 
.A(n_2985),
.B(n_2587),
.C(n_2584),
.Y(n_3647)
);

CKINVDCx20_ASAP7_75t_R g3648 ( 
.A(n_2930),
.Y(n_3648)
);

OAI22xp5_ASAP7_75t_L g3649 ( 
.A1(n_2895),
.A2(n_2680),
.B1(n_2690),
.B2(n_2676),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3422),
.B(n_3428),
.Y(n_3650)
);

O2A1O1Ixp5_ASAP7_75t_L g3651 ( 
.A1(n_3124),
.A2(n_2470),
.B(n_2516),
.C(n_2413),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3422),
.B(n_2805),
.Y(n_3652)
);

INVx3_ASAP7_75t_L g3653 ( 
.A(n_3436),
.Y(n_3653)
);

AOI21x1_ASAP7_75t_L g3654 ( 
.A1(n_2851),
.A2(n_2822),
.B(n_2538),
.Y(n_3654)
);

AND2x4_ASAP7_75t_L g3655 ( 
.A(n_3182),
.B(n_2428),
.Y(n_3655)
);

OAI21xp5_ASAP7_75t_L g3656 ( 
.A1(n_2989),
.A2(n_2405),
.B(n_2643),
.Y(n_3656)
);

BUFx2_ASAP7_75t_R g3657 ( 
.A(n_3302),
.Y(n_3657)
);

INVx3_ASAP7_75t_L g3658 ( 
.A(n_3436),
.Y(n_3658)
);

BUFx8_ASAP7_75t_SL g3659 ( 
.A(n_3144),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3428),
.B(n_2810),
.Y(n_3660)
);

OAI22x1_ASAP7_75t_L g3661 ( 
.A1(n_3017),
.A2(n_2817),
.B1(n_2810),
.B2(n_2200),
.Y(n_3661)
);

AOI21x1_ASAP7_75t_L g3662 ( 
.A1(n_2851),
.A2(n_2822),
.B(n_2538),
.Y(n_3662)
);

INVx6_ASAP7_75t_SL g3663 ( 
.A(n_2968),
.Y(n_3663)
);

OAI21xp5_ASAP7_75t_L g3664 ( 
.A1(n_2981),
.A2(n_2815),
.B(n_2396),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3257),
.Y(n_3665)
);

AOI21xp5_ASAP7_75t_L g3666 ( 
.A1(n_3365),
.A2(n_2269),
.B(n_2268),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_2904),
.Y(n_3667)
);

OAI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_2937),
.A2(n_2815),
.B(n_2396),
.Y(n_3668)
);

INVx3_ASAP7_75t_L g3669 ( 
.A(n_2960),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3441),
.B(n_2817),
.Y(n_3670)
);

AOI21xp5_ASAP7_75t_L g3671 ( 
.A1(n_3365),
.A2(n_2843),
.B(n_3083),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3441),
.B(n_2477),
.Y(n_3672)
);

BUFx3_ASAP7_75t_L g3673 ( 
.A(n_3108),
.Y(n_3673)
);

INVx3_ASAP7_75t_L g3674 ( 
.A(n_2978),
.Y(n_3674)
);

OAI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_2882),
.A2(n_2918),
.B(n_2948),
.Y(n_3675)
);

AOI21xp5_ASAP7_75t_L g3676 ( 
.A1(n_3365),
.A2(n_2337),
.B(n_2269),
.Y(n_3676)
);

HB1xp67_ASAP7_75t_L g3677 ( 
.A(n_2906),
.Y(n_3677)
);

AND2x4_ASAP7_75t_L g3678 ( 
.A(n_3182),
.B(n_2428),
.Y(n_3678)
);

OR2x2_ASAP7_75t_L g3679 ( 
.A(n_3333),
.B(n_2345),
.Y(n_3679)
);

AND2x6_ASAP7_75t_L g3680 ( 
.A(n_3204),
.B(n_2194),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_2908),
.Y(n_3681)
);

INVx5_ASAP7_75t_L g3682 ( 
.A(n_3292),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_2928),
.B(n_2494),
.Y(n_3683)
);

OAI22xp5_ASAP7_75t_L g3684 ( 
.A1(n_2841),
.A2(n_2693),
.B1(n_2708),
.B2(n_2690),
.Y(n_3684)
);

A2O1A1Ixp33_ASAP7_75t_L g3685 ( 
.A1(n_2882),
.A2(n_2965),
.B(n_2979),
.C(n_2887),
.Y(n_3685)
);

OA21x2_ASAP7_75t_L g3686 ( 
.A1(n_2844),
.A2(n_2397),
.B(n_2386),
.Y(n_3686)
);

INVx3_ASAP7_75t_SL g3687 ( 
.A(n_3387),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_SL g3688 ( 
.A(n_2866),
.B(n_2633),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3410),
.B(n_3354),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3257),
.Y(n_3690)
);

AND2x4_ASAP7_75t_L g3691 ( 
.A(n_3204),
.B(n_2428),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_2908),
.Y(n_3692)
);

CKINVDCx20_ASAP7_75t_R g3693 ( 
.A(n_3147),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_2928),
.B(n_2494),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_2976),
.B(n_2510),
.Y(n_3695)
);

AO31x2_ASAP7_75t_L g3696 ( 
.A1(n_3181),
.A2(n_2323),
.A3(n_2328),
.B(n_2318),
.Y(n_3696)
);

OAI22xp33_ASAP7_75t_L g3697 ( 
.A1(n_3066),
.A2(n_2687),
.B1(n_2504),
.B2(n_2190),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_2976),
.B(n_2510),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_2977),
.B(n_2510),
.Y(n_3699)
);

NAND2x1p5_ASAP7_75t_L g3700 ( 
.A(n_3023),
.B(n_2194),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3401),
.A2(n_2361),
.B(n_2337),
.Y(n_3701)
);

OAI21xp5_ASAP7_75t_SL g3702 ( 
.A1(n_3017),
.A2(n_2771),
.B(n_2769),
.Y(n_3702)
);

INVx3_ASAP7_75t_L g3703 ( 
.A(n_2978),
.Y(n_3703)
);

INVx3_ASAP7_75t_L g3704 ( 
.A(n_2978),
.Y(n_3704)
);

O2A1O1Ixp5_ASAP7_75t_SL g3705 ( 
.A1(n_3080),
.A2(n_2516),
.B(n_2470),
.C(n_2401),
.Y(n_3705)
);

OAI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_2918),
.A2(n_2815),
.B(n_2377),
.Y(n_3706)
);

OAI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_2926),
.A2(n_2377),
.B(n_2693),
.Y(n_3707)
);

BUFx2_ASAP7_75t_R g3708 ( 
.A(n_3302),
.Y(n_3708)
);

NOR2xp67_ASAP7_75t_L g3709 ( 
.A(n_3349),
.B(n_2653),
.Y(n_3709)
);

AO31x2_ASAP7_75t_L g3710 ( 
.A1(n_3181),
.A2(n_2328),
.A3(n_2330),
.B(n_2323),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_SL g3711 ( 
.A(n_3348),
.B(n_2633),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3410),
.B(n_2537),
.Y(n_3712)
);

AOI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3073),
.A2(n_2721),
.B1(n_2769),
.B2(n_2633),
.Y(n_3713)
);

INVx1_ASAP7_75t_SL g3714 ( 
.A(n_3392),
.Y(n_3714)
);

NAND2x1_ASAP7_75t_L g3715 ( 
.A(n_3362),
.B(n_2605),
.Y(n_3715)
);

OAI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_2982),
.A2(n_2713),
.B(n_2708),
.Y(n_3716)
);

O2A1O1Ixp33_ASAP7_75t_SL g3717 ( 
.A1(n_3256),
.A2(n_3295),
.B(n_3244),
.C(n_3263),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_2977),
.B(n_2348),
.Y(n_3718)
);

AOI21x1_ASAP7_75t_L g3719 ( 
.A1(n_3432),
.A2(n_3433),
.B(n_2872),
.Y(n_3719)
);

OAI21x1_ASAP7_75t_L g3720 ( 
.A1(n_3398),
.A2(n_2548),
.B(n_2527),
.Y(n_3720)
);

INVx5_ASAP7_75t_L g3721 ( 
.A(n_3292),
.Y(n_3721)
);

AOI21x1_ASAP7_75t_L g3722 ( 
.A1(n_3101),
.A2(n_2538),
.B(n_2536),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3367),
.B(n_2354),
.Y(n_3723)
);

OAI22xp33_ASAP7_75t_L g3724 ( 
.A1(n_3066),
.A2(n_2687),
.B1(n_2504),
.B2(n_2190),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_2919),
.Y(n_3725)
);

INVx3_ASAP7_75t_L g3726 ( 
.A(n_2978),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3354),
.B(n_2537),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3367),
.B(n_2354),
.Y(n_3728)
);

OAI21x1_ASAP7_75t_L g3729 ( 
.A1(n_3398),
.A2(n_2548),
.B(n_2527),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_2919),
.Y(n_3730)
);

A2O1A1Ixp33_ASAP7_75t_L g3731 ( 
.A1(n_3027),
.A2(n_2714),
.B(n_2718),
.C(n_2713),
.Y(n_3731)
);

NOR2xp33_ASAP7_75t_L g3732 ( 
.A(n_2916),
.B(n_2714),
.Y(n_3732)
);

OAI22x1_ASAP7_75t_L g3733 ( 
.A1(n_3023),
.A2(n_2536),
.B1(n_2634),
.B2(n_2540),
.Y(n_3733)
);

BUFx6f_ASAP7_75t_L g3734 ( 
.A(n_2978),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_2920),
.Y(n_3735)
);

AOI21xp5_ASAP7_75t_L g3736 ( 
.A1(n_2993),
.A2(n_2361),
.B(n_2337),
.Y(n_3736)
);

AND2x4_ASAP7_75t_L g3737 ( 
.A(n_3204),
.B(n_2428),
.Y(n_3737)
);

AOI211x1_ASAP7_75t_L g3738 ( 
.A1(n_3399),
.A2(n_2726),
.B(n_2730),
.C(n_2718),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3355),
.B(n_2550),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_2955),
.B(n_3038),
.Y(n_3740)
);

INVx3_ASAP7_75t_L g3741 ( 
.A(n_2978),
.Y(n_3741)
);

AOI221xp5_ASAP7_75t_SL g3742 ( 
.A1(n_3195),
.A2(n_2730),
.B1(n_2726),
.B2(n_2740),
.C(n_2767),
.Y(n_3742)
);

CKINVDCx5p33_ASAP7_75t_R g3743 ( 
.A(n_3098),
.Y(n_3743)
);

OAI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_3437),
.A2(n_2752),
.B1(n_2755),
.B2(n_2740),
.Y(n_3744)
);

OAI21x1_ASAP7_75t_L g3745 ( 
.A1(n_3258),
.A2(n_2548),
.B(n_2527),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_2920),
.Y(n_3746)
);

OA21x2_ASAP7_75t_L g3747 ( 
.A1(n_2844),
.A2(n_2397),
.B(n_2386),
.Y(n_3747)
);

CKINVDCx11_ASAP7_75t_R g3748 ( 
.A(n_3153),
.Y(n_3748)
);

INVx3_ASAP7_75t_L g3749 ( 
.A(n_2980),
.Y(n_3749)
);

CKINVDCx20_ASAP7_75t_R g3750 ( 
.A(n_3051),
.Y(n_3750)
);

AND2x4_ASAP7_75t_L g3751 ( 
.A(n_3204),
.B(n_2428),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_3265),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_2955),
.B(n_2355),
.Y(n_3753)
);

INVx2_ASAP7_75t_SL g3754 ( 
.A(n_3071),
.Y(n_3754)
);

AOI21x1_ASAP7_75t_L g3755 ( 
.A1(n_3116),
.A2(n_2880),
.B(n_3165),
.Y(n_3755)
);

AOI21x1_ASAP7_75t_L g3756 ( 
.A1(n_3262),
.A2(n_2540),
.B(n_2536),
.Y(n_3756)
);

BUFx2_ASAP7_75t_R g3757 ( 
.A(n_3060),
.Y(n_3757)
);

AOI22xp33_ASAP7_75t_SL g3758 ( 
.A1(n_2917),
.A2(n_2514),
.B1(n_2633),
.B2(n_2504),
.Y(n_3758)
);

BUFx6f_ASAP7_75t_L g3759 ( 
.A(n_2980),
.Y(n_3759)
);

AND2x2_ASAP7_75t_L g3760 ( 
.A(n_3355),
.B(n_2550),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3265),
.Y(n_3761)
);

AOI21xp5_ASAP7_75t_L g3762 ( 
.A1(n_2890),
.A2(n_3097),
.B(n_2958),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3038),
.B(n_2355),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_L g3764 ( 
.A(n_2909),
.B(n_2752),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_2945),
.Y(n_3765)
);

INVx3_ASAP7_75t_L g3766 ( 
.A(n_2980),
.Y(n_3766)
);

OR2x2_ASAP7_75t_L g3767 ( 
.A(n_3350),
.B(n_2368),
.Y(n_3767)
);

OA21x2_ASAP7_75t_L g3768 ( 
.A1(n_2858),
.A2(n_2397),
.B(n_2386),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3110),
.B(n_2368),
.Y(n_3769)
);

AOI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_2958),
.A2(n_2640),
.B(n_2634),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3110),
.B(n_2369),
.Y(n_3771)
);

OAI21x1_ASAP7_75t_L g3772 ( 
.A1(n_3340),
.A2(n_2581),
.B(n_2552),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3097),
.A2(n_2685),
.B(n_2640),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3200),
.B(n_2369),
.Y(n_3774)
);

INVx2_ASAP7_75t_SL g3775 ( 
.A(n_3152),
.Y(n_3775)
);

OAI21x1_ASAP7_75t_L g3776 ( 
.A1(n_3341),
.A2(n_2581),
.B(n_2552),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3200),
.B(n_2721),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3005),
.A2(n_2361),
.B(n_2337),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_2945),
.Y(n_3779)
);

AOI21xp5_ASAP7_75t_L g3780 ( 
.A1(n_3090),
.A2(n_3034),
.B(n_3020),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3265),
.Y(n_3781)
);

NOR2xp67_ASAP7_75t_L g3782 ( 
.A(n_3349),
.B(n_2653),
.Y(n_3782)
);

OAI21x1_ASAP7_75t_L g3783 ( 
.A1(n_3341),
.A2(n_2581),
.B(n_2552),
.Y(n_3783)
);

OAI21xp5_ASAP7_75t_L g3784 ( 
.A1(n_2952),
.A2(n_2762),
.B(n_2755),
.Y(n_3784)
);

OA21x2_ASAP7_75t_L g3785 ( 
.A1(n_3224),
.A2(n_2492),
.B(n_2491),
.Y(n_3785)
);

O2A1O1Ixp5_ASAP7_75t_L g3786 ( 
.A1(n_3183),
.A2(n_2587),
.B(n_2624),
.C(n_2584),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_2925),
.B(n_2867),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_2925),
.B(n_2769),
.Y(n_3788)
);

NAND3xp33_ASAP7_75t_L g3789 ( 
.A(n_2943),
.B(n_2767),
.C(n_2762),
.Y(n_3789)
);

AOI211x1_ASAP7_75t_L g3790 ( 
.A1(n_3384),
.A2(n_2492),
.B(n_2546),
.C(n_2491),
.Y(n_3790)
);

BUFx10_ASAP7_75t_L g3791 ( 
.A(n_3362),
.Y(n_3791)
);

OAI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_2885),
.A2(n_2685),
.B(n_2640),
.Y(n_3792)
);

AND2x4_ASAP7_75t_L g3793 ( 
.A(n_3227),
.B(n_3380),
.Y(n_3793)
);

AND3x4_ASAP7_75t_L g3794 ( 
.A(n_3289),
.B(n_2587),
.C(n_2584),
.Y(n_3794)
);

OAI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_2898),
.A2(n_2688),
.B(n_2685),
.Y(n_3795)
);

CKINVDCx20_ASAP7_75t_R g3796 ( 
.A(n_3345),
.Y(n_3796)
);

AOI21xp5_ASAP7_75t_L g3797 ( 
.A1(n_3055),
.A2(n_3078),
.B(n_3440),
.Y(n_3797)
);

HB1xp67_ASAP7_75t_L g3798 ( 
.A(n_3164),
.Y(n_3798)
);

HB1xp67_ASAP7_75t_L g3799 ( 
.A(n_3239),
.Y(n_3799)
);

AOI21xp33_ASAP7_75t_L g3800 ( 
.A1(n_3353),
.A2(n_2673),
.B(n_2663),
.Y(n_3800)
);

BUFx2_ASAP7_75t_SL g3801 ( 
.A(n_3364),
.Y(n_3801)
);

O2A1O1Ixp5_ASAP7_75t_L g3802 ( 
.A1(n_3210),
.A2(n_2584),
.B(n_2624),
.C(n_2587),
.Y(n_3802)
);

CKINVDCx20_ASAP7_75t_R g3803 ( 
.A(n_3250),
.Y(n_3803)
);

AOI21xp5_ASAP7_75t_L g3804 ( 
.A1(n_3440),
.A2(n_2361),
.B(n_2337),
.Y(n_3804)
);

O2A1O1Ixp33_ASAP7_75t_SL g3805 ( 
.A1(n_3021),
.A2(n_2666),
.B(n_2710),
.C(n_2588),
.Y(n_3805)
);

AOI21xp5_ASAP7_75t_L g3806 ( 
.A1(n_3229),
.A2(n_2361),
.B(n_2337),
.Y(n_3806)
);

AOI221xp5_ASAP7_75t_SL g3807 ( 
.A1(n_3425),
.A2(n_2688),
.B1(n_2727),
.B2(n_2837),
.C(n_2738),
.Y(n_3807)
);

OAI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3104),
.A2(n_3224),
.B(n_3150),
.Y(n_3808)
);

NOR2xp33_ASAP7_75t_L g3809 ( 
.A(n_2939),
.B(n_2659),
.Y(n_3809)
);

AOI21xp5_ASAP7_75t_SL g3810 ( 
.A1(n_3196),
.A2(n_2745),
.B(n_2205),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_2869),
.B(n_2663),
.Y(n_3811)
);

OAI21xp5_ASAP7_75t_L g3812 ( 
.A1(n_3260),
.A2(n_2727),
.B(n_2688),
.Y(n_3812)
);

A2O1A1Ixp33_ASAP7_75t_L g3813 ( 
.A1(n_2917),
.A2(n_2727),
.B(n_2502),
.C(n_2428),
.Y(n_3813)
);

O2A1O1Ixp5_ASAP7_75t_L g3814 ( 
.A1(n_3298),
.A2(n_2584),
.B(n_2629),
.C(n_2624),
.Y(n_3814)
);

AND2x6_ASAP7_75t_L g3815 ( 
.A(n_3033),
.B(n_2194),
.Y(n_3815)
);

OA21x2_ASAP7_75t_L g3816 ( 
.A1(n_3222),
.A2(n_2492),
.B(n_2491),
.Y(n_3816)
);

AOI22xp5_ASAP7_75t_L g3817 ( 
.A1(n_3073),
.A2(n_2633),
.B1(n_2190),
.B2(n_2745),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_2879),
.B(n_2673),
.Y(n_3818)
);

BUFx3_ASAP7_75t_L g3819 ( 
.A(n_3108),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_2879),
.B(n_2691),
.Y(n_3820)
);

OAI21xp5_ASAP7_75t_L g3821 ( 
.A1(n_3133),
.A2(n_2387),
.B(n_2310),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_2883),
.B(n_2691),
.Y(n_3822)
);

OAI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3133),
.A2(n_2387),
.B(n_2310),
.Y(n_3823)
);

OAI21x1_ASAP7_75t_SL g3824 ( 
.A1(n_3072),
.A2(n_2772),
.B(n_2701),
.Y(n_3824)
);

AO31x2_ASAP7_75t_L g3825 ( 
.A1(n_2954),
.A2(n_2374),
.A3(n_2380),
.B(n_2356),
.Y(n_3825)
);

CKINVDCx20_ASAP7_75t_R g3826 ( 
.A(n_3312),
.Y(n_3826)
);

BUFx2_ASAP7_75t_L g3827 ( 
.A(n_3109),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3229),
.A2(n_2379),
.B(n_2361),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_2963),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3266),
.Y(n_3830)
);

AOI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_3075),
.A2(n_2379),
.B(n_2361),
.Y(n_3831)
);

BUFx2_ASAP7_75t_L g3832 ( 
.A(n_3109),
.Y(n_3832)
);

OAI21xp33_ASAP7_75t_L g3833 ( 
.A1(n_3088),
.A2(n_2550),
.B(n_2560),
.Y(n_3833)
);

O2A1O1Ixp33_ASAP7_75t_SL g3834 ( 
.A1(n_3389),
.A2(n_2739),
.B(n_2754),
.C(n_2716),
.Y(n_3834)
);

AOI22xp5_ASAP7_75t_L g3835 ( 
.A1(n_2917),
.A2(n_2633),
.B1(n_2190),
.B2(n_2745),
.Y(n_3835)
);

CKINVDCx11_ASAP7_75t_R g3836 ( 
.A(n_3234),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_2883),
.B(n_2716),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_3076),
.A2(n_2382),
.B(n_2379),
.Y(n_3838)
);

A2O1A1Ixp33_ASAP7_75t_L g3839 ( 
.A1(n_3121),
.A2(n_2502),
.B(n_2205),
.C(n_2210),
.Y(n_3839)
);

OAI22xp5_ASAP7_75t_L g3840 ( 
.A1(n_3066),
.A2(n_2550),
.B1(n_2745),
.B2(n_2560),
.Y(n_3840)
);

AO31x2_ASAP7_75t_L g3841 ( 
.A1(n_2954),
.A2(n_2380),
.A3(n_2383),
.B(n_2374),
.Y(n_3841)
);

BUFx2_ASAP7_75t_L g3842 ( 
.A(n_3119),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_2966),
.Y(n_3843)
);

INVx3_ASAP7_75t_L g3844 ( 
.A(n_2980),
.Y(n_3844)
);

OAI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3337),
.A2(n_2550),
.B1(n_2745),
.B2(n_2560),
.Y(n_3845)
);

NAND2x1_ASAP7_75t_L g3846 ( 
.A(n_3362),
.B(n_2605),
.Y(n_3846)
);

BUFx2_ASAP7_75t_L g3847 ( 
.A(n_3119),
.Y(n_3847)
);

NOR2xp33_ASAP7_75t_R g3848 ( 
.A(n_3417),
.B(n_2580),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_SL g3849 ( 
.A(n_3192),
.B(n_2624),
.Y(n_3849)
);

CKINVDCx11_ASAP7_75t_R g3850 ( 
.A(n_3234),
.Y(n_3850)
);

HB1xp67_ASAP7_75t_L g3851 ( 
.A(n_3264),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_2966),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_2974),
.Y(n_3853)
);

OAI21xp33_ASAP7_75t_L g3854 ( 
.A1(n_3161),
.A2(n_2550),
.B(n_2560),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_SL g3855 ( 
.A(n_3192),
.B(n_2624),
.Y(n_3855)
);

AND2x4_ASAP7_75t_L g3856 ( 
.A(n_3227),
.B(n_2560),
.Y(n_3856)
);

NAND3xp33_ASAP7_75t_L g3857 ( 
.A(n_3105),
.B(n_3067),
.C(n_2907),
.Y(n_3857)
);

AND2x2_ASAP7_75t_L g3858 ( 
.A(n_3363),
.B(n_2560),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_2974),
.Y(n_3859)
);

BUFx3_ASAP7_75t_L g3860 ( 
.A(n_3108),
.Y(n_3860)
);

AOI221xp5_ASAP7_75t_L g3861 ( 
.A1(n_3158),
.A2(n_2422),
.B1(n_2455),
.B2(n_2454),
.C(n_2542),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_2984),
.Y(n_3862)
);

AOI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3383),
.A2(n_3061),
.B(n_3059),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3266),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_2900),
.B(n_2754),
.Y(n_3865)
);

CKINVDCx20_ASAP7_75t_R g3866 ( 
.A(n_3336),
.Y(n_3866)
);

OAI21xp5_ASAP7_75t_SL g3867 ( 
.A1(n_3342),
.A2(n_3347),
.B(n_2973),
.Y(n_3867)
);

OAI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3254),
.A2(n_2387),
.B(n_2310),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_2907),
.B(n_2760),
.Y(n_3869)
);

INVx2_ASAP7_75t_L g3870 ( 
.A(n_3266),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_2984),
.Y(n_3871)
);

OR2x2_ASAP7_75t_L g3872 ( 
.A(n_3350),
.B(n_2760),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_2914),
.B(n_2736),
.Y(n_3873)
);

OAI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3077),
.A2(n_3253),
.B(n_3273),
.Y(n_3874)
);

OAI21xp5_ASAP7_75t_SL g3875 ( 
.A1(n_2973),
.A2(n_2629),
.B(n_2659),
.Y(n_3875)
);

AOI21xp5_ASAP7_75t_L g3876 ( 
.A1(n_3307),
.A2(n_2382),
.B(n_2379),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_2914),
.B(n_2736),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_3016),
.B(n_2736),
.Y(n_3878)
);

AOI21x1_ASAP7_75t_L g3879 ( 
.A1(n_3320),
.A2(n_2629),
.B(n_2289),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3016),
.B(n_2736),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_SL g3881 ( 
.A1(n_3125),
.A2(n_2745),
.B(n_2205),
.Y(n_3881)
);

OAI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3077),
.A2(n_2387),
.B(n_2310),
.Y(n_3882)
);

NOR2xp67_ASAP7_75t_SL g3883 ( 
.A(n_3283),
.B(n_2425),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_2992),
.Y(n_3884)
);

NOR2xp33_ASAP7_75t_R g3885 ( 
.A(n_3246),
.B(n_2580),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_3270),
.Y(n_3886)
);

BUFx6f_ASAP7_75t_L g3887 ( 
.A(n_2980),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_2992),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3018),
.B(n_2736),
.Y(n_3889)
);

AOI21xp5_ASAP7_75t_L g3890 ( 
.A1(n_3307),
.A2(n_2382),
.B(n_2379),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_SL g3891 ( 
.A(n_3192),
.B(n_2629),
.Y(n_3891)
);

OAI22xp5_ASAP7_75t_L g3892 ( 
.A1(n_3338),
.A2(n_2745),
.B1(n_2683),
.B2(n_2659),
.Y(n_3892)
);

A2O1A1Ixp33_ASAP7_75t_L g3893 ( 
.A1(n_3148),
.A2(n_2502),
.B(n_2194),
.C(n_2205),
.Y(n_3893)
);

AOI21x1_ASAP7_75t_L g3894 ( 
.A1(n_3330),
.A2(n_2629),
.B(n_2289),
.Y(n_3894)
);

OA21x2_ASAP7_75t_L g3895 ( 
.A1(n_3230),
.A2(n_2578),
.B(n_2577),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3270),
.Y(n_3896)
);

AND2x4_ASAP7_75t_L g3897 ( 
.A(n_3227),
.B(n_2194),
.Y(n_3897)
);

AOI21xp5_ASAP7_75t_L g3898 ( 
.A1(n_3307),
.A2(n_2382),
.B(n_2379),
.Y(n_3898)
);

OA21x2_ASAP7_75t_L g3899 ( 
.A1(n_3232),
.A2(n_2578),
.B(n_2577),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3018),
.B(n_2736),
.Y(n_3900)
);

AO22x2_ASAP7_75t_L g3901 ( 
.A1(n_3314),
.A2(n_2444),
.B1(n_2422),
.B2(n_2542),
.Y(n_3901)
);

AO21x1_ASAP7_75t_L g3902 ( 
.A1(n_2942),
.A2(n_2669),
.B(n_2659),
.Y(n_3902)
);

BUFx6f_ASAP7_75t_L g3903 ( 
.A(n_2994),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3026),
.B(n_2736),
.Y(n_3904)
);

BUFx3_ASAP7_75t_L g3905 ( 
.A(n_3283),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3026),
.B(n_3030),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3030),
.B(n_3037),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_SL g3908 ( 
.A(n_3192),
.B(n_3373),
.Y(n_3908)
);

INVx3_ASAP7_75t_SL g3909 ( 
.A(n_3387),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_3270),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3037),
.B(n_2736),
.Y(n_3911)
);

OAI21xp5_ASAP7_75t_L g3912 ( 
.A1(n_3111),
.A2(n_2387),
.B(n_2310),
.Y(n_3912)
);

AOI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_3307),
.A2(n_2408),
.B(n_2382),
.Y(n_3913)
);

O2A1O1Ixp33_ASAP7_75t_SL g3914 ( 
.A1(n_3180),
.A2(n_2660),
.B(n_2803),
.C(n_2777),
.Y(n_3914)
);

INVx2_ASAP7_75t_SL g3915 ( 
.A(n_3276),
.Y(n_3915)
);

NOR2xp33_ASAP7_75t_L g3916 ( 
.A(n_3031),
.B(n_2659),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_SL g3917 ( 
.A(n_3373),
.B(n_2659),
.Y(n_3917)
);

OR2x2_ASAP7_75t_L g3918 ( 
.A(n_3406),
.B(n_2498),
.Y(n_3918)
);

INVx2_ASAP7_75t_SL g3919 ( 
.A(n_3142),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_2995),
.Y(n_3920)
);

O2A1O1Ixp5_ASAP7_75t_L g3921 ( 
.A1(n_3282),
.A2(n_2597),
.B(n_2528),
.C(n_2689),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_2995),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3040),
.B(n_2738),
.Y(n_3923)
);

INVx2_ASAP7_75t_SL g3924 ( 
.A(n_3142),
.Y(n_3924)
);

A2O1A1Ixp33_ASAP7_75t_L g3925 ( 
.A1(n_3149),
.A2(n_3160),
.B(n_3314),
.C(n_2969),
.Y(n_3925)
);

AOI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3307),
.A2(n_2408),
.B(n_2701),
.Y(n_3926)
);

OAI21xp5_ASAP7_75t_L g3927 ( 
.A1(n_3205),
.A2(n_2387),
.B(n_2310),
.Y(n_3927)
);

AOI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_3170),
.A2(n_2289),
.B(n_2276),
.Y(n_3928)
);

AND2x4_ASAP7_75t_L g3929 ( 
.A(n_3227),
.B(n_2205),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3040),
.B(n_3041),
.Y(n_3930)
);

BUFx3_ASAP7_75t_L g3931 ( 
.A(n_3283),
.Y(n_3931)
);

CKINVDCx20_ASAP7_75t_R g3932 ( 
.A(n_3357),
.Y(n_3932)
);

OAI22xp5_ASAP7_75t_L g3933 ( 
.A1(n_3344),
.A2(n_2669),
.B1(n_2683),
.B2(n_2732),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_2998),
.Y(n_3934)
);

AOI21xp5_ASAP7_75t_SL g3935 ( 
.A1(n_2859),
.A2(n_2275),
.B(n_2210),
.Y(n_3935)
);

NOR2xp33_ASAP7_75t_L g3936 ( 
.A(n_3404),
.B(n_2669),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_3041),
.B(n_2738),
.Y(n_3937)
);

AO21x2_ASAP7_75t_L g3938 ( 
.A1(n_3275),
.A2(n_2228),
.B(n_2224),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3042),
.B(n_2738),
.Y(n_3939)
);

AOI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_2994),
.A2(n_2408),
.B(n_2701),
.Y(n_3940)
);

AOI21xp33_ASAP7_75t_L g3941 ( 
.A1(n_3267),
.A2(n_2250),
.B(n_2229),
.Y(n_3941)
);

BUFx3_ASAP7_75t_L g3942 ( 
.A(n_3332),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3042),
.B(n_2738),
.Y(n_3943)
);

NOR2xp67_ASAP7_75t_L g3944 ( 
.A(n_3349),
.B(n_2653),
.Y(n_3944)
);

O2A1O1Ixp33_ASAP7_75t_SL g3945 ( 
.A1(n_3091),
.A2(n_2803),
.B(n_2823),
.C(n_2804),
.Y(n_3945)
);

AOI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_3376),
.A2(n_2290),
.B(n_2276),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_2998),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3000),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3000),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3047),
.B(n_2738),
.Y(n_3950)
);

INVx3_ASAP7_75t_L g3951 ( 
.A(n_2994),
.Y(n_3951)
);

AOI21xp5_ASAP7_75t_L g3952 ( 
.A1(n_2994),
.A2(n_2408),
.B(n_2772),
.Y(n_3952)
);

BUFx10_ASAP7_75t_L g3953 ( 
.A(n_3362),
.Y(n_3953)
);

INVx2_ASAP7_75t_SL g3954 ( 
.A(n_3221),
.Y(n_3954)
);

NAND3xp33_ASAP7_75t_SL g3955 ( 
.A(n_2868),
.B(n_2956),
.C(n_2951),
.Y(n_3955)
);

NOR2xp33_ASAP7_75t_L g3956 ( 
.A(n_3414),
.B(n_2669),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3002),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3047),
.B(n_3063),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3063),
.B(n_2738),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_SL g3960 ( 
.A(n_3293),
.B(n_2669),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3068),
.B(n_2738),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3068),
.B(n_2837),
.Y(n_3962)
);

INVx1_ASAP7_75t_SL g3963 ( 
.A(n_3131),
.Y(n_3963)
);

CKINVDCx5p33_ASAP7_75t_R g3964 ( 
.A(n_3332),
.Y(n_3964)
);

AOI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_2994),
.A2(n_2408),
.B(n_2772),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3074),
.B(n_2837),
.Y(n_3966)
);

A2O1A1Ixp33_ASAP7_75t_L g3967 ( 
.A1(n_3023),
.A2(n_2210),
.B(n_2275),
.C(n_2732),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3002),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3074),
.B(n_2837),
.Y(n_3969)
);

INVx3_ASAP7_75t_L g3970 ( 
.A(n_2994),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_2942),
.B(n_2837),
.Y(n_3971)
);

AOI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_3003),
.A2(n_2408),
.B(n_2772),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3003),
.A2(n_2408),
.B(n_2791),
.Y(n_3973)
);

OAI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3281),
.A2(n_2387),
.B(n_2310),
.Y(n_3974)
);

AND2x6_ASAP7_75t_L g3975 ( 
.A(n_3033),
.B(n_2210),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3291),
.Y(n_3976)
);

INVx1_ASAP7_75t_SL g3977 ( 
.A(n_3131),
.Y(n_3977)
);

OAI22xp5_ASAP7_75t_L g3978 ( 
.A1(n_3402),
.A2(n_2683),
.B1(n_2669),
.B2(n_2689),
.Y(n_3978)
);

A2O1A1Ixp33_ASAP7_75t_L g3979 ( 
.A1(n_3023),
.A2(n_2210),
.B(n_2275),
.C(n_2683),
.Y(n_3979)
);

OAI21xp5_ASAP7_75t_L g3980 ( 
.A1(n_3281),
.A2(n_2605),
.B(n_2364),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_SL g3981 ( 
.A(n_3300),
.B(n_2683),
.Y(n_3981)
);

OAI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3158),
.A2(n_2605),
.B(n_2364),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_3003),
.A2(n_2807),
.B(n_2791),
.Y(n_3983)
);

O2A1O1Ixp33_ASAP7_75t_SL g3984 ( 
.A1(n_3216),
.A2(n_2823),
.B(n_2804),
.C(n_2250),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_2949),
.B(n_2837),
.Y(n_3985)
);

INVx2_ASAP7_75t_SL g3986 ( 
.A(n_3316),
.Y(n_3986)
);

O2A1O1Ixp5_ASAP7_75t_L g3987 ( 
.A1(n_3391),
.A2(n_2528),
.B(n_2683),
.C(n_2689),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_3291),
.Y(n_3988)
);

AOI21x1_ASAP7_75t_L g3989 ( 
.A1(n_3418),
.A2(n_2317),
.B(n_2290),
.Y(n_3989)
);

BUFx12f_ASAP7_75t_L g3990 ( 
.A(n_3332),
.Y(n_3990)
);

AOI21xp5_ASAP7_75t_L g3991 ( 
.A1(n_3003),
.A2(n_2807),
.B(n_2791),
.Y(n_3991)
);

AND2x2_ASAP7_75t_L g3992 ( 
.A(n_3363),
.B(n_2504),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_2949),
.B(n_2953),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3006),
.Y(n_3994)
);

BUFx3_ASAP7_75t_L g3995 ( 
.A(n_3483),
.Y(n_3995)
);

AOI22xp33_ASAP7_75t_L g3996 ( 
.A1(n_3520),
.A2(n_3517),
.B1(n_3486),
.B2(n_3541),
.Y(n_3996)
);

OAI22xp5_ASAP7_75t_L g3997 ( 
.A1(n_3685),
.A2(n_2862),
.B1(n_2922),
.B2(n_2903),
.Y(n_3997)
);

OAI22xp5_ASAP7_75t_L g3998 ( 
.A1(n_3504),
.A2(n_2862),
.B1(n_3171),
.B2(n_3103),
.Y(n_3998)
);

OA21x2_ASAP7_75t_L g3999 ( 
.A1(n_3450),
.A2(n_3351),
.B(n_3323),
.Y(n_3999)
);

AOI22xp33_ASAP7_75t_L g4000 ( 
.A1(n_3520),
.A2(n_3517),
.B1(n_3486),
.B2(n_3541),
.Y(n_4000)
);

O2A1O1Ixp33_ASAP7_75t_L g4001 ( 
.A1(n_3524),
.A2(n_2936),
.B(n_2931),
.C(n_2953),
.Y(n_4001)
);

O2A1O1Ixp33_ASAP7_75t_L g4002 ( 
.A1(n_3675),
.A2(n_2971),
.B(n_3107),
.C(n_3106),
.Y(n_4002)
);

O2A1O1Ixp33_ASAP7_75t_SL g4003 ( 
.A1(n_3796),
.A2(n_3379),
.B(n_3424),
.C(n_3004),
.Y(n_4003)
);

INVx2_ASAP7_75t_SL g4004 ( 
.A(n_3793),
.Y(n_4004)
);

NOR2xp33_ASAP7_75t_SL g4005 ( 
.A(n_3495),
.B(n_3377),
.Y(n_4005)
);

AO31x2_ASAP7_75t_L g4006 ( 
.A1(n_3626),
.A2(n_3323),
.A3(n_3390),
.B(n_3351),
.Y(n_4006)
);

OAI221xp5_ASAP7_75t_L g4007 ( 
.A1(n_3675),
.A2(n_2934),
.B1(n_2940),
.B2(n_2935),
.C(n_2971),
.Y(n_4007)
);

AO31x2_ASAP7_75t_L g4008 ( 
.A1(n_3626),
.A2(n_3390),
.A3(n_3419),
.B(n_3416),
.Y(n_4008)
);

NOR2xp33_ASAP7_75t_SL g4009 ( 
.A(n_3657),
.B(n_3377),
.Y(n_4009)
);

OAI22xp33_ASAP7_75t_L g4010 ( 
.A1(n_3713),
.A2(n_2862),
.B1(n_3023),
.B2(n_3277),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3463),
.Y(n_4011)
);

BUFx3_ASAP7_75t_L g4012 ( 
.A(n_3483),
.Y(n_4012)
);

AO31x2_ASAP7_75t_L g4013 ( 
.A1(n_3547),
.A2(n_3318),
.A3(n_3305),
.B(n_3308),
.Y(n_4013)
);

O2A1O1Ixp33_ASAP7_75t_L g4014 ( 
.A1(n_3650),
.A2(n_2997),
.B(n_3001),
.C(n_2991),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3505),
.Y(n_4015)
);

O2A1O1Ixp33_ASAP7_75t_SL g4016 ( 
.A1(n_3750),
.A2(n_3932),
.B(n_3650),
.C(n_3693),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3689),
.B(n_3418),
.Y(n_4017)
);

O2A1O1Ixp33_ASAP7_75t_SL g4018 ( 
.A1(n_3648),
.A2(n_3009),
.B(n_3019),
.C(n_3007),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3503),
.B(n_3411),
.Y(n_4019)
);

AOI21xp5_ASAP7_75t_L g4020 ( 
.A1(n_3671),
.A2(n_3215),
.B(n_3228),
.Y(n_4020)
);

BUFx3_ASAP7_75t_L g4021 ( 
.A(n_3483),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3505),
.Y(n_4022)
);

NAND3x1_ASAP7_75t_L g4023 ( 
.A(n_3706),
.B(n_3423),
.C(n_3411),
.Y(n_4023)
);

O2A1O1Ixp33_ASAP7_75t_L g4024 ( 
.A1(n_3874),
.A2(n_3542),
.B(n_3451),
.C(n_3606),
.Y(n_4024)
);

INVx2_ASAP7_75t_SL g4025 ( 
.A(n_3793),
.Y(n_4025)
);

O2A1O1Ixp33_ASAP7_75t_SL g4026 ( 
.A1(n_3455),
.A2(n_3406),
.B(n_3408),
.C(n_3405),
.Y(n_4026)
);

OAI21xp5_ASAP7_75t_L g4027 ( 
.A1(n_3874),
.A2(n_2935),
.B(n_2934),
.Y(n_4027)
);

AO21x1_ASAP7_75t_L g4028 ( 
.A1(n_3547),
.A2(n_2997),
.B(n_2991),
.Y(n_4028)
);

AOI21xp5_ASAP7_75t_L g4029 ( 
.A1(n_3671),
.A2(n_3010),
.B(n_3001),
.Y(n_4029)
);

A2O1A1Ixp33_ASAP7_75t_L g4030 ( 
.A1(n_3867),
.A2(n_3431),
.B(n_3277),
.C(n_3360),
.Y(n_4030)
);

NOR2xp33_ASAP7_75t_L g4031 ( 
.A(n_3659),
.B(n_3423),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3503),
.B(n_3430),
.Y(n_4032)
);

OA21x2_ASAP7_75t_L g4033 ( 
.A1(n_3807),
.A2(n_3315),
.B(n_2896),
.Y(n_4033)
);

HB1xp67_ASAP7_75t_L g4034 ( 
.A(n_3986),
.Y(n_4034)
);

OAI22x1_ASAP7_75t_L g4035 ( 
.A1(n_3608),
.A2(n_3360),
.B1(n_3349),
.B2(n_3435),
.Y(n_4035)
);

AO31x2_ASAP7_75t_L g4036 ( 
.A1(n_3661),
.A2(n_3305),
.A3(n_3308),
.B(n_3291),
.Y(n_4036)
);

NAND2x1p5_ASAP7_75t_L g4037 ( 
.A(n_3587),
.B(n_3349),
.Y(n_4037)
);

BUFx6f_ASAP7_75t_L g4038 ( 
.A(n_3481),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3742),
.B(n_3993),
.Y(n_4039)
);

CKINVDCx20_ASAP7_75t_R g4040 ( 
.A(n_3748),
.Y(n_4040)
);

BUFx8_ASAP7_75t_L g4041 ( 
.A(n_3990),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3507),
.Y(n_4042)
);

AOI21xp5_ASAP7_75t_L g4043 ( 
.A1(n_3762),
.A2(n_3834),
.B(n_3805),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_3742),
.B(n_3430),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3463),
.Y(n_4045)
);

AND2x4_ASAP7_75t_L g4046 ( 
.A(n_3793),
.B(n_3360),
.Y(n_4046)
);

AND2x4_ASAP7_75t_L g4047 ( 
.A(n_3793),
.B(n_3360),
.Y(n_4047)
);

NAND3xp33_ASAP7_75t_SL g4048 ( 
.A(n_3867),
.B(n_3010),
.C(n_3086),
.Y(n_4048)
);

AOI22xp5_ASAP7_75t_L g4049 ( 
.A1(n_3606),
.A2(n_3431),
.B1(n_3127),
.B2(n_3197),
.Y(n_4049)
);

OAI22xp5_ASAP7_75t_L g4050 ( 
.A1(n_3504),
.A2(n_3039),
.B1(n_3057),
.B2(n_3036),
.Y(n_4050)
);

CKINVDCx5p33_ASAP7_75t_R g4051 ( 
.A(n_3476),
.Y(n_4051)
);

BUFx2_ASAP7_75t_R g4052 ( 
.A(n_3500),
.Y(n_4052)
);

OAI21xp5_ASAP7_75t_L g4053 ( 
.A1(n_3857),
.A2(n_2940),
.B(n_3122),
.Y(n_4053)
);

AOI21xp5_ASAP7_75t_L g4054 ( 
.A1(n_3863),
.A2(n_3126),
.B(n_3122),
.Y(n_4054)
);

NAND2x1p5_ASAP7_75t_L g4055 ( 
.A(n_3587),
.B(n_3360),
.Y(n_4055)
);

AO31x2_ASAP7_75t_L g4056 ( 
.A1(n_3661),
.A2(n_3308),
.A3(n_3317),
.B(n_3305),
.Y(n_4056)
);

OAI21x1_ASAP7_75t_L g4057 ( 
.A1(n_3705),
.A2(n_2891),
.B(n_2863),
.Y(n_4057)
);

INVx2_ASAP7_75t_SL g4058 ( 
.A(n_3754),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3993),
.B(n_3434),
.Y(n_4059)
);

NOR2xp33_ASAP7_75t_L g4060 ( 
.A(n_3757),
.B(n_3434),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3507),
.Y(n_4061)
);

O2A1O1Ixp33_ASAP7_75t_SL g4062 ( 
.A1(n_3803),
.A2(n_3408),
.B(n_3405),
.C(n_3065),
.Y(n_4062)
);

BUFx6f_ASAP7_75t_L g4063 ( 
.A(n_3481),
.Y(n_4063)
);

BUFx12f_ASAP7_75t_L g4064 ( 
.A(n_3743),
.Y(n_4064)
);

CKINVDCx11_ASAP7_75t_R g4065 ( 
.A(n_3826),
.Y(n_4065)
);

OAI21x1_ASAP7_75t_L g4066 ( 
.A1(n_3705),
.A2(n_3136),
.B(n_2863),
.Y(n_4066)
);

OAI21xp5_ASAP7_75t_L g4067 ( 
.A1(n_3857),
.A2(n_3140),
.B(n_3126),
.Y(n_4067)
);

AOI21xp5_ASAP7_75t_L g4068 ( 
.A1(n_3863),
.A2(n_3140),
.B(n_2317),
.Y(n_4068)
);

BUFx6f_ASAP7_75t_L g4069 ( 
.A(n_3481),
.Y(n_4069)
);

AOI21xp5_ASAP7_75t_L g4070 ( 
.A1(n_3706),
.A2(n_2317),
.B(n_2290),
.Y(n_4070)
);

BUFx6f_ASAP7_75t_L g4071 ( 
.A(n_3481),
.Y(n_4071)
);

NOR2xp33_ASAP7_75t_L g4072 ( 
.A(n_3757),
.B(n_3395),
.Y(n_4072)
);

AOI21xp33_ASAP7_75t_L g4073 ( 
.A1(n_3535),
.A2(n_3593),
.B(n_3807),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_SL g4074 ( 
.A(n_3738),
.B(n_3519),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3465),
.Y(n_4075)
);

AOI31xp67_ASAP7_75t_L g4076 ( 
.A1(n_3711),
.A2(n_2896),
.A3(n_2902),
.B(n_2881),
.Y(n_4076)
);

AOI21xp5_ASAP7_75t_L g4077 ( 
.A1(n_3808),
.A2(n_2317),
.B(n_2290),
.Y(n_4077)
);

OAI21xp5_ASAP7_75t_L g4078 ( 
.A1(n_3593),
.A2(n_3093),
.B(n_3086),
.Y(n_4078)
);

O2A1O1Ixp33_ASAP7_75t_SL g4079 ( 
.A1(n_3866),
.A2(n_3012),
.B(n_3082),
.C(n_3053),
.Y(n_4079)
);

O2A1O1Ixp33_ASAP7_75t_SL g4080 ( 
.A1(n_3475),
.A2(n_3012),
.B(n_3095),
.C(n_3082),
.Y(n_4080)
);

AOI221xp5_ASAP7_75t_L g4081 ( 
.A1(n_3649),
.A2(n_3093),
.B1(n_3112),
.B2(n_3113),
.C(n_3198),
.Y(n_4081)
);

A2O1A1Ixp33_ASAP7_75t_L g4082 ( 
.A1(n_3495),
.A2(n_3360),
.B(n_3380),
.C(n_3035),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_SL g4083 ( 
.A(n_3738),
.B(n_3377),
.Y(n_4083)
);

A2O1A1Ixp33_ASAP7_75t_L g4084 ( 
.A1(n_3875),
.A2(n_3380),
.B(n_3035),
.C(n_3089),
.Y(n_4084)
);

NAND3xp33_ASAP7_75t_L g4085 ( 
.A(n_3519),
.B(n_3120),
.C(n_3095),
.Y(n_4085)
);

NOR2xp33_ASAP7_75t_L g4086 ( 
.A(n_3657),
.B(n_3395),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_SL g4087 ( 
.A(n_3603),
.B(n_3381),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3465),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_3507),
.Y(n_4089)
);

AOI22xp5_ASAP7_75t_L g4090 ( 
.A1(n_3612),
.A2(n_2968),
.B1(n_3197),
.B2(n_2190),
.Y(n_4090)
);

CKINVDCx20_ASAP7_75t_R g4091 ( 
.A(n_3836),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3906),
.B(n_2873),
.Y(n_4092)
);

BUFx3_ASAP7_75t_L g4093 ( 
.A(n_3483),
.Y(n_4093)
);

OAI22xp33_ASAP7_75t_L g4094 ( 
.A1(n_3553),
.A2(n_3197),
.B1(n_2968),
.B2(n_3397),
.Y(n_4094)
);

OAI21xp5_ASAP7_75t_L g4095 ( 
.A1(n_3490),
.A2(n_3113),
.B(n_3112),
.Y(n_4095)
);

OAI21xp5_ASAP7_75t_L g4096 ( 
.A1(n_3490),
.A2(n_3022),
.B(n_3008),
.Y(n_4096)
);

OAI22x1_ASAP7_75t_L g4097 ( 
.A1(n_3608),
.A2(n_3380),
.B1(n_3069),
.B2(n_3094),
.Y(n_4097)
);

AO31x2_ASAP7_75t_L g4098 ( 
.A1(n_3733),
.A2(n_3329),
.A3(n_3368),
.B(n_3317),
.Y(n_4098)
);

INVx2_ASAP7_75t_L g4099 ( 
.A(n_3574),
.Y(n_4099)
);

O2A1O1Ixp33_ASAP7_75t_L g4100 ( 
.A1(n_3925),
.A2(n_3211),
.B(n_3235),
.C(n_3207),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3496),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3496),
.Y(n_4102)
);

BUFx3_ASAP7_75t_L g4103 ( 
.A(n_3990),
.Y(n_4103)
);

NOR2xp33_ASAP7_75t_L g4104 ( 
.A(n_3708),
.B(n_3166),
.Y(n_4104)
);

BUFx2_ASAP7_75t_L g4105 ( 
.A(n_3827),
.Y(n_4105)
);

OR2x2_ASAP7_75t_L g4106 ( 
.A(n_3545),
.B(n_3381),
.Y(n_4106)
);

HB1xp67_ASAP7_75t_L g4107 ( 
.A(n_3986),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_3906),
.B(n_2873),
.Y(n_4108)
);

NOR2xp33_ASAP7_75t_L g4109 ( 
.A(n_3708),
.B(n_3850),
.Y(n_4109)
);

O2A1O1Ixp33_ASAP7_75t_L g4110 ( 
.A1(n_3808),
.A2(n_3211),
.B(n_3235),
.C(n_3207),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_3907),
.B(n_2941),
.Y(n_4111)
);

OAI21x1_ASAP7_75t_SL g4112 ( 
.A1(n_3475),
.A2(n_3137),
.B(n_3120),
.Y(n_4112)
);

BUFx6f_ASAP7_75t_L g4113 ( 
.A(n_3481),
.Y(n_4113)
);

O2A1O1Ixp33_ASAP7_75t_SL g4114 ( 
.A1(n_3479),
.A2(n_3156),
.B(n_3157),
.C(n_3137),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3907),
.B(n_2941),
.Y(n_4115)
);

BUFx6f_ASAP7_75t_L g4116 ( 
.A(n_3481),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3501),
.Y(n_4117)
);

CKINVDCx6p67_ASAP7_75t_R g4118 ( 
.A(n_3990),
.Y(n_4118)
);

AND2x4_ASAP7_75t_L g4119 ( 
.A(n_3856),
.B(n_3397),
.Y(n_4119)
);

AO31x2_ASAP7_75t_L g4120 ( 
.A1(n_3733),
.A2(n_3329),
.A3(n_3368),
.B(n_3317),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3501),
.Y(n_4121)
);

O2A1O1Ixp33_ASAP7_75t_L g4122 ( 
.A1(n_3479),
.A2(n_3247),
.B(n_3157),
.C(n_3169),
.Y(n_4122)
);

AOI22xp5_ASAP7_75t_L g4123 ( 
.A1(n_3612),
.A2(n_2968),
.B1(n_3197),
.B2(n_2190),
.Y(n_4123)
);

INVx2_ASAP7_75t_L g4124 ( 
.A(n_3574),
.Y(n_4124)
);

AO31x2_ASAP7_75t_L g4125 ( 
.A1(n_3539),
.A2(n_3368),
.A3(n_3372),
.B(n_3329),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_3574),
.Y(n_4126)
);

BUFx2_ASAP7_75t_SL g4127 ( 
.A(n_3902),
.Y(n_4127)
);

AND2x4_ASAP7_75t_L g4128 ( 
.A(n_3856),
.B(n_3397),
.Y(n_4128)
);

AOI21xp5_ASAP7_75t_L g4129 ( 
.A1(n_3780),
.A2(n_2317),
.B(n_2290),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_3627),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3516),
.Y(n_4131)
);

OA21x2_ASAP7_75t_L g4132 ( 
.A1(n_3876),
.A2(n_3315),
.B(n_2896),
.Y(n_4132)
);

INVxp67_ASAP7_75t_L g4133 ( 
.A(n_3443),
.Y(n_4133)
);

AOI21xp5_ASAP7_75t_L g4134 ( 
.A1(n_3780),
.A2(n_2321),
.B(n_2317),
.Y(n_4134)
);

OAI21xp33_ASAP7_75t_L g4135 ( 
.A1(n_3590),
.A2(n_3169),
.B(n_3156),
.Y(n_4135)
);

AO31x2_ASAP7_75t_L g4136 ( 
.A1(n_3539),
.A2(n_3403),
.A3(n_3372),
.B(n_2495),
.Y(n_4136)
);

A2O1A1Ixp33_ASAP7_75t_L g4137 ( 
.A1(n_3875),
.A2(n_3035),
.B(n_3089),
.C(n_3050),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3930),
.B(n_3958),
.Y(n_4138)
);

NOR2xp33_ASAP7_75t_L g4139 ( 
.A(n_3764),
.B(n_3011),
.Y(n_4139)
);

OAI22xp5_ASAP7_75t_L g4140 ( 
.A1(n_3608),
.A2(n_2878),
.B1(n_2915),
.B2(n_2859),
.Y(n_4140)
);

O2A1O1Ixp33_ASAP7_75t_SL g4141 ( 
.A1(n_3955),
.A2(n_3177),
.B(n_3185),
.C(n_3173),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_3627),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3930),
.B(n_3011),
.Y(n_4143)
);

NAND2xp33_ASAP7_75t_L g4144 ( 
.A(n_3854),
.B(n_3003),
.Y(n_4144)
);

INVx4_ASAP7_75t_L g4145 ( 
.A(n_3687),
.Y(n_4145)
);

O2A1O1Ixp33_ASAP7_75t_SL g4146 ( 
.A1(n_3590),
.A2(n_3672),
.B(n_3530),
.C(n_3508),
.Y(n_4146)
);

AO31x2_ASAP7_75t_L g4147 ( 
.A1(n_3617),
.A2(n_3403),
.A3(n_3372),
.B(n_2495),
.Y(n_4147)
);

AO31x2_ASAP7_75t_L g4148 ( 
.A1(n_3617),
.A2(n_3403),
.A3(n_2507),
.B(n_2511),
.Y(n_4148)
);

INVxp67_ASAP7_75t_L g4149 ( 
.A(n_3677),
.Y(n_4149)
);

OAI221xp5_ASAP7_75t_L g4150 ( 
.A1(n_3621),
.A2(n_3188),
.B1(n_3184),
.B2(n_3198),
.C(n_3247),
.Y(n_4150)
);

AOI22xp33_ASAP7_75t_L g4151 ( 
.A1(n_3485),
.A2(n_2504),
.B1(n_3397),
.B2(n_2472),
.Y(n_4151)
);

O2A1O1Ixp33_ASAP7_75t_L g4152 ( 
.A1(n_3621),
.A2(n_3177),
.B(n_3185),
.C(n_3173),
.Y(n_4152)
);

A2O1A1Ixp33_ASAP7_75t_L g4153 ( 
.A1(n_3656),
.A2(n_3445),
.B(n_3868),
.C(n_3817),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3516),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_3958),
.B(n_3029),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_3457),
.B(n_3029),
.Y(n_4156)
);

INVx3_ASAP7_75t_L g4157 ( 
.A(n_3625),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_3627),
.Y(n_4158)
);

AOI21xp5_ASAP7_75t_L g4159 ( 
.A1(n_3521),
.A2(n_2340),
.B(n_2321),
.Y(n_4159)
);

NOR2xp33_ASAP7_75t_L g4160 ( 
.A(n_3732),
.B(n_3145),
.Y(n_4160)
);

OR2x2_ASAP7_75t_L g4161 ( 
.A(n_3545),
.B(n_3393),
.Y(n_4161)
);

OAI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_3560),
.A2(n_3022),
.B(n_3008),
.Y(n_4162)
);

OAI21xp5_ASAP7_75t_L g4163 ( 
.A1(n_3560),
.A2(n_3043),
.B(n_3025),
.Y(n_4163)
);

OAI22xp33_ASAP7_75t_L g4164 ( 
.A1(n_3553),
.A2(n_3197),
.B1(n_2968),
.B2(n_3397),
.Y(n_4164)
);

AND2x4_ASAP7_75t_L g4165 ( 
.A(n_3856),
.B(n_3897),
.Y(n_4165)
);

INVx2_ASAP7_75t_SL g4166 ( 
.A(n_3754),
.Y(n_4166)
);

BUFx6f_ASAP7_75t_L g4167 ( 
.A(n_3482),
.Y(n_4167)
);

AOI211x1_ASAP7_75t_L g4168 ( 
.A1(n_3597),
.A2(n_3145),
.B(n_3159),
.C(n_3167),
.Y(n_4168)
);

NAND2x1_ASAP7_75t_L g4169 ( 
.A(n_3935),
.B(n_3212),
.Y(n_4169)
);

HB1xp67_ASAP7_75t_L g4170 ( 
.A(n_3798),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3526),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3526),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_3529),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_L g4174 ( 
.A1(n_3485),
.A2(n_2504),
.B1(n_2472),
.B2(n_2190),
.Y(n_4174)
);

NOR2xp33_ASAP7_75t_L g4175 ( 
.A(n_3640),
.B(n_3167),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_3529),
.Y(n_4176)
);

O2A1O1Ixp33_ASAP7_75t_L g4177 ( 
.A1(n_3649),
.A2(n_3535),
.B(n_3534),
.C(n_3616),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_3457),
.B(n_3226),
.Y(n_4178)
);

BUFx6f_ASAP7_75t_L g4179 ( 
.A(n_3482),
.Y(n_4179)
);

BUFx3_ASAP7_75t_L g4180 ( 
.A(n_3591),
.Y(n_4180)
);

NAND2x1_ASAP7_75t_L g4181 ( 
.A(n_3935),
.B(n_3810),
.Y(n_4181)
);

AOI221x1_ASAP7_75t_L g4182 ( 
.A1(n_3800),
.A2(n_3208),
.B1(n_3238),
.B2(n_3193),
.C(n_3191),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3536),
.Y(n_4183)
);

OAI22xp5_ASAP7_75t_SL g4184 ( 
.A1(n_3794),
.A2(n_3292),
.B1(n_3138),
.B2(n_2878),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3637),
.Y(n_4185)
);

AND2x4_ASAP7_75t_L g4186 ( 
.A(n_3856),
.B(n_3292),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3536),
.Y(n_4187)
);

AO32x2_ASAP7_75t_L g4188 ( 
.A1(n_3461),
.A2(n_2915),
.A3(n_3064),
.B1(n_2878),
.B2(n_2859),
.Y(n_4188)
);

A2O1A1Ixp33_ASAP7_75t_L g4189 ( 
.A1(n_3656),
.A2(n_3050),
.B(n_3178),
.C(n_3089),
.Y(n_4189)
);

A2O1A1Ixp33_ASAP7_75t_L g4190 ( 
.A1(n_3868),
.A2(n_3050),
.B(n_3190),
.C(n_3178),
.Y(n_4190)
);

O2A1O1Ixp33_ASAP7_75t_SL g4191 ( 
.A1(n_3672),
.A2(n_3193),
.B(n_3208),
.C(n_3191),
.Y(n_4191)
);

AOI21xp5_ASAP7_75t_L g4192 ( 
.A1(n_3531),
.A2(n_2340),
.B(n_2321),
.Y(n_4192)
);

A2O1A1Ixp33_ASAP7_75t_L g4193 ( 
.A1(n_3817),
.A2(n_3190),
.B(n_3259),
.C(n_3178),
.Y(n_4193)
);

NOR2xp33_ASAP7_75t_SL g4194 ( 
.A(n_3964),
.B(n_2915),
.Y(n_4194)
);

A2O1A1Ixp33_ASAP7_75t_L g4195 ( 
.A1(n_3534),
.A2(n_3259),
.B(n_3272),
.C(n_3190),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_3637),
.Y(n_4196)
);

OAI21xp5_ASAP7_75t_L g4197 ( 
.A1(n_3625),
.A2(n_3043),
.B(n_3025),
.Y(n_4197)
);

AOI22xp33_ASAP7_75t_L g4198 ( 
.A1(n_3485),
.A2(n_3638),
.B1(n_3580),
.B2(n_3684),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_3537),
.Y(n_4199)
);

OAI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_3794),
.A2(n_3064),
.B1(n_2886),
.B2(n_3159),
.Y(n_4200)
);

AOI221x1_ASAP7_75t_L g4201 ( 
.A1(n_3800),
.A2(n_3643),
.B1(n_3454),
.B2(n_3941),
.C(n_3668),
.Y(n_4201)
);

INVxp67_ASAP7_75t_SL g4202 ( 
.A(n_3595),
.Y(n_4202)
);

OR2x2_ASAP7_75t_L g4203 ( 
.A(n_3554),
.B(n_3393),
.Y(n_4203)
);

AOI21xp5_ASAP7_75t_L g4204 ( 
.A1(n_3567),
.A2(n_2340),
.B(n_2321),
.Y(n_4204)
);

INVx5_ASAP7_75t_L g4205 ( 
.A(n_3682),
.Y(n_4205)
);

AND2x2_ASAP7_75t_L g4206 ( 
.A(n_3689),
.B(n_3226),
.Y(n_4206)
);

OAI22xp5_ASAP7_75t_L g4207 ( 
.A1(n_3647),
.A2(n_3064),
.B1(n_2886),
.B2(n_2732),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_3462),
.B(n_3212),
.Y(n_4208)
);

INVx5_ASAP7_75t_L g4209 ( 
.A(n_3682),
.Y(n_4209)
);

O2A1O1Ixp33_ASAP7_75t_L g4210 ( 
.A1(n_3616),
.A2(n_3249),
.B(n_3252),
.C(n_3238),
.Y(n_4210)
);

OA21x2_ASAP7_75t_L g4211 ( 
.A1(n_3876),
.A2(n_2902),
.B(n_2881),
.Y(n_4211)
);

INVxp67_ASAP7_75t_SL g4212 ( 
.A(n_3595),
.Y(n_4212)
);

CKINVDCx20_ASAP7_75t_R g4213 ( 
.A(n_3591),
.Y(n_4213)
);

INVx3_ASAP7_75t_L g4214 ( 
.A(n_3989),
.Y(n_4214)
);

INVx2_ASAP7_75t_SL g4215 ( 
.A(n_3775),
.Y(n_4215)
);

OAI22xp33_ASAP7_75t_L g4216 ( 
.A1(n_3623),
.A2(n_2504),
.B1(n_3292),
.B2(n_3272),
.Y(n_4216)
);

AO21x1_ASAP7_75t_L g4217 ( 
.A1(n_3533),
.A2(n_3252),
.B(n_3249),
.Y(n_4217)
);

AOI21xp5_ASAP7_75t_L g4218 ( 
.A1(n_3567),
.A2(n_2359),
.B(n_2340),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_3537),
.Y(n_4219)
);

AOI21xp5_ASAP7_75t_L g4220 ( 
.A1(n_3565),
.A2(n_2411),
.B(n_2359),
.Y(n_4220)
);

A2O1A1Ixp33_ASAP7_75t_L g4221 ( 
.A1(n_3912),
.A2(n_3272),
.B(n_3299),
.C(n_3259),
.Y(n_4221)
);

A2O1A1Ixp33_ASAP7_75t_L g4222 ( 
.A1(n_3912),
.A2(n_3310),
.B(n_3321),
.C(n_3299),
.Y(n_4222)
);

NOR2xp33_ASAP7_75t_L g4223 ( 
.A(n_3523),
.B(n_3394),
.Y(n_4223)
);

O2A1O1Ixp33_ASAP7_75t_SL g4224 ( 
.A1(n_3508),
.A2(n_3297),
.B(n_3303),
.C(n_3286),
.Y(n_4224)
);

INVxp67_ASAP7_75t_SL g4225 ( 
.A(n_3604),
.Y(n_4225)
);

OAI21x1_ASAP7_75t_L g4226 ( 
.A1(n_3447),
.A2(n_3471),
.B(n_3701),
.Y(n_4226)
);

OAI22xp5_ASAP7_75t_L g4227 ( 
.A1(n_3647),
.A2(n_3064),
.B1(n_2732),
.B2(n_2689),
.Y(n_4227)
);

OAI22xp5_ASAP7_75t_L g4228 ( 
.A1(n_3647),
.A2(n_2732),
.B1(n_2689),
.B2(n_3138),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3544),
.Y(n_4229)
);

BUFx2_ASAP7_75t_L g4230 ( 
.A(n_3827),
.Y(n_4230)
);

BUFx2_ASAP7_75t_L g4231 ( 
.A(n_3832),
.Y(n_4231)
);

NOR2xp33_ASAP7_75t_L g4232 ( 
.A(n_3601),
.B(n_3394),
.Y(n_4232)
);

AOI21xp5_ASAP7_75t_L g4233 ( 
.A1(n_3565),
.A2(n_2411),
.B(n_2359),
.Y(n_4233)
);

O2A1O1Ixp33_ASAP7_75t_L g4234 ( 
.A1(n_3604),
.A2(n_3297),
.B(n_3303),
.C(n_3286),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_3637),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_3544),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_3550),
.Y(n_4237)
);

NAND2x1p5_ASAP7_75t_L g4238 ( 
.A(n_3883),
.B(n_2275),
.Y(n_4238)
);

AOI22xp33_ASAP7_75t_L g4239 ( 
.A1(n_3638),
.A2(n_2472),
.B1(n_2500),
.B2(n_2498),
.Y(n_4239)
);

HB1xp67_ASAP7_75t_L g4240 ( 
.A(n_3799),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_3642),
.Y(n_4241)
);

INVx2_ASAP7_75t_SL g4242 ( 
.A(n_3775),
.Y(n_4242)
);

AOI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_3927),
.A2(n_2411),
.B(n_2359),
.Y(n_4243)
);

A2O1A1Ixp33_ASAP7_75t_L g4244 ( 
.A1(n_3618),
.A2(n_3352),
.B(n_3407),
.C(n_3322),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_3462),
.B(n_3219),
.Y(n_4245)
);

AOI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_3927),
.A2(n_2411),
.B(n_2359),
.Y(n_4246)
);

AOI21xp5_ASAP7_75t_L g4247 ( 
.A1(n_3610),
.A2(n_2411),
.B(n_2359),
.Y(n_4247)
);

O2A1O1Ixp33_ASAP7_75t_L g4248 ( 
.A1(n_3613),
.A2(n_3370),
.B(n_3385),
.C(n_3304),
.Y(n_4248)
);

AOI22xp33_ASAP7_75t_L g4249 ( 
.A1(n_3638),
.A2(n_2472),
.B1(n_2500),
.B2(n_2498),
.Y(n_4249)
);

OA21x2_ASAP7_75t_L g4250 ( 
.A1(n_3890),
.A2(n_2902),
.B(n_2881),
.Y(n_4250)
);

AOI21xp5_ASAP7_75t_L g4251 ( 
.A1(n_3610),
.A2(n_3611),
.B(n_3605),
.Y(n_4251)
);

AO21x1_ASAP7_75t_L g4252 ( 
.A1(n_3533),
.A2(n_3370),
.B(n_3304),
.Y(n_4252)
);

BUFx2_ASAP7_75t_L g4253 ( 
.A(n_3832),
.Y(n_4253)
);

NOR2xp33_ASAP7_75t_L g4254 ( 
.A(n_3809),
.B(n_3219),
.Y(n_4254)
);

OAI22x1_ASAP7_75t_L g4255 ( 
.A1(n_3623),
.A2(n_3069),
.B1(n_3094),
.B2(n_3033),
.Y(n_4255)
);

OAI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_3755),
.A2(n_3386),
.B(n_3385),
.Y(n_4256)
);

A2O1A1Ixp33_ASAP7_75t_L g4257 ( 
.A1(n_3602),
.A2(n_3352),
.B(n_3407),
.C(n_3322),
.Y(n_4257)
);

BUFx2_ASAP7_75t_L g4258 ( 
.A(n_3842),
.Y(n_4258)
);

NOR2xp33_ASAP7_75t_L g4259 ( 
.A(n_3557),
.B(n_3261),
.Y(n_4259)
);

OAI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_3755),
.A2(n_3400),
.B(n_3386),
.Y(n_4260)
);

NAND2x1_ASAP7_75t_L g4261 ( 
.A(n_3810),
.B(n_3261),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_3550),
.Y(n_4262)
);

OR2x2_ASAP7_75t_L g4263 ( 
.A(n_3554),
.B(n_3285),
.Y(n_4263)
);

AOI222xp33_ASAP7_75t_L g4264 ( 
.A1(n_3684),
.A2(n_3184),
.B1(n_3188),
.B2(n_3279),
.C1(n_3290),
.C2(n_3274),
.Y(n_4264)
);

INVx1_ASAP7_75t_SL g4265 ( 
.A(n_3557),
.Y(n_4265)
);

AOI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_3664),
.A2(n_2419),
.B(n_2417),
.Y(n_4266)
);

O2A1O1Ixp33_ASAP7_75t_SL g4267 ( 
.A1(n_3530),
.A2(n_3438),
.B(n_3400),
.C(n_3241),
.Y(n_4267)
);

AOI21xp5_ASAP7_75t_L g4268 ( 
.A1(n_3664),
.A2(n_2419),
.B(n_2417),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_3586),
.B(n_3589),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_3586),
.B(n_3285),
.Y(n_4270)
);

AOI22xp5_ASAP7_75t_L g4271 ( 
.A1(n_3744),
.A2(n_3069),
.B1(n_3094),
.B2(n_3033),
.Y(n_4271)
);

NOR2xp33_ASAP7_75t_L g4272 ( 
.A(n_3589),
.B(n_3231),
.Y(n_4272)
);

NOR2xp33_ASAP7_75t_L g4273 ( 
.A(n_3592),
.B(n_3231),
.Y(n_4273)
);

OAI21xp5_ASAP7_75t_L g4274 ( 
.A1(n_3613),
.A2(n_3438),
.B(n_3269),
.Y(n_4274)
);

AOI221x1_ASAP7_75t_L g4275 ( 
.A1(n_3643),
.A2(n_3290),
.B1(n_3255),
.B2(n_3269),
.C(n_3271),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3573),
.Y(n_4276)
);

AO32x2_ASAP7_75t_L g4277 ( 
.A1(n_3461),
.A2(n_2329),
.A3(n_2357),
.B1(n_2312),
.B2(n_2489),
.Y(n_4277)
);

INVxp67_ASAP7_75t_SL g4278 ( 
.A(n_3615),
.Y(n_4278)
);

INVxp67_ASAP7_75t_SL g4279 ( 
.A(n_3615),
.Y(n_4279)
);

AOI21x1_ASAP7_75t_L g4280 ( 
.A1(n_3719),
.A2(n_2923),
.B(n_2911),
.Y(n_4280)
);

NOR2xp33_ASAP7_75t_L g4281 ( 
.A(n_3592),
.B(n_3231),
.Y(n_4281)
);

INVx3_ASAP7_75t_L g4282 ( 
.A(n_3989),
.Y(n_4282)
);

NAND2xp5_ASAP7_75t_L g4283 ( 
.A(n_3641),
.B(n_3255),
.Y(n_4283)
);

OAI22xp5_ASAP7_75t_L g4284 ( 
.A1(n_3603),
.A2(n_2732),
.B1(n_2689),
.B2(n_3352),
.Y(n_4284)
);

A2O1A1Ixp33_ASAP7_75t_L g4285 ( 
.A1(n_3833),
.A2(n_3407),
.B(n_3094),
.C(n_3128),
.Y(n_4285)
);

BUFx3_ASAP7_75t_L g4286 ( 
.A(n_3591),
.Y(n_4286)
);

BUFx2_ASAP7_75t_L g4287 ( 
.A(n_3842),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_3641),
.B(n_3271),
.Y(n_4288)
);

INVx2_ASAP7_75t_L g4289 ( 
.A(n_3642),
.Y(n_4289)
);

INVx1_ASAP7_75t_SL g4290 ( 
.A(n_3714),
.Y(n_4290)
);

OAI21x1_ASAP7_75t_L g4291 ( 
.A1(n_3776),
.A2(n_3335),
.B(n_3334),
.Y(n_4291)
);

AOI21xp5_ASAP7_75t_L g4292 ( 
.A1(n_3585),
.A2(n_3828),
.B(n_3806),
.Y(n_4292)
);

BUFx6f_ASAP7_75t_L g4293 ( 
.A(n_3482),
.Y(n_4293)
);

OAI21xp5_ASAP7_75t_L g4294 ( 
.A1(n_3620),
.A2(n_3287),
.B(n_3274),
.Y(n_4294)
);

AOI22xp5_ASAP7_75t_L g4295 ( 
.A1(n_3744),
.A2(n_3128),
.B1(n_3129),
.B2(n_3069),
.Y(n_4295)
);

AO31x2_ASAP7_75t_L g4296 ( 
.A1(n_3548),
.A2(n_2507),
.A3(n_2511),
.B(n_2486),
.Y(n_4296)
);

AND2x4_ASAP7_75t_L g4297 ( 
.A(n_3897),
.B(n_3128),
.Y(n_4297)
);

AOI21xp5_ASAP7_75t_L g4298 ( 
.A1(n_3585),
.A2(n_2419),
.B(n_3287),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_3573),
.Y(n_4299)
);

O2A1O1Ixp33_ASAP7_75t_SL g4300 ( 
.A1(n_3464),
.A2(n_3439),
.B(n_3335),
.C(n_3339),
.Y(n_4300)
);

INVx5_ASAP7_75t_L g4301 ( 
.A(n_3682),
.Y(n_4301)
);

AND2x2_ASAP7_75t_L g4302 ( 
.A(n_3459),
.B(n_3335),
.Y(n_4302)
);

A2O1A1Ixp33_ASAP7_75t_L g4303 ( 
.A1(n_3833),
.A2(n_3128),
.B(n_3129),
.C(n_3135),
.Y(n_4303)
);

AO32x2_ASAP7_75t_L g4304 ( 
.A1(n_3478),
.A2(n_2489),
.A3(n_2357),
.B1(n_2329),
.B2(n_2312),
.Y(n_4304)
);

A2O1A1Ixp33_ASAP7_75t_L g4305 ( 
.A1(n_3582),
.A2(n_3135),
.B(n_3129),
.C(n_3141),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_3642),
.Y(n_4306)
);

NAND2x1p5_ASAP7_75t_L g4307 ( 
.A(n_3883),
.B(n_2275),
.Y(n_4307)
);

BUFx10_ASAP7_75t_L g4308 ( 
.A(n_3482),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_3459),
.B(n_3339),
.Y(n_4309)
);

NOR2xp33_ASAP7_75t_L g4310 ( 
.A(n_3714),
.B(n_3231),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_3512),
.B(n_3339),
.Y(n_4311)
);

AOI21xp33_ASAP7_75t_L g4312 ( 
.A1(n_3789),
.A2(n_3306),
.B(n_3296),
.Y(n_4312)
);

AO32x2_ASAP7_75t_L g4313 ( 
.A1(n_3478),
.A2(n_2357),
.A3(n_2329),
.B1(n_2312),
.B2(n_2489),
.Y(n_4313)
);

OAI21xp5_ASAP7_75t_L g4314 ( 
.A1(n_3620),
.A2(n_3306),
.B(n_3296),
.Y(n_4314)
);

INVx3_ASAP7_75t_L g4315 ( 
.A(n_3715),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_3583),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_3645),
.Y(n_4317)
);

HB1xp67_ASAP7_75t_L g4318 ( 
.A(n_3851),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_3788),
.B(n_3740),
.Y(n_4319)
);

OR2x2_ASAP7_75t_L g4320 ( 
.A(n_3777),
.B(n_3683),
.Y(n_4320)
);

O2A1O1Ixp33_ASAP7_75t_SL g4321 ( 
.A1(n_3464),
.A2(n_3439),
.B(n_3278),
.C(n_3426),
.Y(n_4321)
);

AOI21xp5_ASAP7_75t_L g4322 ( 
.A1(n_3828),
.A2(n_3548),
.B(n_3786),
.Y(n_4322)
);

AND2x6_ASAP7_75t_L g4323 ( 
.A(n_3473),
.B(n_2275),
.Y(n_4323)
);

AO31x2_ASAP7_75t_L g4324 ( 
.A1(n_3840),
.A2(n_2507),
.A3(n_2511),
.B(n_2524),
.Y(n_4324)
);

OAI21x1_ASAP7_75t_L g4325 ( 
.A1(n_3783),
.A2(n_3439),
.B(n_3189),
.Y(n_4325)
);

CKINVDCx6p67_ASAP7_75t_R g4326 ( 
.A(n_3687),
.Y(n_4326)
);

AOI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_3802),
.A2(n_3311),
.B(n_2702),
.Y(n_4327)
);

AO31x2_ASAP7_75t_L g4328 ( 
.A1(n_3840),
.A2(n_2507),
.A3(n_2511),
.B(n_2524),
.Y(n_4328)
);

BUFx2_ASAP7_75t_L g4329 ( 
.A(n_3847),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_3583),
.Y(n_4330)
);

NAND2x2_ASAP7_75t_L g4331 ( 
.A(n_3484),
.B(n_3278),
.Y(n_4331)
);

AOI22xp5_ASAP7_75t_L g4332 ( 
.A1(n_3561),
.A2(n_3135),
.B1(n_3141),
.B2(n_2959),
.Y(n_4332)
);

A2O1A1Ixp33_ASAP7_75t_L g4333 ( 
.A1(n_3598),
.A2(n_3141),
.B(n_2927),
.C(n_2999),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_3588),
.Y(n_4334)
);

AO21x1_ASAP7_75t_L g4335 ( 
.A1(n_3559),
.A2(n_3311),
.B(n_2959),
.Y(n_4335)
);

OR2x2_ASAP7_75t_L g4336 ( 
.A(n_3777),
.B(n_2911),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_3788),
.B(n_3439),
.Y(n_4337)
);

O2A1O1Ixp33_ASAP7_75t_L g4338 ( 
.A1(n_3622),
.A2(n_3045),
.B(n_2923),
.C(n_2924),
.Y(n_4338)
);

AOI22xp33_ASAP7_75t_L g4339 ( 
.A1(n_3580),
.A2(n_2472),
.B1(n_2498),
.B2(n_2500),
.Y(n_4339)
);

AOI22xp33_ASAP7_75t_L g4340 ( 
.A1(n_3580),
.A2(n_2472),
.B1(n_2498),
.B2(n_2500),
.Y(n_4340)
);

CKINVDCx5p33_ASAP7_75t_R g4341 ( 
.A(n_3609),
.Y(n_4341)
);

AOI21xp5_ASAP7_75t_L g4342 ( 
.A1(n_3945),
.A2(n_2702),
.B(n_2653),
.Y(n_4342)
);

O2A1O1Ixp33_ASAP7_75t_L g4343 ( 
.A1(n_3622),
.A2(n_3099),
.B(n_2987),
.C(n_2924),
.Y(n_4343)
);

OAI22xp5_ASAP7_75t_L g4344 ( 
.A1(n_3551),
.A2(n_2927),
.B1(n_2959),
.B2(n_2999),
.Y(n_4344)
);

NOR2xp33_ASAP7_75t_L g4345 ( 
.A(n_3740),
.B(n_3607),
.Y(n_4345)
);

O2A1O1Ixp33_ASAP7_75t_SL g4346 ( 
.A1(n_3469),
.A2(n_3426),
.B(n_3278),
.C(n_3233),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_L g4347 ( 
.A(n_3716),
.B(n_3787),
.Y(n_4347)
);

OAI22xp33_ASAP7_75t_L g4348 ( 
.A1(n_3561),
.A2(n_2472),
.B1(n_2498),
.B2(n_2500),
.Y(n_4348)
);

OAI22xp33_ASAP7_75t_L g4349 ( 
.A1(n_3835),
.A2(n_2500),
.B1(n_2498),
.B2(n_2580),
.Y(n_4349)
);

AOI22xp5_ASAP7_75t_L g4350 ( 
.A1(n_3789),
.A2(n_2959),
.B1(n_2927),
.B2(n_3013),
.Y(n_4350)
);

O2A1O1Ixp33_ASAP7_75t_L g4351 ( 
.A1(n_3635),
.A2(n_3100),
.B(n_2987),
.C(n_3015),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_3588),
.Y(n_4352)
);

AOI22xp33_ASAP7_75t_L g4353 ( 
.A1(n_3454),
.A2(n_2500),
.B1(n_3280),
.B2(n_3309),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_3645),
.Y(n_4354)
);

AO31x2_ASAP7_75t_L g4355 ( 
.A1(n_3902),
.A2(n_2555),
.A3(n_2524),
.B(n_2541),
.Y(n_4355)
);

OR2x2_ASAP7_75t_L g4356 ( 
.A(n_3683),
.B(n_2957),
.Y(n_4356)
);

AO32x2_ASAP7_75t_L g4357 ( 
.A1(n_3915),
.A2(n_3924),
.A3(n_3954),
.B1(n_3919),
.B2(n_3933),
.Y(n_4357)
);

AOI22xp33_ASAP7_75t_L g4358 ( 
.A1(n_3758),
.A2(n_3309),
.B1(n_3280),
.B2(n_2927),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_3787),
.B(n_3049),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_3594),
.Y(n_4360)
);

NOR2xp33_ASAP7_75t_L g4361 ( 
.A(n_3607),
.B(n_3278),
.Y(n_4361)
);

O2A1O1Ixp33_ASAP7_75t_SL g4362 ( 
.A1(n_3469),
.A2(n_3426),
.B(n_3233),
.C(n_2809),
.Y(n_4362)
);

AND2x4_ASAP7_75t_L g4363 ( 
.A(n_3897),
.B(n_2999),
.Y(n_4363)
);

BUFx8_ASAP7_75t_L g4364 ( 
.A(n_3569),
.Y(n_4364)
);

BUFx5_ASAP7_75t_L g4365 ( 
.A(n_3815),
.Y(n_4365)
);

AOI221x1_ASAP7_75t_L g4366 ( 
.A1(n_3941),
.A2(n_2837),
.B1(n_2254),
.B2(n_2253),
.C(n_2264),
.Y(n_4366)
);

INVx3_ASAP7_75t_L g4367 ( 
.A(n_3715),
.Y(n_4367)
);

AND2x4_ASAP7_75t_L g4368 ( 
.A(n_3897),
.B(n_2999),
.Y(n_4368)
);

AOI21xp5_ASAP7_75t_L g4369 ( 
.A1(n_3821),
.A2(n_3823),
.B(n_3797),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_3718),
.B(n_3049),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_3594),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_3718),
.B(n_3049),
.Y(n_4372)
);

HB1xp67_ASAP7_75t_L g4373 ( 
.A(n_3847),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_3614),
.Y(n_4374)
);

AND2x4_ASAP7_75t_L g4375 ( 
.A(n_3929),
.B(n_3013),
.Y(n_4375)
);

O2A1O1Ixp33_ASAP7_75t_SL g4376 ( 
.A1(n_3908),
.A2(n_3497),
.B(n_3514),
.C(n_3849),
.Y(n_4376)
);

AOI221x1_ASAP7_75t_L g4377 ( 
.A1(n_3668),
.A2(n_2837),
.B1(n_2254),
.B2(n_2264),
.C(n_2265),
.Y(n_4377)
);

AND2x2_ASAP7_75t_L g4378 ( 
.A(n_3512),
.B(n_3049),
.Y(n_4378)
);

OAI21xp33_ASAP7_75t_L g4379 ( 
.A1(n_3723),
.A2(n_3728),
.B(n_3644),
.Y(n_4379)
);

NOR2xp33_ASAP7_75t_L g4380 ( 
.A(n_3679),
.B(n_3426),
.Y(n_4380)
);

AOI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_3797),
.A2(n_2702),
.B(n_2653),
.Y(n_4381)
);

AOI21xp5_ASAP7_75t_L g4382 ( 
.A1(n_3795),
.A2(n_2702),
.B(n_2528),
.Y(n_4382)
);

AOI22xp5_ASAP7_75t_L g4383 ( 
.A1(n_3558),
.A2(n_3013),
.B1(n_3309),
.B2(n_3280),
.Y(n_4383)
);

BUFx6f_ASAP7_75t_L g4384 ( 
.A(n_3482),
.Y(n_4384)
);

AND2x4_ASAP7_75t_L g4385 ( 
.A(n_3929),
.B(n_3013),
.Y(n_4385)
);

AOI22xp33_ASAP7_75t_L g4386 ( 
.A1(n_3835),
.A2(n_3280),
.B1(n_3309),
.B2(n_2840),
.Y(n_4386)
);

AOI21xp5_ASAP7_75t_L g4387 ( 
.A1(n_3792),
.A2(n_2528),
.B(n_2312),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_3614),
.Y(n_4388)
);

AO31x2_ASAP7_75t_L g4389 ( 
.A1(n_3559),
.A2(n_2524),
.A3(n_2539),
.B(n_2529),
.Y(n_4389)
);

OR2x2_ASAP7_75t_L g4390 ( 
.A(n_3694),
.B(n_2961),
.Y(n_4390)
);

AOI221xp5_ASAP7_75t_L g4391 ( 
.A1(n_3723),
.A2(n_2961),
.B1(n_3024),
.B2(n_3045),
.C(n_3015),
.Y(n_4391)
);

INVx2_ASAP7_75t_L g4392 ( 
.A(n_3645),
.Y(n_4392)
);

BUFx3_ASAP7_75t_L g4393 ( 
.A(n_3591),
.Y(n_4393)
);

A2O1A1Ixp33_ASAP7_75t_L g4394 ( 
.A1(n_3599),
.A2(n_2358),
.B(n_2412),
.C(n_3015),
.Y(n_4394)
);

OAI22xp33_ASAP7_75t_L g4395 ( 
.A1(n_3728),
.A2(n_2809),
.B1(n_2580),
.B2(n_2562),
.Y(n_4395)
);

INVx2_ASAP7_75t_L g4396 ( 
.A(n_3665),
.Y(n_4396)
);

CKINVDCx5p33_ASAP7_75t_R g4397 ( 
.A(n_3848),
.Y(n_4397)
);

OAI22xp5_ASAP7_75t_L g4398 ( 
.A1(n_3456),
.A2(n_3436),
.B1(n_3412),
.B2(n_3396),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_3449),
.B(n_3049),
.Y(n_4399)
);

BUFx2_ASAP7_75t_L g4400 ( 
.A(n_3480),
.Y(n_4400)
);

OAI21xp5_ASAP7_75t_L g4401 ( 
.A1(n_3635),
.A2(n_2528),
.B(n_2605),
.Y(n_4401)
);

OR2x6_ASAP7_75t_L g4402 ( 
.A(n_3881),
.B(n_2840),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_3633),
.B(n_3049),
.Y(n_4403)
);

INVx1_ASAP7_75t_SL g4404 ( 
.A(n_3872),
.Y(n_4404)
);

OA21x2_ASAP7_75t_L g4405 ( 
.A1(n_3898),
.A2(n_3024),
.B(n_2986),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_3449),
.B(n_3134),
.Y(n_4406)
);

AOI221xp5_ASAP7_75t_L g4407 ( 
.A1(n_3784),
.A2(n_3045),
.B1(n_3048),
.B2(n_3087),
.C(n_3092),
.Y(n_4407)
);

AOI21xp5_ASAP7_75t_L g4408 ( 
.A1(n_3792),
.A2(n_3882),
.B(n_3984),
.Y(n_4408)
);

INVx3_ASAP7_75t_L g4409 ( 
.A(n_3846),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_3633),
.B(n_3134),
.Y(n_4410)
);

AND2x2_ASAP7_75t_L g4411 ( 
.A(n_3634),
.B(n_3134),
.Y(n_4411)
);

AOI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_3882),
.A2(n_3472),
.B(n_3470),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_3624),
.Y(n_4413)
);

OAI22xp33_ASAP7_75t_L g4414 ( 
.A1(n_3812),
.A2(n_2809),
.B1(n_2561),
.B2(n_2563),
.Y(n_4414)
);

AOI22xp33_ASAP7_75t_SL g4415 ( 
.A1(n_3901),
.A2(n_3233),
.B1(n_2809),
.B2(n_2840),
.Y(n_4415)
);

AO32x2_ASAP7_75t_L g4416 ( 
.A1(n_3915),
.A2(n_2489),
.A3(n_2357),
.B1(n_2296),
.B2(n_3092),
.Y(n_4416)
);

O2A1O1Ixp33_ASAP7_75t_L g4417 ( 
.A1(n_3652),
.A2(n_3048),
.B(n_3087),
.C(n_3092),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_3624),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_3667),
.Y(n_4419)
);

AOI22xp5_ASAP7_75t_L g4420 ( 
.A1(n_3632),
.A2(n_2261),
.B1(n_2592),
.B2(n_2840),
.Y(n_4420)
);

NOR2x1_ASAP7_75t_L g4421 ( 
.A(n_3702),
.B(n_2425),
.Y(n_4421)
);

AOI22xp33_ASAP7_75t_SL g4422 ( 
.A1(n_3901),
.A2(n_3233),
.B1(n_2840),
.B2(n_2261),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_L g4423 ( 
.A(n_3753),
.B(n_3134),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_3667),
.Y(n_4424)
);

BUFx12f_ASAP7_75t_L g4425 ( 
.A(n_3484),
.Y(n_4425)
);

NOR2xp67_ASAP7_75t_SL g4426 ( 
.A(n_3801),
.B(n_2334),
.Y(n_4426)
);

O2A1O1Ixp33_ASAP7_75t_SL g4427 ( 
.A1(n_3497),
.A2(n_2412),
.B(n_2358),
.C(n_3214),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_L g4428 ( 
.A(n_3753),
.B(n_3134),
.Y(n_4428)
);

INVxp67_ASAP7_75t_SL g4429 ( 
.A(n_3660),
.Y(n_4429)
);

BUFx6f_ASAP7_75t_L g4430 ( 
.A(n_3482),
.Y(n_4430)
);

NOR2x1_ASAP7_75t_SL g4431 ( 
.A(n_3801),
.B(n_3134),
.Y(n_4431)
);

NOR2xp33_ASAP7_75t_L g4432 ( 
.A(n_3679),
.B(n_3155),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_3681),
.Y(n_4433)
);

AOI22xp5_ASAP7_75t_L g4434 ( 
.A1(n_3731),
.A2(n_2261),
.B1(n_2592),
.B2(n_2840),
.Y(n_4434)
);

HB1xp67_ASAP7_75t_L g4435 ( 
.A(n_3963),
.Y(n_4435)
);

NAND2x1p5_ASAP7_75t_L g4436 ( 
.A(n_3682),
.B(n_2334),
.Y(n_4436)
);

O2A1O1Ixp33_ASAP7_75t_L g4437 ( 
.A1(n_3660),
.A2(n_3172),
.B(n_3099),
.C(n_3100),
.Y(n_4437)
);

BUFx12f_ASAP7_75t_L g4438 ( 
.A(n_3484),
.Y(n_4438)
);

A2O1A1Ixp33_ASAP7_75t_L g4439 ( 
.A1(n_3812),
.A2(n_2358),
.B(n_2412),
.C(n_3099),
.Y(n_4439)
);

INVx3_ASAP7_75t_L g4440 ( 
.A(n_3846),
.Y(n_4440)
);

A2O1A1Ixp33_ASAP7_75t_L g4441 ( 
.A1(n_3546),
.A2(n_2358),
.B(n_2412),
.C(n_3220),
.Y(n_4441)
);

OAI21xp5_ASAP7_75t_L g4442 ( 
.A1(n_3670),
.A2(n_3549),
.B(n_3522),
.Y(n_4442)
);

OA21x2_ASAP7_75t_L g4443 ( 
.A1(n_3913),
.A2(n_3123),
.B(n_3139),
.Y(n_4443)
);

AO32x2_ASAP7_75t_L g4444 ( 
.A1(n_3919),
.A2(n_3123),
.A3(n_3139),
.B1(n_3172),
.B2(n_3176),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_L g4445 ( 
.A(n_3763),
.B(n_3155),
.Y(n_4445)
);

CKINVDCx9p33_ASAP7_75t_R g4446 ( 
.A(n_3480),
.Y(n_4446)
);

OR2x2_ASAP7_75t_L g4447 ( 
.A(n_3694),
.B(n_3176),
.Y(n_4447)
);

BUFx2_ASAP7_75t_L g4448 ( 
.A(n_3510),
.Y(n_4448)
);

INVxp67_ASAP7_75t_L g4449 ( 
.A(n_3924),
.Y(n_4449)
);

OAI22xp33_ASAP7_75t_L g4450 ( 
.A1(n_3845),
.A2(n_2576),
.B1(n_2416),
.B2(n_2431),
.Y(n_4450)
);

AO32x2_ASAP7_75t_L g4451 ( 
.A1(n_3954),
.A2(n_3176),
.A3(n_3220),
.B1(n_3236),
.B2(n_3175),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_3681),
.Y(n_4452)
);

INVx2_ASAP7_75t_L g4453 ( 
.A(n_3665),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_3665),
.Y(n_4454)
);

NAND3xp33_ASAP7_75t_L g4455 ( 
.A(n_3549),
.B(n_3412),
.C(n_3396),
.Y(n_4455)
);

O2A1O1Ixp33_ASAP7_75t_SL g4456 ( 
.A1(n_3514),
.A2(n_2358),
.B(n_2412),
.C(n_3375),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_3763),
.B(n_3155),
.Y(n_4457)
);

OR2x2_ASAP7_75t_L g4458 ( 
.A(n_3767),
.B(n_3236),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_3634),
.B(n_3155),
.Y(n_4459)
);

INVx2_ASAP7_75t_L g4460 ( 
.A(n_3690),
.Y(n_4460)
);

OAI22xp33_ASAP7_75t_L g4461 ( 
.A1(n_3845),
.A2(n_2562),
.B1(n_2416),
.B2(n_2431),
.Y(n_4461)
);

OAI21x1_ASAP7_75t_L g4462 ( 
.A1(n_3636),
.A2(n_2529),
.B(n_2607),
.Y(n_4462)
);

OAI22xp5_ASAP7_75t_L g4463 ( 
.A1(n_3444),
.A2(n_3412),
.B1(n_3396),
.B2(n_3375),
.Y(n_4463)
);

INVx2_ASAP7_75t_L g4464 ( 
.A(n_3690),
.Y(n_4464)
);

CKINVDCx11_ASAP7_75t_R g4465 ( 
.A(n_3687),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_3692),
.Y(n_4466)
);

NAND2x1p5_ASAP7_75t_L g4467 ( 
.A(n_3682),
.B(n_2334),
.Y(n_4467)
);

AO32x2_ASAP7_75t_L g4468 ( 
.A1(n_3933),
.A2(n_3375),
.A3(n_3301),
.B1(n_3155),
.B2(n_3168),
.Y(n_4468)
);

BUFx4f_ASAP7_75t_SL g4469 ( 
.A(n_3493),
.Y(n_4469)
);

AO32x2_ASAP7_75t_L g4470 ( 
.A1(n_3978),
.A2(n_3301),
.A3(n_3240),
.B1(n_3155),
.B2(n_3168),
.Y(n_4470)
);

O2A1O1Ixp33_ASAP7_75t_SL g4471 ( 
.A1(n_3855),
.A2(n_2412),
.B(n_2358),
.C(n_3214),
.Y(n_4471)
);

O2A1O1Ixp33_ASAP7_75t_SL g4472 ( 
.A1(n_3891),
.A2(n_2412),
.B(n_2358),
.C(n_3214),
.Y(n_4472)
);

O2A1O1Ixp33_ASAP7_75t_L g4473 ( 
.A1(n_3509),
.A2(n_2478),
.B(n_2273),
.C(n_2274),
.Y(n_4473)
);

NOR2xp33_ASAP7_75t_L g4474 ( 
.A(n_3767),
.B(n_3168),
.Y(n_4474)
);

HB1xp67_ASAP7_75t_L g4475 ( 
.A(n_3963),
.Y(n_4475)
);

BUFx4f_ASAP7_75t_SL g4476 ( 
.A(n_3493),
.Y(n_4476)
);

O2A1O1Ixp33_ASAP7_75t_SL g4477 ( 
.A1(n_3960),
.A2(n_3301),
.B(n_3168),
.C(n_3175),
.Y(n_4477)
);

O2A1O1Ixp33_ASAP7_75t_SL g4478 ( 
.A1(n_3917),
.A2(n_3301),
.B(n_3168),
.C(n_3175),
.Y(n_4478)
);

CKINVDCx16_ASAP7_75t_R g4479 ( 
.A(n_3885),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_3769),
.B(n_3168),
.Y(n_4480)
);

INVx2_ASAP7_75t_L g4481 ( 
.A(n_3690),
.Y(n_4481)
);

O2A1O1Ixp5_ASAP7_75t_L g4482 ( 
.A1(n_3509),
.A2(n_2480),
.B(n_2283),
.C(n_2285),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_3692),
.Y(n_4483)
);

CKINVDCx20_ASAP7_75t_R g4484 ( 
.A(n_3493),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_3769),
.B(n_3175),
.Y(n_4485)
);

AOI22xp33_ASAP7_75t_L g4486 ( 
.A1(n_3901),
.A2(n_3663),
.B1(n_3724),
.B2(n_3697),
.Y(n_4486)
);

O2A1O1Ixp33_ASAP7_75t_SL g4487 ( 
.A1(n_3977),
.A2(n_3301),
.B(n_3175),
.C(n_3201),
.Y(n_4487)
);

A2O1A1Ixp33_ASAP7_75t_L g4488 ( 
.A1(n_3784),
.A2(n_2565),
.B(n_2598),
.C(n_2576),
.Y(n_4488)
);

A2O1A1Ixp33_ASAP7_75t_L g4489 ( 
.A1(n_3518),
.A2(n_2565),
.B(n_2598),
.C(n_2576),
.Y(n_4489)
);

NOR2x1_ASAP7_75t_SL g4490 ( 
.A(n_3892),
.B(n_3175),
.Y(n_4490)
);

INVx2_ASAP7_75t_L g4491 ( 
.A(n_3752),
.Y(n_4491)
);

NOR2xp67_ASAP7_75t_L g4492 ( 
.A(n_3682),
.B(n_3240),
.Y(n_4492)
);

BUFx3_ASAP7_75t_L g4493 ( 
.A(n_3673),
.Y(n_4493)
);

OAI22xp5_ASAP7_75t_L g4494 ( 
.A1(n_3491),
.A2(n_3240),
.B1(n_3223),
.B2(n_3214),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_3725),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_3771),
.B(n_3201),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_L g4497 ( 
.A(n_3771),
.B(n_3201),
.Y(n_4497)
);

O2A1O1Ixp33_ASAP7_75t_SL g4498 ( 
.A1(n_3977),
.A2(n_3240),
.B(n_3201),
.C(n_3203),
.Y(n_4498)
);

AOI22xp5_ASAP7_75t_L g4499 ( 
.A1(n_3511),
.A2(n_2261),
.B1(n_2592),
.B2(n_2563),
.Y(n_4499)
);

AOI22xp33_ASAP7_75t_L g4500 ( 
.A1(n_3663),
.A2(n_2285),
.B1(n_2286),
.B2(n_2297),
.Y(n_4500)
);

OAI22xp33_ASAP7_75t_L g4501 ( 
.A1(n_3892),
.A2(n_2591),
.B1(n_2474),
.B2(n_2501),
.Y(n_4501)
);

AOI22xp5_ASAP7_75t_L g4502 ( 
.A1(n_3552),
.A2(n_2592),
.B1(n_2563),
.B2(n_2562),
.Y(n_4502)
);

AO31x2_ASAP7_75t_L g4503 ( 
.A1(n_3562),
.A2(n_2529),
.A3(n_2623),
.B(n_2611),
.Y(n_4503)
);

INVx2_ASAP7_75t_SL g4504 ( 
.A(n_3929),
.Y(n_4504)
);

O2A1O1Ixp33_ASAP7_75t_SL g4505 ( 
.A1(n_3978),
.A2(n_3240),
.B(n_3223),
.C(n_3214),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_3725),
.Y(n_4506)
);

AO31x2_ASAP7_75t_L g4507 ( 
.A1(n_3581),
.A2(n_2614),
.A3(n_2623),
.B(n_2611),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_3774),
.B(n_3201),
.Y(n_4508)
);

BUFx6f_ASAP7_75t_L g4509 ( 
.A(n_3515),
.Y(n_4509)
);

AOI22xp33_ASAP7_75t_L g4510 ( 
.A1(n_3663),
.A2(n_3631),
.B1(n_3473),
.B2(n_3721),
.Y(n_4510)
);

OAI22x1_ASAP7_75t_L g4511 ( 
.A1(n_3510),
.A2(n_2286),
.B1(n_2297),
.B2(n_2301),
.Y(n_4511)
);

OAI21x1_ASAP7_75t_L g4512 ( 
.A1(n_3636),
.A2(n_2795),
.B(n_2614),
.Y(n_4512)
);

AOI22xp33_ASAP7_75t_L g4513 ( 
.A1(n_3663),
.A2(n_2301),
.B1(n_2303),
.B2(n_2306),
.Y(n_4513)
);

NOR2xp67_ASAP7_75t_SL g4514 ( 
.A(n_3452),
.B(n_2334),
.Y(n_4514)
);

OAI22xp33_ASAP7_75t_L g4515 ( 
.A1(n_3721),
.A2(n_2565),
.B1(n_2474),
.B2(n_2448),
.Y(n_4515)
);

INVx5_ASAP7_75t_L g4516 ( 
.A(n_3721),
.Y(n_4516)
);

INVx1_ASAP7_75t_SL g4517 ( 
.A(n_3872),
.Y(n_4517)
);

INVx2_ASAP7_75t_SL g4518 ( 
.A(n_3929),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_3730),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_3774),
.B(n_3201),
.Y(n_4520)
);

CKINVDCx11_ASAP7_75t_R g4521 ( 
.A(n_3909),
.Y(n_4521)
);

O2A1O1Ixp5_ASAP7_75t_L g4522 ( 
.A1(n_3651),
.A2(n_3921),
.B(n_3688),
.C(n_3987),
.Y(n_4522)
);

INVx5_ASAP7_75t_SL g4523 ( 
.A(n_3527),
.Y(n_4523)
);

AND2x2_ASAP7_75t_L g4524 ( 
.A(n_3712),
.B(n_3203),
.Y(n_4524)
);

OAI22xp33_ASAP7_75t_L g4525 ( 
.A1(n_3721),
.A2(n_2565),
.B1(n_2474),
.B2(n_2448),
.Y(n_4525)
);

INVxp67_ASAP7_75t_L g4526 ( 
.A(n_3568),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_3695),
.B(n_3203),
.Y(n_4527)
);

OAI22xp5_ASAP7_75t_L g4528 ( 
.A1(n_3936),
.A2(n_3223),
.B1(n_3206),
.B2(n_3203),
.Y(n_4528)
);

BUFx2_ASAP7_75t_L g4529 ( 
.A(n_3525),
.Y(n_4529)
);

INVx2_ASAP7_75t_L g4530 ( 
.A(n_3752),
.Y(n_4530)
);

O2A1O1Ixp33_ASAP7_75t_SL g4531 ( 
.A1(n_3453),
.A2(n_3223),
.B(n_3206),
.C(n_3203),
.Y(n_4531)
);

AO31x2_ASAP7_75t_L g4532 ( 
.A1(n_3629),
.A2(n_2637),
.A3(n_2623),
.B(n_2614),
.Y(n_4532)
);

A2O1A1Ixp33_ASAP7_75t_L g4533 ( 
.A1(n_3629),
.A2(n_2562),
.B(n_2604),
.C(n_2598),
.Y(n_4533)
);

AND2x2_ASAP7_75t_L g4534 ( 
.A(n_3712),
.B(n_3203),
.Y(n_4534)
);

NOR2xp33_ASAP7_75t_L g4535 ( 
.A(n_3956),
.B(n_3206),
.Y(n_4535)
);

A2O1A1Ixp33_ASAP7_75t_L g4536 ( 
.A1(n_3839),
.A2(n_3813),
.B(n_3974),
.C(n_3814),
.Y(n_4536)
);

AOI22xp5_ASAP7_75t_L g4537 ( 
.A1(n_3488),
.A2(n_2592),
.B1(n_2562),
.B2(n_2604),
.Y(n_4537)
);

AOI22xp33_ASAP7_75t_L g4538 ( 
.A1(n_3473),
.A2(n_2324),
.B1(n_2350),
.B2(n_2352),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_3730),
.Y(n_4539)
);

INVx3_ASAP7_75t_L g4540 ( 
.A(n_3515),
.Y(n_4540)
);

AOI21xp5_ASAP7_75t_SL g4541 ( 
.A1(n_3967),
.A2(n_3979),
.B(n_3893),
.Y(n_4541)
);

A2O1A1Ixp33_ASAP7_75t_L g4542 ( 
.A1(n_3974),
.A2(n_2576),
.B(n_2604),
.C(n_2598),
.Y(n_4542)
);

AOI22xp33_ASAP7_75t_L g4543 ( 
.A1(n_3473),
.A2(n_2350),
.B1(n_2352),
.B2(n_2353),
.Y(n_4543)
);

INVx2_ASAP7_75t_L g4544 ( 
.A(n_3752),
.Y(n_4544)
);

INVx2_ASAP7_75t_L g4545 ( 
.A(n_3761),
.Y(n_4545)
);

BUFx6f_ASAP7_75t_L g4546 ( 
.A(n_3515),
.Y(n_4546)
);

AO31x2_ASAP7_75t_L g4547 ( 
.A1(n_3926),
.A2(n_2644),
.A3(n_2637),
.B(n_2839),
.Y(n_4547)
);

O2A1O1Ixp33_ASAP7_75t_SL g4548 ( 
.A1(n_3453),
.A2(n_3223),
.B(n_3206),
.C(n_2567),
.Y(n_4548)
);

AND2x4_ASAP7_75t_L g4549 ( 
.A(n_3628),
.B(n_3206),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_3735),
.Y(n_4550)
);

AO31x2_ASAP7_75t_L g4551 ( 
.A1(n_3770),
.A2(n_2839),
.A3(n_2826),
.B(n_2821),
.Y(n_4551)
);

HB1xp67_ASAP7_75t_L g4552 ( 
.A(n_3971),
.Y(n_4552)
);

CKINVDCx5p33_ASAP7_75t_R g4553 ( 
.A(n_3673),
.Y(n_4553)
);

INVx2_ASAP7_75t_SL g4554 ( 
.A(n_3909),
.Y(n_4554)
);

CKINVDCx6p67_ASAP7_75t_R g4555 ( 
.A(n_3909),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_3735),
.Y(n_4556)
);

AOI21xp5_ASAP7_75t_L g4557 ( 
.A1(n_3666),
.A2(n_3676),
.B(n_3773),
.Y(n_4557)
);

OAI21x1_ASAP7_75t_L g4558 ( 
.A1(n_3719),
.A2(n_2731),
.B(n_2826),
.Y(n_4558)
);

CKINVDCx11_ASAP7_75t_R g4559 ( 
.A(n_3673),
.Y(n_4559)
);

AOI31xp67_ASAP7_75t_L g4560 ( 
.A1(n_3761),
.A2(n_2839),
.A3(n_2826),
.B(n_2821),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_3695),
.B(n_2612),
.Y(n_4561)
);

BUFx10_ASAP7_75t_L g4562 ( 
.A(n_3515),
.Y(n_4562)
);

BUFx6f_ASAP7_75t_L g4563 ( 
.A(n_3515),
.Y(n_4563)
);

CKINVDCx9p33_ASAP7_75t_R g4564 ( 
.A(n_3556),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_3746),
.Y(n_4565)
);

O2A1O1Ixp33_ASAP7_75t_SL g4566 ( 
.A1(n_3460),
.A2(n_2567),
.B(n_2479),
.C(n_2371),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_3746),
.Y(n_4567)
);

AOI22xp33_ASAP7_75t_L g4568 ( 
.A1(n_3631),
.A2(n_2353),
.B1(n_2360),
.B2(n_2535),
.Y(n_4568)
);

OR2x2_ASAP7_75t_L g4569 ( 
.A(n_3698),
.B(n_2577),
.Y(n_4569)
);

NAND3xp33_ASAP7_75t_L g4570 ( 
.A(n_3790),
.B(n_2612),
.C(n_2647),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_3765),
.Y(n_4571)
);

BUFx6f_ASAP7_75t_L g4572 ( 
.A(n_3515),
.Y(n_4572)
);

OR2x6_ASAP7_75t_L g4573 ( 
.A(n_3700),
.B(n_2416),
.Y(n_4573)
);

AND2x2_ASAP7_75t_L g4574 ( 
.A(n_3727),
.B(n_2612),
.Y(n_4574)
);

NOR2xp33_ASAP7_75t_SL g4575 ( 
.A(n_3474),
.B(n_2371),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_3727),
.B(n_2612),
.Y(n_4576)
);

HB1xp67_ASAP7_75t_L g4577 ( 
.A(n_4552),
.Y(n_4577)
);

BUFx3_ASAP7_75t_L g4578 ( 
.A(n_4364),
.Y(n_4578)
);

A2O1A1Ixp33_ASAP7_75t_L g4579 ( 
.A1(n_3996),
.A2(n_3980),
.B(n_3556),
.C(n_3982),
.Y(n_4579)
);

AND2x4_ASAP7_75t_L g4580 ( 
.A(n_4490),
.B(n_3628),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4468),
.B(n_3569),
.Y(n_4581)
);

HB1xp67_ASAP7_75t_L g4582 ( 
.A(n_4373),
.Y(n_4582)
);

AOI21xp5_ASAP7_75t_L g4583 ( 
.A1(n_4169),
.A2(n_3816),
.B(n_3804),
.Y(n_4583)
);

OAI21x1_ASAP7_75t_SL g4584 ( 
.A1(n_4024),
.A2(n_3894),
.B(n_3879),
.Y(n_4584)
);

BUFx12f_ASAP7_75t_L g4585 ( 
.A(n_4065),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4468),
.B(n_3569),
.Y(n_4586)
);

HB1xp67_ASAP7_75t_L g4587 ( 
.A(n_4170),
.Y(n_4587)
);

INVx3_ASAP7_75t_L g4588 ( 
.A(n_4549),
.Y(n_4588)
);

AOI21xp5_ASAP7_75t_L g4589 ( 
.A1(n_4169),
.A2(n_3816),
.B(n_3804),
.Y(n_4589)
);

INVxp67_ASAP7_75t_L g4590 ( 
.A(n_4074),
.Y(n_4590)
);

AO21x2_ASAP7_75t_L g4591 ( 
.A1(n_4028),
.A2(n_3584),
.B(n_3600),
.Y(n_4591)
);

HB1xp67_ASAP7_75t_L g4592 ( 
.A(n_4240),
.Y(n_4592)
);

BUFx2_ASAP7_75t_L g4593 ( 
.A(n_4357),
.Y(n_4593)
);

NAND2x1p5_ASAP7_75t_L g4594 ( 
.A(n_4181),
.B(n_3721),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4011),
.Y(n_4595)
);

OAI21xp5_ASAP7_75t_L g4596 ( 
.A1(n_4000),
.A2(n_3707),
.B(n_3861),
.Y(n_4596)
);

INVx1_ASAP7_75t_SL g4597 ( 
.A(n_4446),
.Y(n_4597)
);

INVx2_ASAP7_75t_L g4598 ( 
.A(n_4444),
.Y(n_4598)
);

INVx2_ASAP7_75t_L g4599 ( 
.A(n_4444),
.Y(n_4599)
);

AND2x4_ASAP7_75t_L g4600 ( 
.A(n_4490),
.B(n_4165),
.Y(n_4600)
);

OAI21xp5_ASAP7_75t_L g4601 ( 
.A1(n_4177),
.A2(n_3861),
.B(n_3532),
.Y(n_4601)
);

AO21x2_ASAP7_75t_L g4602 ( 
.A1(n_4028),
.A2(n_3584),
.B(n_3600),
.Y(n_4602)
);

AND2x4_ASAP7_75t_L g4603 ( 
.A(n_4165),
.B(n_3639),
.Y(n_4603)
);

OAI21x1_ASAP7_75t_L g4604 ( 
.A1(n_4226),
.A2(n_3662),
.B(n_3654),
.Y(n_4604)
);

NOR2xp67_ASAP7_75t_L g4605 ( 
.A(n_4157),
.B(n_3721),
.Y(n_4605)
);

AOI21x1_ASAP7_75t_L g4606 ( 
.A1(n_4280),
.A2(n_4226),
.B(n_4201),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4011),
.Y(n_4607)
);

A2O1A1Ixp33_ASAP7_75t_L g4608 ( 
.A1(n_4135),
.A2(n_3980),
.B(n_3982),
.C(n_3474),
.Y(n_4608)
);

OAI22xp5_ASAP7_75t_L g4609 ( 
.A1(n_4135),
.A2(n_3790),
.B1(n_3918),
.B2(n_3698),
.Y(n_4609)
);

AO21x2_ASAP7_75t_L g4610 ( 
.A1(n_4217),
.A2(n_3584),
.B(n_3600),
.Y(n_4610)
);

AO21x2_ASAP7_75t_L g4611 ( 
.A1(n_4217),
.A2(n_3584),
.B(n_3600),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4468),
.B(n_3569),
.Y(n_4612)
);

AOI21xp5_ASAP7_75t_L g4613 ( 
.A1(n_4369),
.A2(n_3816),
.B(n_3532),
.Y(n_4613)
);

NOR2xp33_ASAP7_75t_L g4614 ( 
.A(n_4379),
.B(n_3487),
.Y(n_4614)
);

AOI21x1_ASAP7_75t_L g4615 ( 
.A1(n_4201),
.A2(n_3555),
.B(n_3722),
.Y(n_4615)
);

OAI21x1_ASAP7_75t_L g4616 ( 
.A1(n_4292),
.A2(n_4066),
.B(n_4057),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4045),
.Y(n_4617)
);

OR2x6_ASAP7_75t_L g4618 ( 
.A(n_4181),
.B(n_4127),
.Y(n_4618)
);

OAI21x1_ASAP7_75t_L g4619 ( 
.A1(n_4057),
.A2(n_3555),
.B(n_3639),
.Y(n_4619)
);

OAI21x1_ASAP7_75t_L g4620 ( 
.A1(n_4066),
.A2(n_3722),
.B(n_3446),
.Y(n_4620)
);

AO21x2_ASAP7_75t_L g4621 ( 
.A1(n_4252),
.A2(n_3938),
.B(n_3540),
.Y(n_4621)
);

INVx4_ASAP7_75t_L g4622 ( 
.A(n_4326),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_L g4623 ( 
.A(n_4202),
.B(n_3572),
.Y(n_4623)
);

INVx6_ASAP7_75t_L g4624 ( 
.A(n_4041),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4045),
.Y(n_4625)
);

AO21x2_ASAP7_75t_L g4626 ( 
.A1(n_4073),
.A2(n_3938),
.B(n_3540),
.Y(n_4626)
);

BUFx8_ASAP7_75t_SL g4627 ( 
.A(n_4040),
.Y(n_4627)
);

AOI22x1_ASAP7_75t_L g4628 ( 
.A1(n_4043),
.A2(n_4322),
.B1(n_4127),
.B2(n_4479),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4075),
.Y(n_4629)
);

HB1xp67_ASAP7_75t_L g4630 ( 
.A(n_4318),
.Y(n_4630)
);

OAI21x1_ASAP7_75t_L g4631 ( 
.A1(n_4557),
.A2(n_3736),
.B(n_3458),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4212),
.B(n_4225),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4075),
.Y(n_4633)
);

INVx1_ASAP7_75t_SL g4634 ( 
.A(n_4564),
.Y(n_4634)
);

OAI21xp5_ASAP7_75t_L g4635 ( 
.A1(n_4048),
.A2(n_3477),
.B(n_3785),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4088),
.Y(n_4636)
);

NAND3xp33_ASAP7_75t_L g4637 ( 
.A(n_4379),
.B(n_3477),
.C(n_3466),
.Y(n_4637)
);

AO31x2_ASAP7_75t_L g4638 ( 
.A1(n_4335),
.A2(n_3877),
.A3(n_3873),
.B(n_3779),
.Y(n_4638)
);

AND2x4_ASAP7_75t_L g4639 ( 
.A(n_4165),
.B(n_3992),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4468),
.B(n_3569),
.Y(n_4640)
);

AO21x1_ASAP7_75t_L g4641 ( 
.A1(n_4039),
.A2(n_3489),
.B(n_3487),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_L g4642 ( 
.A(n_4278),
.B(n_3572),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_4279),
.B(n_4429),
.Y(n_4643)
);

NOR2xp33_ASAP7_75t_L g4644 ( 
.A(n_4347),
.B(n_3489),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_4444),
.Y(n_4645)
);

OAI21x1_ASAP7_75t_L g4646 ( 
.A1(n_4325),
.A2(n_3578),
.B(n_3756),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4088),
.Y(n_4647)
);

AO21x2_ASAP7_75t_L g4648 ( 
.A1(n_4335),
.A2(n_3938),
.B(n_3540),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_4444),
.Y(n_4649)
);

OAI21x1_ASAP7_75t_L g4650 ( 
.A1(n_4214),
.A2(n_3778),
.B(n_3772),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4101),
.Y(n_4651)
);

AO31x2_ASAP7_75t_L g4652 ( 
.A1(n_4182),
.A2(n_4275),
.A3(n_4366),
.B(n_4511),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4101),
.Y(n_4653)
);

OAI22xp5_ASAP7_75t_L g4654 ( 
.A1(n_4168),
.A2(n_3918),
.B1(n_3699),
.B2(n_3858),
.Y(n_4654)
);

OR2x2_ASAP7_75t_L g4655 ( 
.A(n_4442),
.B(n_3971),
.Y(n_4655)
);

OAI21x1_ASAP7_75t_L g4656 ( 
.A1(n_4214),
.A2(n_3772),
.B(n_3745),
.Y(n_4656)
);

INVx2_ASAP7_75t_SL g4657 ( 
.A(n_4364),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4102),
.Y(n_4658)
);

INVx3_ASAP7_75t_L g4659 ( 
.A(n_4549),
.Y(n_4659)
);

OR2x2_ASAP7_75t_L g4660 ( 
.A(n_4044),
.B(n_3985),
.Y(n_4660)
);

BUFx3_ASAP7_75t_L g4661 ( 
.A(n_4364),
.Y(n_4661)
);

OAI21x1_ASAP7_75t_L g4662 ( 
.A1(n_4214),
.A2(n_4282),
.B(n_4291),
.Y(n_4662)
);

NOR2x1_ASAP7_75t_SL g4663 ( 
.A(n_4228),
.B(n_3879),
.Y(n_4663)
);

HB1xp67_ASAP7_75t_L g4664 ( 
.A(n_4435),
.Y(n_4664)
);

BUFx2_ASAP7_75t_R g4665 ( 
.A(n_3995),
.Y(n_4665)
);

OR2x6_ASAP7_75t_L g4666 ( 
.A(n_4035),
.B(n_3700),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4014),
.B(n_3575),
.Y(n_4667)
);

OAI21x1_ASAP7_75t_L g4668 ( 
.A1(n_4282),
.A2(n_3838),
.B(n_3831),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4102),
.Y(n_4669)
);

INVx2_ASAP7_75t_L g4670 ( 
.A(n_4444),
.Y(n_4670)
);

BUFx2_ASAP7_75t_SL g4671 ( 
.A(n_4492),
.Y(n_4671)
);

BUFx6f_ASAP7_75t_L g4672 ( 
.A(n_4468),
.Y(n_4672)
);

AND2x4_ASAP7_75t_L g4673 ( 
.A(n_4165),
.B(n_3992),
.Y(n_4673)
);

OA21x2_ASAP7_75t_L g4674 ( 
.A1(n_4275),
.A2(n_4377),
.B(n_4533),
.Y(n_4674)
);

NOR2xp33_ASAP7_75t_L g4675 ( 
.A(n_4019),
.B(n_3460),
.Y(n_4675)
);

AND2x2_ASAP7_75t_L g4676 ( 
.A(n_4470),
.B(n_3569),
.Y(n_4676)
);

OR2x6_ASAP7_75t_L g4677 ( 
.A(n_4035),
.B(n_3700),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4117),
.Y(n_4678)
);

NOR2xp33_ASAP7_75t_L g4679 ( 
.A(n_4032),
.B(n_3466),
.Y(n_4679)
);

AOI21xp5_ASAP7_75t_L g4680 ( 
.A1(n_4541),
.A2(n_3816),
.B(n_3747),
.Y(n_4680)
);

INVx4_ASAP7_75t_L g4681 ( 
.A(n_4326),
.Y(n_4681)
);

BUFx2_ASAP7_75t_R g4682 ( 
.A(n_3995),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4029),
.B(n_3575),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4526),
.B(n_3492),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4117),
.Y(n_4685)
);

AND2x4_ASAP7_75t_L g4686 ( 
.A(n_4046),
.B(n_4047),
.Y(n_4686)
);

HB1xp67_ASAP7_75t_L g4687 ( 
.A(n_4475),
.Y(n_4687)
);

HB1xp67_ASAP7_75t_L g4688 ( 
.A(n_4105),
.Y(n_4688)
);

HB1xp67_ASAP7_75t_L g4689 ( 
.A(n_4105),
.Y(n_4689)
);

INVx2_ASAP7_75t_L g4690 ( 
.A(n_4451),
.Y(n_4690)
);

BUFx4f_ASAP7_75t_SL g4691 ( 
.A(n_4040),
.Y(n_4691)
);

OAI21x1_ASAP7_75t_SL g4692 ( 
.A1(n_4431),
.A2(n_3894),
.B(n_3824),
.Y(n_4692)
);

OAI22xp5_ASAP7_75t_L g4693 ( 
.A1(n_4168),
.A2(n_3699),
.B1(n_3858),
.B2(n_3760),
.Y(n_4693)
);

NAND2x1p5_ASAP7_75t_L g4694 ( 
.A(n_4205),
.B(n_3709),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4054),
.B(n_3492),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4121),
.Y(n_4696)
);

NAND2x1p5_ASAP7_75t_L g4697 ( 
.A(n_4205),
.B(n_3709),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4451),
.Y(n_4698)
);

NOR2x1_ASAP7_75t_SL g4699 ( 
.A(n_4207),
.B(n_3566),
.Y(n_4699)
);

CKINVDCx5p33_ASAP7_75t_R g4700 ( 
.A(n_4064),
.Y(n_4700)
);

AO21x2_ASAP7_75t_L g4701 ( 
.A1(n_4558),
.A2(n_3938),
.B(n_3540),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4121),
.Y(n_4702)
);

AND2x2_ASAP7_75t_L g4703 ( 
.A(n_4470),
.B(n_3739),
.Y(n_4703)
);

CKINVDCx20_ASAP7_75t_R g4704 ( 
.A(n_4091),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4131),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4131),
.Y(n_4706)
);

INVx4_ASAP7_75t_L g4707 ( 
.A(n_4555),
.Y(n_4707)
);

OAI21x1_ASAP7_75t_SL g4708 ( 
.A1(n_4431),
.A2(n_3824),
.B(n_3576),
.Y(n_4708)
);

OAI21xp5_ASAP7_75t_L g4709 ( 
.A1(n_4122),
.A2(n_3477),
.B(n_3785),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4274),
.B(n_4294),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4314),
.B(n_3502),
.Y(n_4711)
);

AND2x4_ASAP7_75t_L g4712 ( 
.A(n_4046),
.B(n_3655),
.Y(n_4712)
);

OAI21xp5_ASAP7_75t_L g4713 ( 
.A1(n_4210),
.A2(n_3477),
.B(n_3785),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4154),
.Y(n_4714)
);

BUFx2_ASAP7_75t_R g4715 ( 
.A(n_4012),
.Y(n_4715)
);

AOI22xp33_ASAP7_75t_L g4716 ( 
.A1(n_3997),
.A2(n_3785),
.B1(n_3527),
.B2(n_3686),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4451),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4154),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4451),
.Y(n_4719)
);

NAND2x1p5_ASAP7_75t_L g4720 ( 
.A(n_4205),
.B(n_3782),
.Y(n_4720)
);

INVx2_ASAP7_75t_SL g4721 ( 
.A(n_4364),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4171),
.Y(n_4722)
);

A2O1A1Ixp33_ASAP7_75t_L g4723 ( 
.A1(n_4030),
.A2(n_4198),
.B(n_4153),
.C(n_4536),
.Y(n_4723)
);

NAND2x1p5_ASAP7_75t_L g4724 ( 
.A(n_4205),
.B(n_3782),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4171),
.Y(n_4725)
);

OAI21xp5_ASAP7_75t_L g4726 ( 
.A1(n_4023),
.A2(n_3468),
.B(n_3467),
.Y(n_4726)
);

BUFx6f_ASAP7_75t_L g4727 ( 
.A(n_4470),
.Y(n_4727)
);

AO22x2_ASAP7_75t_L g4728 ( 
.A1(n_4251),
.A2(n_4157),
.B1(n_4085),
.B2(n_4112),
.Y(n_4728)
);

INVx2_ASAP7_75t_L g4729 ( 
.A(n_4451),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4172),
.Y(n_4730)
);

AOI21x1_ASAP7_75t_L g4731 ( 
.A1(n_4549),
.A2(n_3768),
.B(n_3940),
.Y(n_4731)
);

HB1xp67_ASAP7_75t_L g4732 ( 
.A(n_4230),
.Y(n_4732)
);

INVx2_ASAP7_75t_L g4733 ( 
.A(n_4560),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4172),
.Y(n_4734)
);

AOI21xp5_ASAP7_75t_L g4735 ( 
.A1(n_4541),
.A2(n_3965),
.B(n_3952),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4173),
.Y(n_4736)
);

INVx3_ASAP7_75t_L g4737 ( 
.A(n_4211),
.Y(n_4737)
);

AND2x2_ASAP7_75t_L g4738 ( 
.A(n_4470),
.B(n_3739),
.Y(n_4738)
);

AND2x2_ASAP7_75t_L g4739 ( 
.A(n_4470),
.B(n_3760),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4560),
.Y(n_4740)
);

AO31x2_ASAP7_75t_L g4741 ( 
.A1(n_4097),
.A2(n_3843),
.A3(n_3852),
.B(n_3829),
.Y(n_4741)
);

INVx2_ASAP7_75t_L g4742 ( 
.A(n_4211),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4173),
.Y(n_4743)
);

AOI21xp5_ASAP7_75t_L g4744 ( 
.A1(n_4114),
.A2(n_3973),
.B(n_3972),
.Y(n_4744)
);

AND2x4_ASAP7_75t_L g4745 ( 
.A(n_4046),
.B(n_3655),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4176),
.Y(n_4746)
);

BUFx8_ASAP7_75t_L g4747 ( 
.A(n_4188),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4067),
.B(n_3502),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4176),
.Y(n_4749)
);

HB1xp67_ASAP7_75t_L g4750 ( 
.A(n_4230),
.Y(n_4750)
);

NAND2x1p5_ASAP7_75t_L g4751 ( 
.A(n_4205),
.B(n_3944),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_L g4752 ( 
.A(n_4053),
.B(n_3506),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4183),
.Y(n_4753)
);

HB1xp67_ASAP7_75t_L g4754 ( 
.A(n_4231),
.Y(n_4754)
);

OAI22xp5_ASAP7_75t_L g4755 ( 
.A1(n_4023),
.A2(n_3916),
.B1(n_3543),
.B2(n_3563),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4357),
.B(n_3494),
.Y(n_4756)
);

INVx2_ASAP7_75t_L g4757 ( 
.A(n_4211),
.Y(n_4757)
);

AO21x2_ASAP7_75t_L g4758 ( 
.A1(n_4558),
.A2(n_4260),
.B(n_4256),
.Y(n_4758)
);

NOR2xp33_ASAP7_75t_L g4759 ( 
.A(n_4018),
.B(n_4139),
.Y(n_4759)
);

INVx1_ASAP7_75t_SL g4760 ( 
.A(n_4400),
.Y(n_4760)
);

HB1xp67_ASAP7_75t_L g4761 ( 
.A(n_4231),
.Y(n_4761)
);

BUFx6f_ASAP7_75t_L g4762 ( 
.A(n_4205),
.Y(n_4762)
);

AND2x4_ASAP7_75t_L g4763 ( 
.A(n_4046),
.B(n_3655),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4183),
.Y(n_4764)
);

NOR2xp67_ASAP7_75t_L g4765 ( 
.A(n_4157),
.B(n_3448),
.Y(n_4765)
);

INVx1_ASAP7_75t_SL g4766 ( 
.A(n_4400),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4078),
.B(n_3506),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4187),
.Y(n_4768)
);

INVx6_ASAP7_75t_L g4769 ( 
.A(n_4041),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4187),
.Y(n_4770)
);

OAI21xp5_ASAP7_75t_L g4771 ( 
.A1(n_4027),
.A2(n_3468),
.B(n_3467),
.Y(n_4771)
);

CKINVDCx11_ASAP7_75t_R g4772 ( 
.A(n_4091),
.Y(n_4772)
);

AOI21xp5_ASAP7_75t_L g4773 ( 
.A1(n_4080),
.A2(n_4505),
.B(n_4381),
.Y(n_4773)
);

INVxp67_ASAP7_75t_L g4774 ( 
.A(n_4034),
.Y(n_4774)
);

CKINVDCx5p33_ASAP7_75t_R g4775 ( 
.A(n_4064),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4199),
.Y(n_4776)
);

OR2x2_ASAP7_75t_L g4777 ( 
.A(n_4404),
.B(n_3985),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4199),
.Y(n_4778)
);

A2O1A1Ixp33_ASAP7_75t_L g4779 ( 
.A1(n_4001),
.A2(n_3944),
.B(n_3528),
.C(n_3928),
.Y(n_4779)
);

OR2x2_ASAP7_75t_L g4780 ( 
.A(n_4517),
.B(n_3878),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4219),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4219),
.Y(n_4782)
);

BUFx2_ASAP7_75t_L g4783 ( 
.A(n_4357),
.Y(n_4783)
);

BUFx2_ASAP7_75t_L g4784 ( 
.A(n_4357),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4229),
.Y(n_4785)
);

OAI21xp5_ASAP7_75t_L g4786 ( 
.A1(n_4020),
.A2(n_3818),
.B(n_3811),
.Y(n_4786)
);

AOI21xp5_ASAP7_75t_L g4787 ( 
.A1(n_4033),
.A2(n_3768),
.B(n_3983),
.Y(n_4787)
);

NAND2x1p5_ASAP7_75t_L g4788 ( 
.A(n_4209),
.B(n_3452),
.Y(n_4788)
);

AO21x2_ASAP7_75t_L g4789 ( 
.A1(n_4112),
.A2(n_3527),
.B(n_3498),
.Y(n_4789)
);

NOR2xp67_ASAP7_75t_L g4790 ( 
.A(n_4097),
.B(n_3448),
.Y(n_4790)
);

OA21x2_ASAP7_75t_L g4791 ( 
.A1(n_4522),
.A2(n_4412),
.B(n_4482),
.Y(n_4791)
);

INVx2_ASAP7_75t_L g4792 ( 
.A(n_4211),
.Y(n_4792)
);

NOR2xp33_ASAP7_75t_L g4793 ( 
.A(n_4016),
.B(n_3568),
.Y(n_4793)
);

NOR2xp33_ASAP7_75t_L g4794 ( 
.A(n_4026),
.B(n_3571),
.Y(n_4794)
);

OA21x2_ASAP7_75t_L g4795 ( 
.A1(n_4455),
.A2(n_3729),
.B(n_3720),
.Y(n_4795)
);

OAI21xp5_ASAP7_75t_L g4796 ( 
.A1(n_4085),
.A2(n_3818),
.B(n_3811),
.Y(n_4796)
);

HB1xp67_ASAP7_75t_L g4797 ( 
.A(n_4253),
.Y(n_4797)
);

AOI21xp5_ASAP7_75t_L g4798 ( 
.A1(n_4033),
.A2(n_3768),
.B(n_3991),
.Y(n_4798)
);

INVx2_ASAP7_75t_L g4799 ( 
.A(n_4250),
.Y(n_4799)
);

CKINVDCx5p33_ASAP7_75t_R g4800 ( 
.A(n_4051),
.Y(n_4800)
);

AO21x2_ASAP7_75t_L g4801 ( 
.A1(n_4462),
.A2(n_3527),
.B(n_3498),
.Y(n_4801)
);

BUFx2_ASAP7_75t_L g4802 ( 
.A(n_4357),
.Y(n_4802)
);

AO31x2_ASAP7_75t_L g4803 ( 
.A1(n_4255),
.A2(n_3852),
.A3(n_3853),
.B(n_3843),
.Y(n_4803)
);

INVx3_ASAP7_75t_L g4804 ( 
.A(n_4250),
.Y(n_4804)
);

AOI21xp5_ASAP7_75t_L g4805 ( 
.A1(n_4033),
.A2(n_3768),
.B(n_3946),
.Y(n_4805)
);

AND2x4_ASAP7_75t_L g4806 ( 
.A(n_4047),
.B(n_3655),
.Y(n_4806)
);

NAND2x1p5_ASAP7_75t_L g4807 ( 
.A(n_4209),
.B(n_3452),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4229),
.Y(n_4808)
);

INVx3_ASAP7_75t_L g4809 ( 
.A(n_4250),
.Y(n_4809)
);

OAI21xp5_ASAP7_75t_L g4810 ( 
.A1(n_4100),
.A2(n_4081),
.B(n_4141),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4236),
.Y(n_4811)
);

HB1xp67_ASAP7_75t_L g4812 ( 
.A(n_4253),
.Y(n_4812)
);

CKINVDCx20_ASAP7_75t_R g4813 ( 
.A(n_4213),
.Y(n_4813)
);

AND2x2_ASAP7_75t_L g4814 ( 
.A(n_4206),
.B(n_3494),
.Y(n_4814)
);

INVx3_ASAP7_75t_L g4815 ( 
.A(n_4250),
.Y(n_4815)
);

OAI21xp5_ASAP7_75t_L g4816 ( 
.A1(n_4408),
.A2(n_4049),
.B(n_4007),
.Y(n_4816)
);

NOR2xp67_ASAP7_75t_L g4817 ( 
.A(n_4455),
.B(n_3448),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4206),
.B(n_3494),
.Y(n_4818)
);

AO21x2_ASAP7_75t_L g4819 ( 
.A1(n_4512),
.A2(n_4096),
.B(n_4197),
.Y(n_4819)
);

BUFx6f_ASAP7_75t_L g4820 ( 
.A(n_4209),
.Y(n_4820)
);

AO222x2_ASAP7_75t_SL g4821 ( 
.A1(n_4448),
.A2(n_3704),
.B1(n_3970),
.B2(n_3951),
.C1(n_3844),
.C2(n_3766),
.Y(n_4821)
);

AOI21xp5_ASAP7_75t_L g4822 ( 
.A1(n_4033),
.A2(n_3579),
.B(n_3914),
.Y(n_4822)
);

AOI21xp33_ASAP7_75t_SL g4823 ( 
.A1(n_4109),
.A2(n_3570),
.B(n_3499),
.Y(n_4823)
);

INVx2_ASAP7_75t_L g4824 ( 
.A(n_4405),
.Y(n_4824)
);

AND2x4_ASAP7_75t_L g4825 ( 
.A(n_4047),
.B(n_4186),
.Y(n_4825)
);

OR2x2_ASAP7_75t_L g4826 ( 
.A(n_4356),
.B(n_3878),
.Y(n_4826)
);

BUFx3_ASAP7_75t_L g4827 ( 
.A(n_4365),
.Y(n_4827)
);

OA21x2_ASAP7_75t_L g4828 ( 
.A1(n_4327),
.A2(n_3830),
.B(n_3781),
.Y(n_4828)
);

HB1xp67_ASAP7_75t_L g4829 ( 
.A(n_4258),
.Y(n_4829)
);

NOR2xp33_ASAP7_75t_L g4830 ( 
.A(n_4031),
.B(n_3571),
.Y(n_4830)
);

AOI22xp33_ASAP7_75t_L g4831 ( 
.A1(n_4264),
.A2(n_3680),
.B1(n_3631),
.B2(n_3815),
.Y(n_4831)
);

INVx3_ASAP7_75t_L g4832 ( 
.A(n_4405),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_L g4833 ( 
.A(n_4138),
.B(n_4345),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4236),
.Y(n_4834)
);

AO21x2_ASAP7_75t_L g4835 ( 
.A1(n_4570),
.A2(n_3864),
.B(n_3830),
.Y(n_4835)
);

BUFx6f_ASAP7_75t_L g4836 ( 
.A(n_4209),
.Y(n_4836)
);

AO21x2_ASAP7_75t_L g4837 ( 
.A1(n_4570),
.A2(n_3870),
.B(n_3864),
.Y(n_4837)
);

AOI21xp5_ASAP7_75t_L g4838 ( 
.A1(n_4146),
.A2(n_3579),
.B(n_3880),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_4234),
.B(n_3880),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4237),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4237),
.Y(n_4841)
);

NOR2xp33_ASAP7_75t_L g4842 ( 
.A(n_4060),
.B(n_3981),
.Y(n_4842)
);

INVx2_ASAP7_75t_L g4843 ( 
.A(n_4405),
.Y(n_4843)
);

AOI21x1_ASAP7_75t_L g4844 ( 
.A1(n_4083),
.A2(n_3630),
.B(n_3579),
.Y(n_4844)
);

INVx2_ASAP7_75t_L g4845 ( 
.A(n_4405),
.Y(n_4845)
);

AND2x4_ASAP7_75t_L g4846 ( 
.A(n_4047),
.B(n_3678),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4262),
.Y(n_4847)
);

NAND2x1p5_ASAP7_75t_L g4848 ( 
.A(n_4209),
.B(n_3452),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4262),
.Y(n_4849)
);

INVx2_ASAP7_75t_L g4850 ( 
.A(n_4443),
.Y(n_4850)
);

NOR2x1_ASAP7_75t_SL g4851 ( 
.A(n_4227),
.B(n_3576),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4276),
.Y(n_4852)
);

AO31x2_ASAP7_75t_L g4853 ( 
.A1(n_4255),
.A2(n_4082),
.A3(n_4488),
.B(n_4200),
.Y(n_4853)
);

OA21x2_ASAP7_75t_L g4854 ( 
.A1(n_4068),
.A2(n_3870),
.B(n_3864),
.Y(n_4854)
);

NAND2xp5_ASAP7_75t_L g4855 ( 
.A(n_4248),
.B(n_3889),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4017),
.B(n_4004),
.Y(n_4856)
);

AOI21xp5_ASAP7_75t_L g4857 ( 
.A1(n_4531),
.A2(n_3579),
.B(n_3889),
.Y(n_4857)
);

BUFx6f_ASAP7_75t_L g4858 ( 
.A(n_4209),
.Y(n_4858)
);

INVx2_ASAP7_75t_L g4859 ( 
.A(n_4443),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4319),
.B(n_3900),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4017),
.B(n_3494),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4276),
.Y(n_4862)
);

NOR2xp67_ASAP7_75t_L g4863 ( 
.A(n_4301),
.B(n_3448),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4299),
.Y(n_4864)
);

AOI21x1_ASAP7_75t_L g4865 ( 
.A1(n_3999),
.A2(n_3630),
.B(n_3870),
.Y(n_4865)
);

INVx2_ASAP7_75t_L g4866 ( 
.A(n_4443),
.Y(n_4866)
);

OA21x2_ASAP7_75t_L g4867 ( 
.A1(n_4162),
.A2(n_3896),
.B(n_3886),
.Y(n_4867)
);

AND2x4_ASAP7_75t_L g4868 ( 
.A(n_4186),
.B(n_3678),
.Y(n_4868)
);

AO21x1_ASAP7_75t_L g4869 ( 
.A1(n_4338),
.A2(n_3822),
.B(n_3820),
.Y(n_4869)
);

NAND2xp5_ASAP7_75t_L g4870 ( 
.A(n_4320),
.B(n_3900),
.Y(n_4870)
);

HB1xp67_ASAP7_75t_L g4871 ( 
.A(n_4258),
.Y(n_4871)
);

NAND2x1p5_ASAP7_75t_L g4872 ( 
.A(n_4301),
.B(n_3576),
.Y(n_4872)
);

AND2x2_ASAP7_75t_L g4873 ( 
.A(n_4004),
.B(n_4025),
.Y(n_4873)
);

INVx3_ASAP7_75t_L g4874 ( 
.A(n_4443),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4299),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4316),
.Y(n_4876)
);

OAI21xp5_ASAP7_75t_L g4877 ( 
.A1(n_4049),
.A2(n_3822),
.B(n_3820),
.Y(n_4877)
);

INVx2_ASAP7_75t_SL g4878 ( 
.A(n_4308),
.Y(n_4878)
);

INVx2_ASAP7_75t_L g4879 ( 
.A(n_4098),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_L g4880 ( 
.A(n_4320),
.B(n_3904),
.Y(n_4880)
);

NOR2xp33_ASAP7_75t_L g4881 ( 
.A(n_4072),
.B(n_3717),
.Y(n_4881)
);

OA21x2_ASAP7_75t_L g4882 ( 
.A1(n_4163),
.A2(n_3896),
.B(n_3886),
.Y(n_4882)
);

OAI21x1_ASAP7_75t_L g4883 ( 
.A1(n_4343),
.A2(n_3577),
.B(n_3513),
.Y(n_4883)
);

BUFx3_ASAP7_75t_L g4884 ( 
.A(n_4365),
.Y(n_4884)
);

AND2x2_ASAP7_75t_L g4885 ( 
.A(n_4025),
.B(n_3494),
.Y(n_4885)
);

OAI21x1_ASAP7_75t_L g4886 ( 
.A1(n_4351),
.A2(n_3653),
.B(n_3577),
.Y(n_4886)
);

AO31x2_ASAP7_75t_L g4887 ( 
.A1(n_4285),
.A2(n_4084),
.A3(n_4303),
.B(n_4222),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4316),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_L g4889 ( 
.A(n_4417),
.B(n_3904),
.Y(n_4889)
);

AOI21xp5_ASAP7_75t_L g4890 ( 
.A1(n_4300),
.A2(n_3923),
.B(n_3911),
.Y(n_4890)
);

AO21x1_ASAP7_75t_L g4891 ( 
.A1(n_4437),
.A2(n_3865),
.B(n_3837),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4330),
.Y(n_4892)
);

OAI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4095),
.A2(n_3865),
.B(n_3837),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4330),
.Y(n_4894)
);

INVxp67_ASAP7_75t_L g4895 ( 
.A(n_4107),
.Y(n_4895)
);

OA21x2_ASAP7_75t_L g4896 ( 
.A1(n_4407),
.A2(n_3896),
.B(n_3886),
.Y(n_4896)
);

AND2x2_ASAP7_75t_L g4897 ( 
.A(n_4504),
.B(n_3494),
.Y(n_4897)
);

INVx1_ASAP7_75t_SL g4898 ( 
.A(n_4448),
.Y(n_4898)
);

A2O1A1Ixp33_ASAP7_75t_L g4899 ( 
.A1(n_4005),
.A2(n_3631),
.B(n_3751),
.C(n_3691),
.Y(n_4899)
);

OAI21xp5_ASAP7_75t_L g4900 ( 
.A1(n_4152),
.A2(n_3869),
.B(n_3911),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4334),
.Y(n_4901)
);

AOI22xp5_ASAP7_75t_L g4902 ( 
.A1(n_3998),
.A2(n_3680),
.B1(n_3815),
.B2(n_3975),
.Y(n_4902)
);

NAND2xp5_ASAP7_75t_L g4903 ( 
.A(n_4059),
.B(n_3923),
.Y(n_4903)
);

AND2x4_ASAP7_75t_L g4904 ( 
.A(n_4186),
.B(n_3678),
.Y(n_4904)
);

BUFx2_ASAP7_75t_R g4905 ( 
.A(n_4012),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4334),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_L g4907 ( 
.A(n_4110),
.B(n_3937),
.Y(n_4907)
);

AOI21xp5_ASAP7_75t_L g4908 ( 
.A1(n_4487),
.A2(n_4498),
.B(n_4144),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4106),
.B(n_3937),
.Y(n_4909)
);

OAI21x1_ASAP7_75t_L g4910 ( 
.A1(n_4129),
.A2(n_4134),
.B(n_4382),
.Y(n_4910)
);

HB1xp67_ASAP7_75t_L g4911 ( 
.A(n_4287),
.Y(n_4911)
);

HB1xp67_ASAP7_75t_L g4912 ( 
.A(n_4287),
.Y(n_4912)
);

INVx3_ASAP7_75t_L g4913 ( 
.A(n_4389),
.Y(n_4913)
);

AND2x2_ASAP7_75t_L g4914 ( 
.A(n_4504),
.B(n_4518),
.Y(n_4914)
);

AO21x2_ASAP7_75t_L g4915 ( 
.A1(n_4312),
.A2(n_3976),
.B(n_3910),
.Y(n_4915)
);

AOI21xp5_ASAP7_75t_L g4916 ( 
.A1(n_4144),
.A2(n_3943),
.B(n_3939),
.Y(n_4916)
);

NAND2x1p5_ASAP7_75t_L g4917 ( 
.A(n_4301),
.B(n_3576),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4352),
.Y(n_4918)
);

AOI21xp5_ASAP7_75t_L g4919 ( 
.A1(n_4267),
.A2(n_3943),
.B(n_3939),
.Y(n_4919)
);

AO21x2_ASAP7_75t_L g4920 ( 
.A1(n_4348),
.A2(n_3976),
.B(n_3910),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_L g4921 ( 
.A(n_4106),
.B(n_3950),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4352),
.Y(n_4922)
);

NAND3xp33_ASAP7_75t_L g4923 ( 
.A(n_4002),
.B(n_3869),
.C(n_3950),
.Y(n_4923)
);

INVx2_ASAP7_75t_L g4924 ( 
.A(n_4098),
.Y(n_4924)
);

NOR2xp33_ASAP7_75t_L g4925 ( 
.A(n_4087),
.B(n_3853),
.Y(n_4925)
);

BUFx2_ASAP7_75t_R g4926 ( 
.A(n_4021),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4360),
.Y(n_4927)
);

AO31x2_ASAP7_75t_L g4928 ( 
.A1(n_4221),
.A2(n_3948),
.A3(n_3862),
.B(n_3871),
.Y(n_4928)
);

AND2x4_ASAP7_75t_L g4929 ( 
.A(n_4186),
.B(n_3678),
.Y(n_4929)
);

AND2x4_ASAP7_75t_L g4930 ( 
.A(n_4315),
.B(n_3691),
.Y(n_4930)
);

OR2x2_ASAP7_75t_L g4931 ( 
.A(n_4356),
.B(n_3959),
.Y(n_4931)
);

BUFx3_ASAP7_75t_L g4932 ( 
.A(n_4365),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4360),
.Y(n_4933)
);

OA21x2_ASAP7_75t_L g4934 ( 
.A1(n_4391),
.A2(n_3976),
.B(n_3910),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4371),
.Y(n_4935)
);

INVx2_ASAP7_75t_L g4936 ( 
.A(n_4098),
.Y(n_4936)
);

NAND2x1p5_ASAP7_75t_L g4937 ( 
.A(n_4301),
.B(n_3646),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4371),
.Y(n_4938)
);

OR2x2_ASAP7_75t_L g4939 ( 
.A(n_4390),
.B(n_3959),
.Y(n_4939)
);

INVx2_ASAP7_75t_L g4940 ( 
.A(n_4098),
.Y(n_4940)
);

NAND2x1p5_ASAP7_75t_L g4941 ( 
.A(n_4301),
.B(n_3646),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4374),
.Y(n_4942)
);

OAI21x1_ASAP7_75t_L g4943 ( 
.A1(n_4159),
.A2(n_4192),
.B(n_4261),
.Y(n_4943)
);

AOI22xp5_ASAP7_75t_L g4944 ( 
.A1(n_4005),
.A2(n_3680),
.B1(n_3815),
.B2(n_3975),
.Y(n_4944)
);

INVx1_ASAP7_75t_SL g4945 ( 
.A(n_4529),
.Y(n_4945)
);

CKINVDCx5p33_ASAP7_75t_R g4946 ( 
.A(n_4051),
.Y(n_4946)
);

INVx2_ASAP7_75t_L g4947 ( 
.A(n_4098),
.Y(n_4947)
);

OAI21x1_ASAP7_75t_L g4948 ( 
.A1(n_4261),
.A2(n_3669),
.B(n_3658),
.Y(n_4948)
);

AOI21xp5_ASAP7_75t_L g4949 ( 
.A1(n_4224),
.A2(n_3962),
.B(n_3961),
.Y(n_4949)
);

AO21x2_ASAP7_75t_L g4950 ( 
.A1(n_4501),
.A2(n_3988),
.B(n_3962),
.Y(n_4950)
);

AOI21xp5_ASAP7_75t_L g4951 ( 
.A1(n_4489),
.A2(n_3966),
.B(n_3961),
.Y(n_4951)
);

AO21x2_ASAP7_75t_L g4952 ( 
.A1(n_4414),
.A2(n_3988),
.B(n_3969),
.Y(n_4952)
);

NAND2x1p5_ASAP7_75t_L g4953 ( 
.A(n_4301),
.B(n_3646),
.Y(n_4953)
);

NAND2x1p5_ASAP7_75t_L g4954 ( 
.A(n_4516),
.B(n_3646),
.Y(n_4954)
);

OAI21xp5_ASAP7_75t_L g4955 ( 
.A1(n_4191),
.A2(n_3966),
.B(n_3862),
.Y(n_4955)
);

INVx2_ASAP7_75t_L g4956 ( 
.A(n_4120),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4473),
.B(n_4569),
.Y(n_4957)
);

INVx2_ASAP7_75t_SL g4958 ( 
.A(n_4308),
.Y(n_4958)
);

AO21x2_ASAP7_75t_L g4959 ( 
.A1(n_4450),
.A2(n_2400),
.B(n_2360),
.Y(n_4959)
);

OR2x6_ASAP7_75t_L g4960 ( 
.A(n_4247),
.B(n_3691),
.Y(n_4960)
);

OR2x6_ASAP7_75t_L g4961 ( 
.A(n_4037),
.B(n_3691),
.Y(n_4961)
);

AO31x2_ASAP7_75t_L g4962 ( 
.A1(n_4305),
.A2(n_3994),
.A3(n_3968),
.B(n_3957),
.Y(n_4962)
);

INVx2_ASAP7_75t_L g4963 ( 
.A(n_4120),
.Y(n_4963)
);

AOI21xp5_ASAP7_75t_L g4964 ( 
.A1(n_4477),
.A2(n_4376),
.B(n_4478),
.Y(n_4964)
);

CKINVDCx5p33_ASAP7_75t_R g4965 ( 
.A(n_4052),
.Y(n_4965)
);

OAI21x1_ASAP7_75t_SL g4966 ( 
.A1(n_4421),
.A2(n_3871),
.B(n_3859),
.Y(n_4966)
);

OAI21x1_ASAP7_75t_L g4967 ( 
.A1(n_4037),
.A2(n_3703),
.B(n_3674),
.Y(n_4967)
);

OAI21x1_ASAP7_75t_L g4968 ( 
.A1(n_4037),
.A2(n_3703),
.B(n_3674),
.Y(n_4968)
);

OA21x2_ASAP7_75t_L g4969 ( 
.A1(n_4486),
.A2(n_3888),
.B(n_3884),
.Y(n_4969)
);

OAI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4150),
.A2(n_3888),
.B(n_3884),
.Y(n_4970)
);

OAI21x1_ASAP7_75t_L g4971 ( 
.A1(n_4055),
.A2(n_3704),
.B(n_3703),
.Y(n_4971)
);

OAI21xp5_ASAP7_75t_L g4972 ( 
.A1(n_4439),
.A2(n_3922),
.B(n_3920),
.Y(n_4972)
);

HB1xp67_ASAP7_75t_L g4973 ( 
.A(n_4329),
.Y(n_4973)
);

OR2x2_ASAP7_75t_L g4974 ( 
.A(n_4390),
.B(n_3825),
.Y(n_4974)
);

AND2x4_ASAP7_75t_L g4975 ( 
.A(n_4315),
.B(n_3737),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4374),
.Y(n_4976)
);

NAND2x1p5_ASAP7_75t_L g4977 ( 
.A(n_4516),
.B(n_3819),
.Y(n_4977)
);

INVx1_ASAP7_75t_L g4978 ( 
.A(n_4388),
.Y(n_4978)
);

OA21x2_ASAP7_75t_L g4979 ( 
.A1(n_4298),
.A2(n_3934),
.B(n_3920),
.Y(n_4979)
);

CKINVDCx5p33_ASAP7_75t_R g4980 ( 
.A(n_4559),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_L g4981 ( 
.A(n_4569),
.B(n_3934),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4388),
.Y(n_4982)
);

OAI21x1_ASAP7_75t_L g4983 ( 
.A1(n_4055),
.A2(n_4467),
.B(n_4436),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_L g4984 ( 
.A(n_4447),
.B(n_3947),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4413),
.Y(n_4985)
);

OA21x2_ASAP7_75t_L g4986 ( 
.A1(n_4441),
.A2(n_3948),
.B(n_3947),
.Y(n_4986)
);

NAND2x1p5_ASAP7_75t_L g4987 ( 
.A(n_4516),
.B(n_4421),
.Y(n_4987)
);

AOI21x1_ASAP7_75t_L g4988 ( 
.A1(n_4132),
.A2(n_3630),
.B(n_3619),
.Y(n_4988)
);

OA21x2_ASAP7_75t_L g4989 ( 
.A1(n_4542),
.A2(n_3949),
.B(n_3957),
.Y(n_4989)
);

INVx1_ASAP7_75t_L g4990 ( 
.A(n_4413),
.Y(n_4990)
);

OA21x2_ASAP7_75t_L g4991 ( 
.A1(n_4239),
.A2(n_3949),
.B(n_3751),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_L g4992 ( 
.A(n_4447),
.B(n_3825),
.Y(n_4992)
);

OR2x2_ASAP7_75t_L g4993 ( 
.A(n_4336),
.B(n_3825),
.Y(n_4993)
);

AOI22x1_ASAP7_75t_L g4994 ( 
.A1(n_4479),
.A2(n_3903),
.B1(n_3887),
.B2(n_3538),
.Y(n_4994)
);

OR2x6_ASAP7_75t_L g4995 ( 
.A(n_4402),
.B(n_3737),
.Y(n_4995)
);

CKINVDCx5p33_ASAP7_75t_R g4996 ( 
.A(n_4465),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4283),
.B(n_4288),
.Y(n_4997)
);

AOI22xp33_ASAP7_75t_L g4998 ( 
.A1(n_4050),
.A2(n_3680),
.B1(n_3975),
.B2(n_3815),
.Y(n_4998)
);

INVx2_ASAP7_75t_L g4999 ( 
.A(n_4120),
.Y(n_4999)
);

OR2x6_ASAP7_75t_L g5000 ( 
.A(n_4402),
.B(n_3737),
.Y(n_5000)
);

BUFx3_ASAP7_75t_L g5001 ( 
.A(n_4365),
.Y(n_5001)
);

INVx3_ASAP7_75t_L g5002 ( 
.A(n_4389),
.Y(n_5002)
);

INVx3_ASAP7_75t_L g5003 ( 
.A(n_4389),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4418),
.B(n_3825),
.Y(n_5004)
);

INVx4_ASAP7_75t_L g5005 ( 
.A(n_4555),
.Y(n_5005)
);

AOI21xp33_ASAP7_75t_SL g5006 ( 
.A1(n_4397),
.A2(n_3951),
.B(n_3749),
.Y(n_5006)
);

OR2x2_ASAP7_75t_L g5007 ( 
.A(n_4336),
.B(n_3825),
.Y(n_5007)
);

OR2x6_ASAP7_75t_L g5008 ( 
.A(n_4402),
.B(n_3737),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4418),
.B(n_4419),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4419),
.Y(n_5010)
);

BUFx2_ASAP7_75t_R g5011 ( 
.A(n_4021),
.Y(n_5011)
);

NOR2xp33_ASAP7_75t_L g5012 ( 
.A(n_4175),
.B(n_3538),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4424),
.Y(n_5013)
);

OAI21x1_ASAP7_75t_L g5014 ( 
.A1(n_4463),
.A2(n_3726),
.B(n_3844),
.Y(n_5014)
);

OAI21x1_ASAP7_75t_L g5015 ( 
.A1(n_4494),
.A2(n_3726),
.B(n_3844),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_SL g5016 ( 
.A(n_4365),
.B(n_3538),
.Y(n_5016)
);

AO21x2_ASAP7_75t_L g5017 ( 
.A1(n_4461),
.A2(n_2535),
.B(n_2400),
.Y(n_5017)
);

OA21x2_ASAP7_75t_L g5018 ( 
.A1(n_4249),
.A2(n_3751),
.B(n_2402),
.Y(n_5018)
);

BUFx3_ASAP7_75t_L g5019 ( 
.A(n_4365),
.Y(n_5019)
);

NAND2xp5_ASAP7_75t_L g5020 ( 
.A(n_4424),
.B(n_3825),
.Y(n_5020)
);

AND2x4_ASAP7_75t_L g5021 ( 
.A(n_4315),
.B(n_4367),
.Y(n_5021)
);

OAI21x1_ASAP7_75t_L g5022 ( 
.A1(n_4398),
.A2(n_3766),
.B(n_3741),
.Y(n_5022)
);

INVxp67_ASAP7_75t_SL g5023 ( 
.A(n_4132),
.Y(n_5023)
);

NOR2xp33_ASAP7_75t_SL g5024 ( 
.A(n_4516),
.B(n_3819),
.Y(n_5024)
);

OAI21xp5_ASAP7_75t_L g5025 ( 
.A1(n_4195),
.A2(n_3619),
.B(n_3895),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4433),
.Y(n_5026)
);

NAND2xp5_ASAP7_75t_L g5027 ( 
.A(n_4433),
.B(n_4452),
.Y(n_5027)
);

INVx2_ASAP7_75t_L g5028 ( 
.A(n_4120),
.Y(n_5028)
);

HB1xp67_ASAP7_75t_L g5029 ( 
.A(n_4329),
.Y(n_5029)
);

BUFx8_ASAP7_75t_L g5030 ( 
.A(n_4188),
.Y(n_5030)
);

INVx3_ASAP7_75t_SL g5031 ( 
.A(n_4118),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_4452),
.B(n_3841),
.Y(n_5032)
);

AO21x2_ASAP7_75t_L g5033 ( 
.A1(n_4216),
.A2(n_2531),
.B(n_2402),
.Y(n_5033)
);

OAI21xp5_ASAP7_75t_L g5034 ( 
.A1(n_4271),
.A2(n_3895),
.B(n_3899),
.Y(n_5034)
);

AND2x4_ASAP7_75t_L g5035 ( 
.A(n_4367),
.B(n_3751),
.Y(n_5035)
);

INVx3_ASAP7_75t_L g5036 ( 
.A(n_4389),
.Y(n_5036)
);

INVx2_ASAP7_75t_L g5037 ( 
.A(n_4120),
.Y(n_5037)
);

OA21x2_ASAP7_75t_L g5038 ( 
.A1(n_4339),
.A2(n_2531),
.B(n_2407),
.Y(n_5038)
);

OAI21x1_ASAP7_75t_L g5039 ( 
.A1(n_4220),
.A2(n_4233),
.B(n_4077),
.Y(n_5039)
);

AOI21xp5_ASAP7_75t_L g5040 ( 
.A1(n_4515),
.A2(n_3895),
.B(n_3899),
.Y(n_5040)
);

BUFx6f_ASAP7_75t_L g5041 ( 
.A(n_4516),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_4466),
.B(n_4483),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_4466),
.Y(n_5043)
);

OA21x2_ASAP7_75t_L g5044 ( 
.A1(n_4340),
.A2(n_2525),
.B(n_2407),
.Y(n_5044)
);

INVx4_ASAP7_75t_L g5045 ( 
.A(n_4145),
.Y(n_5045)
);

INVx2_ASAP7_75t_L g5046 ( 
.A(n_4547),
.Y(n_5046)
);

HB1xp67_ASAP7_75t_L g5047 ( 
.A(n_4132),
.Y(n_5047)
);

HB1xp67_ASAP7_75t_L g5048 ( 
.A(n_4483),
.Y(n_5048)
);

INVx8_ASAP7_75t_L g5049 ( 
.A(n_4425),
.Y(n_5049)
);

CKINVDCx6p67_ASAP7_75t_R g5050 ( 
.A(n_4118),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4495),
.Y(n_5051)
);

OAI21x1_ASAP7_75t_L g5052 ( 
.A1(n_4387),
.A2(n_3970),
.B(n_3844),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4495),
.Y(n_5053)
);

INVx2_ASAP7_75t_L g5054 ( 
.A(n_4547),
.Y(n_5054)
);

HB1xp67_ASAP7_75t_L g5055 ( 
.A(n_4506),
.Y(n_5055)
);

INVx5_ASAP7_75t_L g5056 ( 
.A(n_4516),
.Y(n_5056)
);

INVx2_ASAP7_75t_L g5057 ( 
.A(n_4547),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4506),
.Y(n_5058)
);

AOI21xp5_ASAP7_75t_L g5059 ( 
.A1(n_4525),
.A2(n_3899),
.B(n_3970),
.Y(n_5059)
);

INVx2_ASAP7_75t_SL g5060 ( 
.A(n_4308),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4519),
.Y(n_5061)
);

NAND2x1p5_ASAP7_75t_L g5062 ( 
.A(n_4514),
.B(n_3819),
.Y(n_5062)
);

OAI21xp5_ASAP7_75t_L g5063 ( 
.A1(n_4271),
.A2(n_3975),
.B(n_3815),
.Y(n_5063)
);

NAND2x1p5_ASAP7_75t_L g5064 ( 
.A(n_4514),
.B(n_4426),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4519),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_4547),
.Y(n_5066)
);

CKINVDCx14_ASAP7_75t_R g5067 ( 
.A(n_4521),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_4539),
.Y(n_5068)
);

INVx2_ASAP7_75t_L g5069 ( 
.A(n_4547),
.Y(n_5069)
);

OAI21x1_ASAP7_75t_SL g5070 ( 
.A1(n_4401),
.A2(n_3942),
.B(n_3860),
.Y(n_5070)
);

BUFx12f_ASAP7_75t_L g5071 ( 
.A(n_4041),
.Y(n_5071)
);

BUFx6f_ASAP7_75t_L g5072 ( 
.A(n_4038),
.Y(n_5072)
);

NAND2xp5_ASAP7_75t_L g5073 ( 
.A(n_4539),
.B(n_3841),
.Y(n_5073)
);

CKINVDCx11_ASAP7_75t_R g5074 ( 
.A(n_4213),
.Y(n_5074)
);

BUFx12f_ASAP7_75t_L g5075 ( 
.A(n_4041),
.Y(n_5075)
);

AOI21x1_ASAP7_75t_L g5076 ( 
.A1(n_4426),
.A2(n_2517),
.B(n_2414),
.Y(n_5076)
);

INVx2_ASAP7_75t_L g5077 ( 
.A(n_4036),
.Y(n_5077)
);

OAI21xp5_ASAP7_75t_L g5078 ( 
.A1(n_4295),
.A2(n_3815),
.B(n_3975),
.Y(n_5078)
);

INVx2_ASAP7_75t_SL g5079 ( 
.A(n_4562),
.Y(n_5079)
);

INVx2_ASAP7_75t_L g5080 ( 
.A(n_4036),
.Y(n_5080)
);

HB1xp67_ASAP7_75t_L g5081 ( 
.A(n_4587),
.Y(n_5081)
);

BUFx3_ASAP7_75t_L g5082 ( 
.A(n_4585),
.Y(n_5082)
);

AOI21xp5_ASAP7_75t_L g5083 ( 
.A1(n_4810),
.A2(n_4003),
.B(n_4079),
.Y(n_5083)
);

AO21x2_ASAP7_75t_L g5084 ( 
.A1(n_4606),
.A2(n_4022),
.B(n_4015),
.Y(n_5084)
);

OR2x2_ASAP7_75t_L g5085 ( 
.A(n_4660),
.B(n_4263),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_L g5086 ( 
.A(n_4794),
.B(n_4265),
.Y(n_5086)
);

NAND2xp5_ASAP7_75t_L g5087 ( 
.A(n_4794),
.B(n_4290),
.Y(n_5087)
);

INVx2_ASAP7_75t_L g5088 ( 
.A(n_4854),
.Y(n_5088)
);

AND2x4_ASAP7_75t_L g5089 ( 
.A(n_4600),
.B(n_4363),
.Y(n_5089)
);

NOR2xp33_ASAP7_75t_L g5090 ( 
.A(n_4585),
.B(n_4103),
.Y(n_5090)
);

AOI21xp5_ASAP7_75t_L g5091 ( 
.A1(n_4810),
.A2(n_4723),
.B(n_4596),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_4614),
.B(n_4223),
.Y(n_5092)
);

OAI221xp5_ASAP7_75t_L g5093 ( 
.A1(n_4723),
.A2(n_4353),
.B1(n_4415),
.B2(n_4151),
.C(n_4174),
.Y(n_5093)
);

AOI222xp33_ASAP7_75t_L g5094 ( 
.A1(n_4596),
.A2(n_4523),
.B1(n_4094),
.B2(n_4164),
.C1(n_4349),
.C2(n_4104),
.Y(n_5094)
);

AO21x2_ASAP7_75t_L g5095 ( 
.A1(n_4606),
.A2(n_4061),
.B(n_4042),
.Y(n_5095)
);

OA21x2_ASAP7_75t_L g5096 ( 
.A1(n_4680),
.A2(n_4061),
.B(n_4042),
.Y(n_5096)
);

AND2x2_ASAP7_75t_L g5097 ( 
.A(n_4703),
.B(n_4529),
.Y(n_5097)
);

BUFx2_ASAP7_75t_L g5098 ( 
.A(n_4741),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4595),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_4595),
.Y(n_5100)
);

AOI21xp5_ASAP7_75t_L g5101 ( 
.A1(n_4601),
.A2(n_4456),
.B(n_4427),
.Y(n_5101)
);

BUFx2_ASAP7_75t_L g5102 ( 
.A(n_4741),
.Y(n_5102)
);

NAND2xp5_ASAP7_75t_L g5103 ( 
.A(n_4614),
.B(n_4232),
.Y(n_5103)
);

AOI21xp5_ASAP7_75t_L g5104 ( 
.A1(n_4601),
.A2(n_4321),
.B(n_4062),
.Y(n_5104)
);

BUFx10_ASAP7_75t_L g5105 ( 
.A(n_4624),
.Y(n_5105)
);

NAND2xp5_ASAP7_75t_L g5106 ( 
.A(n_4644),
.B(n_4675),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_4633),
.Y(n_5107)
);

NAND2xp5_ASAP7_75t_SL g5108 ( 
.A(n_4641),
.B(n_4365),
.Y(n_5108)
);

OAI21x1_ASAP7_75t_L g5109 ( 
.A1(n_4680),
.A2(n_4440),
.B(n_4409),
.Y(n_5109)
);

OAI21xp5_ASAP7_75t_L g5110 ( 
.A1(n_4816),
.A2(n_4350),
.B(n_4295),
.Y(n_5110)
);

AND2x4_ASAP7_75t_L g5111 ( 
.A(n_4600),
.B(n_4363),
.Y(n_5111)
);

INVx2_ASAP7_75t_L g5112 ( 
.A(n_4854),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4633),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_4644),
.B(n_4133),
.Y(n_5114)
);

NAND2xp5_ASAP7_75t_L g5115 ( 
.A(n_4675),
.B(n_4149),
.Y(n_5115)
);

INVx2_ASAP7_75t_L g5116 ( 
.A(n_4854),
.Y(n_5116)
);

OAI21x1_ASAP7_75t_L g5117 ( 
.A1(n_4662),
.A2(n_4440),
.B(n_4409),
.Y(n_5117)
);

OA21x2_ASAP7_75t_L g5118 ( 
.A1(n_4635),
.A2(n_4099),
.B(n_4089),
.Y(n_5118)
);

AOI21xp5_ASAP7_75t_L g5119 ( 
.A1(n_4964),
.A2(n_4137),
.B(n_4333),
.Y(n_5119)
);

INVx2_ASAP7_75t_L g5120 ( 
.A(n_4854),
.Y(n_5120)
);

OAI221xp5_ASAP7_75t_L g5121 ( 
.A1(n_4816),
.A2(n_4086),
.B1(n_4332),
.B2(n_4350),
.C(n_4422),
.Y(n_5121)
);

NAND2xp5_ASAP7_75t_L g5122 ( 
.A(n_4679),
.B(n_4092),
.Y(n_5122)
);

AO21x2_ASAP7_75t_L g5123 ( 
.A1(n_4606),
.A2(n_4099),
.B(n_4089),
.Y(n_5123)
);

NAND2xp5_ASAP7_75t_L g5124 ( 
.A(n_4679),
.B(n_4108),
.Y(n_5124)
);

CKINVDCx5p33_ASAP7_75t_R g5125 ( 
.A(n_4627),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_L g5126 ( 
.A(n_4667),
.B(n_4111),
.Y(n_5126)
);

OAI21xp5_ASAP7_75t_L g5127 ( 
.A1(n_4590),
.A2(n_4449),
.B(n_4269),
.Y(n_5127)
);

AOI22xp33_ASAP7_75t_L g5128 ( 
.A1(n_4593),
.A2(n_4010),
.B1(n_4123),
.B2(n_4090),
.Y(n_5128)
);

NOR2xp67_ASAP7_75t_SL g5129 ( 
.A(n_5071),
.B(n_4093),
.Y(n_5129)
);

AOI21x1_ASAP7_75t_L g5130 ( 
.A1(n_4615),
.A2(n_4126),
.B(n_4124),
.Y(n_5130)
);

OAI22xp5_ASAP7_75t_SL g5131 ( 
.A1(n_5067),
.A2(n_4484),
.B1(n_4397),
.B2(n_4093),
.Y(n_5131)
);

AOI21xp5_ASAP7_75t_L g5132 ( 
.A1(n_4964),
.A2(n_4184),
.B(n_4471),
.Y(n_5132)
);

HB1xp67_ASAP7_75t_L g5133 ( 
.A(n_4587),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_5048),
.Y(n_5134)
);

BUFx3_ASAP7_75t_L g5135 ( 
.A(n_4585),
.Y(n_5135)
);

AOI21xp5_ASAP7_75t_L g5136 ( 
.A1(n_4735),
.A2(n_4184),
.B(n_4472),
.Y(n_5136)
);

OR2x6_ASAP7_75t_L g5137 ( 
.A(n_4594),
.B(n_4402),
.Y(n_5137)
);

AO31x2_ASAP7_75t_L g5138 ( 
.A1(n_4641),
.A2(n_4244),
.A3(n_4257),
.B(n_4394),
.Y(n_5138)
);

OAI21xp5_ASAP7_75t_L g5139 ( 
.A1(n_4590),
.A2(n_4166),
.B(n_4058),
.Y(n_5139)
);

OA21x2_ASAP7_75t_L g5140 ( 
.A1(n_4635),
.A2(n_4126),
.B(n_4124),
.Y(n_5140)
);

INVx2_ASAP7_75t_L g5141 ( 
.A(n_4854),
.Y(n_5141)
);

AOI21x1_ASAP7_75t_L g5142 ( 
.A1(n_4615),
.A2(n_4142),
.B(n_4130),
.Y(n_5142)
);

AND2x4_ASAP7_75t_L g5143 ( 
.A(n_4600),
.B(n_4363),
.Y(n_5143)
);

OAI21x1_ASAP7_75t_L g5144 ( 
.A1(n_4662),
.A2(n_4440),
.B(n_4409),
.Y(n_5144)
);

INVx2_ASAP7_75t_SL g5145 ( 
.A(n_4624),
.Y(n_5145)
);

HB1xp67_ASAP7_75t_L g5146 ( 
.A(n_4592),
.Y(n_5146)
);

OAI21xp5_ASAP7_75t_L g5147 ( 
.A1(n_4796),
.A2(n_4166),
.B(n_4058),
.Y(n_5147)
);

OA21x2_ASAP7_75t_L g5148 ( 
.A1(n_4709),
.A2(n_4142),
.B(n_4130),
.Y(n_5148)
);

HB1xp67_ASAP7_75t_L g5149 ( 
.A(n_4592),
.Y(n_5149)
);

NAND2xp5_ASAP7_75t_L g5150 ( 
.A(n_4667),
.B(n_4115),
.Y(n_5150)
);

NAND3xp33_ASAP7_75t_L g5151 ( 
.A(n_4628),
.B(n_4259),
.C(n_4242),
.Y(n_5151)
);

AOI22xp33_ASAP7_75t_L g5152 ( 
.A1(n_4593),
.A2(n_4090),
.B1(n_4123),
.B2(n_4386),
.Y(n_5152)
);

AOI322xp5_ASAP7_75t_L g5153 ( 
.A1(n_4593),
.A2(n_4160),
.A3(n_4009),
.B1(n_4332),
.B2(n_4254),
.C1(n_4341),
.C2(n_4143),
.Y(n_5153)
);

INVx3_ASAP7_75t_L g5154 ( 
.A(n_4672),
.Y(n_5154)
);

INVx2_ASAP7_75t_L g5155 ( 
.A(n_4854),
.Y(n_5155)
);

A2O1A1Ixp33_ASAP7_75t_L g5156 ( 
.A1(n_4783),
.A2(n_4190),
.B(n_4189),
.C(n_4193),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_L g5157 ( 
.A(n_4683),
.B(n_4155),
.Y(n_5157)
);

BUFx8_ASAP7_75t_L g5158 ( 
.A(n_4585),
.Y(n_5158)
);

OR2x2_ASAP7_75t_L g5159 ( 
.A(n_4660),
.B(n_4263),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_5048),
.Y(n_5160)
);

AOI22xp33_ASAP7_75t_L g5161 ( 
.A1(n_4783),
.A2(n_4523),
.B1(n_4365),
.B2(n_4358),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_4636),
.Y(n_5162)
);

OA21x2_ASAP7_75t_L g5163 ( 
.A1(n_4709),
.A2(n_4185),
.B(n_4158),
.Y(n_5163)
);

AOI21xp5_ASAP7_75t_L g5164 ( 
.A1(n_4735),
.A2(n_4548),
.B(n_4362),
.Y(n_5164)
);

INVx2_ASAP7_75t_L g5165 ( 
.A(n_4879),
.Y(n_5165)
);

INVx2_ASAP7_75t_L g5166 ( 
.A(n_4879),
.Y(n_5166)
);

AND2x2_ASAP7_75t_L g5167 ( 
.A(n_4703),
.B(n_4518),
.Y(n_5167)
);

HB1xp67_ASAP7_75t_L g5168 ( 
.A(n_4630),
.Y(n_5168)
);

OAI21x1_ASAP7_75t_L g5169 ( 
.A1(n_4662),
.A2(n_4540),
.B(n_4185),
.Y(n_5169)
);

OR2x2_ASAP7_75t_L g5170 ( 
.A(n_4660),
.B(n_4161),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_4636),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_4647),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_5055),
.Y(n_5173)
);

OA21x2_ASAP7_75t_L g5174 ( 
.A1(n_4713),
.A2(n_4196),
.B(n_4158),
.Y(n_5174)
);

AOI22xp33_ASAP7_75t_L g5175 ( 
.A1(n_4783),
.A2(n_4523),
.B1(n_3680),
.B2(n_4383),
.Y(n_5175)
);

AOI21xp5_ASAP7_75t_L g5176 ( 
.A1(n_4796),
.A2(n_4346),
.B(n_4566),
.Y(n_5176)
);

INVx2_ASAP7_75t_L g5177 ( 
.A(n_4879),
.Y(n_5177)
);

INVx2_ASAP7_75t_L g5178 ( 
.A(n_4879),
.Y(n_5178)
);

AND2x4_ASAP7_75t_L g5179 ( 
.A(n_4600),
.B(n_4363),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_L g5180 ( 
.A(n_4683),
.B(n_4161),
.Y(n_5180)
);

INVxp67_ASAP7_75t_L g5181 ( 
.A(n_4793),
.Y(n_5181)
);

AO21x2_ASAP7_75t_L g5182 ( 
.A1(n_4713),
.A2(n_4235),
.B(n_4196),
.Y(n_5182)
);

NAND2xp5_ASAP7_75t_L g5183 ( 
.A(n_4710),
.B(n_4203),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_L g5184 ( 
.A(n_4710),
.B(n_4203),
.Y(n_5184)
);

AND2x2_ASAP7_75t_L g5185 ( 
.A(n_4703),
.B(n_4738),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_4647),
.Y(n_5186)
);

INVx3_ASAP7_75t_L g5187 ( 
.A(n_4672),
.Y(n_5187)
);

A2O1A1Ixp33_ASAP7_75t_L g5188 ( 
.A1(n_4784),
.A2(n_4383),
.B(n_4502),
.C(n_4434),
.Y(n_5188)
);

OAI22xp5_ASAP7_75t_L g5189 ( 
.A1(n_4579),
.A2(n_4784),
.B1(n_4802),
.B2(n_4759),
.Y(n_5189)
);

OR2x2_ASAP7_75t_L g5190 ( 
.A(n_4907),
.B(n_4208),
.Y(n_5190)
);

A2O1A1Ixp33_ASAP7_75t_L g5191 ( 
.A1(n_4784),
.A2(n_4502),
.B(n_4434),
.C(n_4499),
.Y(n_5191)
);

AOI22xp5_ASAP7_75t_L g5192 ( 
.A1(n_4756),
.A2(n_4499),
.B1(n_4284),
.B2(n_4341),
.Y(n_5192)
);

AND2x2_ASAP7_75t_L g5193 ( 
.A(n_4738),
.B(n_4302),
.Y(n_5193)
);

AOI22xp33_ASAP7_75t_L g5194 ( 
.A1(n_4802),
.A2(n_4523),
.B1(n_3680),
.B2(n_4513),
.Y(n_5194)
);

AOI22xp33_ASAP7_75t_L g5195 ( 
.A1(n_4802),
.A2(n_3680),
.B1(n_4500),
.B2(n_4128),
.Y(n_5195)
);

AOI21xp5_ASAP7_75t_L g5196 ( 
.A1(n_4579),
.A2(n_4395),
.B(n_4246),
.Y(n_5196)
);

OR2x6_ASAP7_75t_L g5197 ( 
.A(n_4594),
.B(n_4204),
.Y(n_5197)
);

AOI22xp33_ASAP7_75t_L g5198 ( 
.A1(n_4969),
.A2(n_3680),
.B1(n_4128),
.B2(n_4119),
.Y(n_5198)
);

OAI21xp5_ASAP7_75t_L g5199 ( 
.A1(n_4628),
.A2(n_4242),
.B(n_4215),
.Y(n_5199)
);

AOI22xp33_ASAP7_75t_SL g5200 ( 
.A1(n_4756),
.A2(n_4581),
.B1(n_4612),
.B2(n_4586),
.Y(n_5200)
);

AO21x2_ASAP7_75t_L g5201 ( 
.A1(n_4637),
.A2(n_4241),
.B(n_4235),
.Y(n_5201)
);

AO21x2_ASAP7_75t_L g5202 ( 
.A1(n_4637),
.A2(n_4289),
.B(n_4241),
.Y(n_5202)
);

AOI22xp33_ASAP7_75t_L g5203 ( 
.A1(n_4969),
.A2(n_4128),
.B1(n_4119),
.B2(n_4218),
.Y(n_5203)
);

AOI221xp5_ASAP7_75t_L g5204 ( 
.A1(n_4756),
.A2(n_4156),
.B1(n_4178),
.B2(n_4550),
.C(n_4571),
.Y(n_5204)
);

AOI21xp5_ASAP7_75t_L g5205 ( 
.A1(n_4728),
.A2(n_4243),
.B(n_4344),
.Y(n_5205)
);

AO31x2_ASAP7_75t_L g5206 ( 
.A1(n_4641),
.A2(n_4306),
.A3(n_4317),
.B(n_4289),
.Y(n_5206)
);

AOI21xp5_ASAP7_75t_SL g5207 ( 
.A1(n_4618),
.A2(n_4103),
.B(n_4180),
.Y(n_5207)
);

HB1xp67_ASAP7_75t_L g5208 ( 
.A(n_4630),
.Y(n_5208)
);

A2O1A1Ixp33_ASAP7_75t_L g5209 ( 
.A1(n_4726),
.A2(n_4537),
.B(n_4070),
.C(n_4268),
.Y(n_5209)
);

BUFx12f_ASAP7_75t_L g5210 ( 
.A(n_4772),
.Y(n_5210)
);

AOI22xp5_ASAP7_75t_L g5211 ( 
.A1(n_4728),
.A2(n_4323),
.B1(n_4128),
.B2(n_4119),
.Y(n_5211)
);

AOI21xp5_ASAP7_75t_L g5212 ( 
.A1(n_4728),
.A2(n_4266),
.B(n_4535),
.Y(n_5212)
);

OAI21xp5_ASAP7_75t_SL g5213 ( 
.A1(n_4821),
.A2(n_4586),
.B(n_4581),
.Y(n_5213)
);

OAI321xp33_ASAP7_75t_L g5214 ( 
.A1(n_4672),
.A2(n_4727),
.A3(n_4615),
.B1(n_4726),
.B2(n_4716),
.C(n_4612),
.Y(n_5214)
);

INVx4_ASAP7_75t_SL g5215 ( 
.A(n_4624),
.Y(n_5215)
);

OAI21x1_ASAP7_75t_L g5216 ( 
.A1(n_4908),
.A2(n_4540),
.B(n_4317),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_4695),
.B(n_4215),
.Y(n_5217)
);

NOR2xp33_ASAP7_75t_SL g5218 ( 
.A(n_4665),
.B(n_4180),
.Y(n_5218)
);

CKINVDCx11_ASAP7_75t_R g5219 ( 
.A(n_4772),
.Y(n_5219)
);

OAI221xp5_ASAP7_75t_L g5220 ( 
.A1(n_4628),
.A2(n_4716),
.B1(n_4970),
.B2(n_4893),
.C(n_5034),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_4695),
.B(n_4337),
.Y(n_5221)
);

OAI221xp5_ASAP7_75t_L g5222 ( 
.A1(n_4970),
.A2(n_4893),
.B1(n_5034),
.B2(n_4786),
.C(n_4609),
.Y(n_5222)
);

AO31x2_ASAP7_75t_L g5223 ( 
.A1(n_4869),
.A2(n_4306),
.A3(n_4392),
.B(n_4354),
.Y(n_5223)
);

HB1xp67_ASAP7_75t_L g5224 ( 
.A(n_4664),
.Y(n_5224)
);

AOI222xp33_ASAP7_75t_L g5225 ( 
.A1(n_4609),
.A2(n_4561),
.B1(n_4538),
.B2(n_4543),
.C1(n_4568),
.C2(n_4006),
.Y(n_5225)
);

HB1xp67_ASAP7_75t_L g5226 ( 
.A(n_4664),
.Y(n_5226)
);

AOI21xp5_ASAP7_75t_L g5227 ( 
.A1(n_4728),
.A2(n_4119),
.B(n_4554),
.Y(n_5227)
);

OAI22xp5_ASAP7_75t_L g5228 ( 
.A1(n_4759),
.A2(n_4634),
.B1(n_4597),
.B2(n_4728),
.Y(n_5228)
);

AOI21xp5_ASAP7_75t_L g5229 ( 
.A1(n_4728),
.A2(n_4554),
.B(n_4528),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_5055),
.Y(n_5230)
);

OA21x2_ASAP7_75t_L g5231 ( 
.A1(n_4805),
.A2(n_4886),
.B(n_4883),
.Y(n_5231)
);

NAND2xp5_ASAP7_75t_L g5232 ( 
.A(n_4748),
.B(n_4432),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_4607),
.Y(n_5233)
);

NAND2xp5_ASAP7_75t_L g5234 ( 
.A(n_4748),
.B(n_4474),
.Y(n_5234)
);

CKINVDCx6p67_ASAP7_75t_R g5235 ( 
.A(n_5071),
.Y(n_5235)
);

OR2x2_ASAP7_75t_L g5236 ( 
.A(n_4907),
.B(n_4245),
.Y(n_5236)
);

INVx1_ASAP7_75t_L g5237 ( 
.A(n_4607),
.Y(n_5237)
);

BUFx12f_ASAP7_75t_L g5238 ( 
.A(n_5074),
.Y(n_5238)
);

AOI21xp5_ASAP7_75t_L g5239 ( 
.A1(n_4773),
.A2(n_4140),
.B(n_4342),
.Y(n_5239)
);

NAND3xp33_ASAP7_75t_L g5240 ( 
.A(n_4791),
.B(n_4270),
.C(n_4361),
.Y(n_5240)
);

OAI21x1_ASAP7_75t_L g5241 ( 
.A1(n_4908),
.A2(n_4540),
.B(n_4392),
.Y(n_5241)
);

OR2x2_ASAP7_75t_L g5242 ( 
.A(n_4957),
.B(n_4370),
.Y(n_5242)
);

NAND2xp5_ASAP7_75t_L g5243 ( 
.A(n_4767),
.B(n_4550),
.Y(n_5243)
);

AOI22xp33_ASAP7_75t_SL g5244 ( 
.A1(n_4581),
.A2(n_4323),
.B1(n_4006),
.B2(n_4008),
.Y(n_5244)
);

OR2x2_ASAP7_75t_L g5245 ( 
.A(n_4957),
.B(n_4372),
.Y(n_5245)
);

AO31x2_ASAP7_75t_L g5246 ( 
.A1(n_4869),
.A2(n_4396),
.A3(n_4453),
.B(n_4354),
.Y(n_5246)
);

AOI21xp5_ASAP7_75t_L g5247 ( 
.A1(n_4773),
.A2(n_4380),
.B(n_4273),
.Y(n_5247)
);

OA21x2_ASAP7_75t_L g5248 ( 
.A1(n_4805),
.A2(n_4453),
.B(n_4396),
.Y(n_5248)
);

AOI21x1_ASAP7_75t_L g5249 ( 
.A1(n_5047),
.A2(n_4460),
.B(n_4454),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_4607),
.Y(n_5250)
);

AOI21xp5_ASAP7_75t_L g5251 ( 
.A1(n_4608),
.A2(n_4281),
.B(n_4272),
.Y(n_5251)
);

INVx4_ASAP7_75t_SL g5252 ( 
.A(n_4624),
.Y(n_5252)
);

AOI21xp33_ASAP7_75t_L g5253 ( 
.A1(n_4791),
.A2(n_4310),
.B(n_4420),
.Y(n_5253)
);

OAI22xp5_ASAP7_75t_L g5254 ( 
.A1(n_4597),
.A2(n_4331),
.B1(n_4484),
.B2(n_4537),
.Y(n_5254)
);

AOI22xp33_ASAP7_75t_L g5255 ( 
.A1(n_4969),
.A2(n_3975),
.B1(n_3815),
.B2(n_4323),
.Y(n_5255)
);

AOI21xp5_ASAP7_75t_L g5256 ( 
.A1(n_4608),
.A2(n_4406),
.B(n_4399),
.Y(n_5256)
);

AND2x2_ASAP7_75t_SL g5257 ( 
.A(n_4674),
.B(n_4145),
.Y(n_5257)
);

BUFx3_ASAP7_75t_L g5258 ( 
.A(n_4627),
.Y(n_5258)
);

INVx4_ASAP7_75t_SL g5259 ( 
.A(n_4624),
.Y(n_5259)
);

INVx2_ASAP7_75t_L g5260 ( 
.A(n_4924),
.Y(n_5260)
);

NOR2xp33_ASAP7_75t_L g5261 ( 
.A(n_4691),
.B(n_4286),
.Y(n_5261)
);

AOI21xp5_ASAP7_75t_L g5262 ( 
.A1(n_4786),
.A2(n_4359),
.B(n_4194),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_4651),
.Y(n_5263)
);

AND3x2_ASAP7_75t_L g5264 ( 
.A(n_4881),
.B(n_4575),
.C(n_4297),
.Y(n_5264)
);

BUFx6f_ASAP7_75t_L g5265 ( 
.A(n_5071),
.Y(n_5265)
);

OAI221xp5_ASAP7_75t_L g5266 ( 
.A1(n_4791),
.A2(n_4510),
.B1(n_4458),
.B2(n_4420),
.C(n_4428),
.Y(n_5266)
);

BUFx2_ASAP7_75t_L g5267 ( 
.A(n_4741),
.Y(n_5267)
);

OAI21xp33_ASAP7_75t_SL g5268 ( 
.A1(n_4586),
.A2(n_4640),
.B(n_4612),
.Y(n_5268)
);

OR2x2_ASAP7_75t_L g5269 ( 
.A(n_4655),
.B(n_4458),
.Y(n_5269)
);

INVx6_ASAP7_75t_L g5270 ( 
.A(n_5071),
.Y(n_5270)
);

AOI21xp5_ASAP7_75t_L g5271 ( 
.A1(n_4899),
.A2(n_4375),
.B(n_4368),
.Y(n_5271)
);

OAI21xp5_ASAP7_75t_L g5272 ( 
.A1(n_4791),
.A2(n_4076),
.B(n_4556),
.Y(n_5272)
);

AND2x4_ASAP7_75t_L g5273 ( 
.A(n_4600),
.B(n_4368),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_4767),
.B(n_4556),
.Y(n_5274)
);

OAI22xp5_ASAP7_75t_L g5275 ( 
.A1(n_4634),
.A2(n_4331),
.B1(n_4307),
.B2(n_4238),
.Y(n_5275)
);

AOI22xp33_ASAP7_75t_L g5276 ( 
.A1(n_4969),
.A2(n_3975),
.B1(n_4323),
.B2(n_4460),
.Y(n_5276)
);

AND2x2_ASAP7_75t_L g5277 ( 
.A(n_4738),
.B(n_4302),
.Y(n_5277)
);

OR2x2_ASAP7_75t_L g5278 ( 
.A(n_4655),
.B(n_4527),
.Y(n_5278)
);

OR2x6_ASAP7_75t_L g5279 ( 
.A(n_4594),
.B(n_4238),
.Y(n_5279)
);

BUFx10_ASAP7_75t_L g5280 ( 
.A(n_4624),
.Y(n_5280)
);

AOI21xp5_ASAP7_75t_L g5281 ( 
.A1(n_4899),
.A2(n_4375),
.B(n_4368),
.Y(n_5281)
);

OAI21x1_ASAP7_75t_L g5282 ( 
.A1(n_4883),
.A2(n_4464),
.B(n_4454),
.Y(n_5282)
);

NOR2xp33_ASAP7_75t_L g5283 ( 
.A(n_4691),
.B(n_4286),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_4651),
.Y(n_5284)
);

AOI32xp33_ASAP7_75t_L g5285 ( 
.A1(n_4640),
.A2(n_4576),
.A3(n_4574),
.B1(n_4524),
.B2(n_4459),
.Y(n_5285)
);

AO22x2_ASAP7_75t_L g5286 ( 
.A1(n_4690),
.A2(n_4464),
.B1(n_4491),
.B2(n_4481),
.Y(n_5286)
);

NOR2xp33_ASAP7_75t_SL g5287 ( 
.A(n_4665),
.B(n_4393),
.Y(n_5287)
);

HB1xp67_ASAP7_75t_L g5288 ( 
.A(n_4687),
.Y(n_5288)
);

INVx2_ASAP7_75t_L g5289 ( 
.A(n_4924),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_4653),
.Y(n_5290)
);

OAI21xp33_ASAP7_75t_L g5291 ( 
.A1(n_4640),
.A2(n_4445),
.B(n_4423),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_4653),
.Y(n_5292)
);

A2O1A1Ixp33_ASAP7_75t_L g5293 ( 
.A1(n_4676),
.A2(n_4008),
.B(n_4006),
.C(n_4393),
.Y(n_5293)
);

AOI22xp5_ASAP7_75t_L g5294 ( 
.A1(n_4793),
.A2(n_4323),
.B1(n_3975),
.B2(n_4331),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_4658),
.Y(n_5295)
);

OAI22xp5_ASAP7_75t_L g5296 ( 
.A1(n_4831),
.A2(n_4238),
.B1(n_4307),
.B2(n_4297),
.Y(n_5296)
);

AOI22xp5_ASAP7_75t_L g5297 ( 
.A1(n_4676),
.A2(n_4323),
.B1(n_4573),
.B2(n_4485),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_4658),
.Y(n_5298)
);

INVx2_ASAP7_75t_SL g5299 ( 
.A(n_4769),
.Y(n_5299)
);

AOI21xp5_ASAP7_75t_L g5300 ( 
.A1(n_4779),
.A2(n_4375),
.B(n_4368),
.Y(n_5300)
);

OR2x2_ASAP7_75t_L g5301 ( 
.A(n_4655),
.B(n_4457),
.Y(n_5301)
);

INVx2_ASAP7_75t_SL g5302 ( 
.A(n_4769),
.Y(n_5302)
);

NAND2x1p5_ASAP7_75t_L g5303 ( 
.A(n_5056),
.B(n_4994),
.Y(n_5303)
);

AOI21xp5_ASAP7_75t_L g5304 ( 
.A1(n_4779),
.A2(n_4385),
.B(n_4375),
.Y(n_5304)
);

OR2x6_ASAP7_75t_L g5305 ( 
.A(n_4594),
.B(n_4307),
.Y(n_5305)
);

AO21x2_ASAP7_75t_L g5306 ( 
.A1(n_5023),
.A2(n_4491),
.B(n_4481),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_4669),
.Y(n_5307)
);

OAI22xp5_ASAP7_75t_L g5308 ( 
.A1(n_4831),
.A2(n_4297),
.B1(n_4385),
.B2(n_4476),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_4669),
.Y(n_5309)
);

AOI21xp5_ASAP7_75t_L g5310 ( 
.A1(n_4618),
.A2(n_4385),
.B(n_4145),
.Y(n_5310)
);

NAND2xp5_ASAP7_75t_SL g5311 ( 
.A(n_4672),
.B(n_4553),
.Y(n_5311)
);

OAI221xp5_ASAP7_75t_L g5312 ( 
.A1(n_4791),
.A2(n_4496),
.B1(n_4508),
.B2(n_4480),
.C(n_4520),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_4685),
.Y(n_5313)
);

BUFx8_ASAP7_75t_L g5314 ( 
.A(n_5075),
.Y(n_5314)
);

AND2x2_ASAP7_75t_L g5315 ( 
.A(n_4739),
.B(n_4309),
.Y(n_5315)
);

NAND2xp5_ASAP7_75t_L g5316 ( 
.A(n_4752),
.B(n_4833),
.Y(n_5316)
);

INVx2_ASAP7_75t_L g5317 ( 
.A(n_4924),
.Y(n_5317)
);

OR2x2_ASAP7_75t_L g5318 ( 
.A(n_4839),
.B(n_4497),
.Y(n_5318)
);

BUFx10_ASAP7_75t_L g5319 ( 
.A(n_4769),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_4685),
.Y(n_5320)
);

BUFx2_ASAP7_75t_L g5321 ( 
.A(n_4741),
.Y(n_5321)
);

AOI22xp33_ASAP7_75t_L g5322 ( 
.A1(n_4969),
.A2(n_4323),
.B1(n_4530),
.B2(n_4544),
.Y(n_5322)
);

AND2x4_ASAP7_75t_L g5323 ( 
.A(n_4790),
.B(n_4385),
.Y(n_5323)
);

AOI21x1_ASAP7_75t_L g5324 ( 
.A1(n_5047),
.A2(n_4544),
.B(n_4530),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_4696),
.Y(n_5325)
);

CKINVDCx12_ASAP7_75t_R g5326 ( 
.A(n_5067),
.Y(n_5326)
);

INVx2_ASAP7_75t_L g5327 ( 
.A(n_4924),
.Y(n_5327)
);

AOI21xp5_ASAP7_75t_L g5328 ( 
.A1(n_4618),
.A2(n_4297),
.B(n_4573),
.Y(n_5328)
);

INVx1_ASAP7_75t_L g5329 ( 
.A(n_4696),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_4714),
.Y(n_5330)
);

OR2x2_ASAP7_75t_L g5331 ( 
.A(n_4839),
.B(n_4565),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_4714),
.Y(n_5332)
);

OR2x6_ASAP7_75t_L g5333 ( 
.A(n_4618),
.B(n_4573),
.Y(n_5333)
);

AND2x2_ASAP7_75t_L g5334 ( 
.A(n_4739),
.B(n_4309),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_4730),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_4730),
.Y(n_5336)
);

AND2x2_ASAP7_75t_L g5337 ( 
.A(n_4739),
.B(n_4311),
.Y(n_5337)
);

AND2x2_ASAP7_75t_L g5338 ( 
.A(n_4861),
.B(n_4311),
.Y(n_5338)
);

OAI221xp5_ASAP7_75t_L g5339 ( 
.A1(n_4791),
.A2(n_4545),
.B1(n_4571),
.B2(n_4565),
.C(n_4567),
.Y(n_5339)
);

OAI21x1_ASAP7_75t_L g5340 ( 
.A1(n_4883),
.A2(n_4545),
.B(n_4567),
.Y(n_5340)
);

NAND3xp33_ASAP7_75t_L g5341 ( 
.A(n_5025),
.B(n_4553),
.C(n_4063),
.Y(n_5341)
);

INVx1_ASAP7_75t_L g5342 ( 
.A(n_4617),
.Y(n_5342)
);

NAND2xp5_ASAP7_75t_L g5343 ( 
.A(n_4752),
.B(n_4574),
.Y(n_5343)
);

OA21x2_ASAP7_75t_L g5344 ( 
.A1(n_4886),
.A2(n_4798),
.B(n_4787),
.Y(n_5344)
);

AOI22xp33_ASAP7_75t_L g5345 ( 
.A1(n_4969),
.A2(n_4438),
.B1(n_4425),
.B2(n_3931),
.Y(n_5345)
);

BUFx4f_ASAP7_75t_SL g5346 ( 
.A(n_4704),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_4617),
.Y(n_5347)
);

INVxp67_ASAP7_75t_SL g5348 ( 
.A(n_4869),
.Y(n_5348)
);

AND2x2_ASAP7_75t_L g5349 ( 
.A(n_4861),
.B(n_4378),
.Y(n_5349)
);

BUFx3_ASAP7_75t_L g5350 ( 
.A(n_4704),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_4617),
.Y(n_5351)
);

AOI22xp33_ASAP7_75t_L g5352 ( 
.A1(n_4920),
.A2(n_4438),
.B1(n_3942),
.B2(n_3931),
.Y(n_5352)
);

AND2x2_ASAP7_75t_L g5353 ( 
.A(n_4861),
.B(n_4378),
.Y(n_5353)
);

AOI21xp5_ASAP7_75t_L g5354 ( 
.A1(n_4618),
.A2(n_4573),
.B(n_4575),
.Y(n_5354)
);

OAI21xp5_ASAP7_75t_L g5355 ( 
.A1(n_4676),
.A2(n_4076),
.B(n_4576),
.Y(n_5355)
);

INVx2_ASAP7_75t_SL g5356 ( 
.A(n_4769),
.Y(n_5356)
);

NAND2xp5_ASAP7_75t_L g5357 ( 
.A(n_4833),
.B(n_4403),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_4734),
.Y(n_5358)
);

NAND2xp5_ASAP7_75t_L g5359 ( 
.A(n_4711),
.B(n_4403),
.Y(n_5359)
);

AOI321xp33_ASAP7_75t_L g5360 ( 
.A1(n_4613),
.A2(n_4006),
.A3(n_4008),
.B1(n_4355),
.B2(n_4136),
.C(n_4389),
.Y(n_5360)
);

AO31x2_ASAP7_75t_L g5361 ( 
.A1(n_4891),
.A2(n_2509),
.A3(n_2415),
.B(n_2480),
.Y(n_5361)
);

AO31x2_ASAP7_75t_L g5362 ( 
.A1(n_4891),
.A2(n_2509),
.A3(n_2478),
.B(n_2473),
.Y(n_5362)
);

AOI21xp33_ASAP7_75t_L g5363 ( 
.A1(n_4584),
.A2(n_4493),
.B(n_4063),
.Y(n_5363)
);

NAND2xp5_ASAP7_75t_L g5364 ( 
.A(n_4711),
.B(n_4410),
.Y(n_5364)
);

INVx3_ASAP7_75t_L g5365 ( 
.A(n_4672),
.Y(n_5365)
);

AO31x2_ASAP7_75t_L g5366 ( 
.A1(n_4891),
.A2(n_2471),
.A3(n_2463),
.B(n_2460),
.Y(n_5366)
);

CKINVDCx5p33_ASAP7_75t_R g5367 ( 
.A(n_5074),
.Y(n_5367)
);

AND2x2_ASAP7_75t_L g5368 ( 
.A(n_4814),
.B(n_4410),
.Y(n_5368)
);

AOI221xp5_ASAP7_75t_L g5369 ( 
.A1(n_5023),
.A2(n_4006),
.B1(n_4008),
.B2(n_4524),
.C(n_4411),
.Y(n_5369)
);

INVx1_ASAP7_75t_L g5370 ( 
.A(n_4734),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_4736),
.Y(n_5371)
);

AOI21x1_ASAP7_75t_L g5372 ( 
.A1(n_4765),
.A2(n_4459),
.B(n_4411),
.Y(n_5372)
);

OR2x6_ASAP7_75t_L g5373 ( 
.A(n_4618),
.B(n_3860),
.Y(n_5373)
);

BUFx2_ASAP7_75t_L g5374 ( 
.A(n_4741),
.Y(n_5374)
);

AOI21xp5_ASAP7_75t_L g5375 ( 
.A1(n_4618),
.A2(n_4493),
.B(n_3905),
.Y(n_5375)
);

O2A1O1Ixp33_ASAP7_75t_L g5376 ( 
.A1(n_4584),
.A2(n_4008),
.B(n_4534),
.C(n_3942),
.Y(n_5376)
);

AOI21xp5_ASAP7_75t_L g5377 ( 
.A1(n_4821),
.A2(n_3860),
.B(n_3905),
.Y(n_5377)
);

OA21x2_ASAP7_75t_L g5378 ( 
.A1(n_4886),
.A2(n_4534),
.B(n_4532),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_4736),
.Y(n_5379)
);

OAI211xp5_ASAP7_75t_L g5380 ( 
.A1(n_4672),
.A2(n_4727),
.B(n_4838),
.C(n_4613),
.Y(n_5380)
);

A2O1A1Ixp33_ASAP7_75t_L g5381 ( 
.A1(n_5039),
.A2(n_4136),
.B(n_4125),
.C(n_3905),
.Y(n_5381)
);

NAND2xp5_ASAP7_75t_L g5382 ( 
.A(n_4925),
.B(n_4771),
.Y(n_5382)
);

INVxp67_ASAP7_75t_L g5383 ( 
.A(n_4925),
.Y(n_5383)
);

O2A1O1Ixp33_ASAP7_75t_L g5384 ( 
.A1(n_4584),
.A2(n_3931),
.B(n_4355),
.C(n_4013),
.Y(n_5384)
);

CKINVDCx6p67_ASAP7_75t_R g5385 ( 
.A(n_5075),
.Y(n_5385)
);

OAI21x1_ASAP7_75t_L g5386 ( 
.A1(n_5014),
.A2(n_2644),
.B(n_2792),
.Y(n_5386)
);

BUFx3_ASAP7_75t_L g5387 ( 
.A(n_4980),
.Y(n_5387)
);

AOI21xp5_ASAP7_75t_L g5388 ( 
.A1(n_4755),
.A2(n_5078),
.B(n_5063),
.Y(n_5388)
);

AOI21xp5_ASAP7_75t_L g5389 ( 
.A1(n_4755),
.A2(n_4572),
.B(n_4546),
.Y(n_5389)
);

INVx2_ASAP7_75t_L g5390 ( 
.A(n_4936),
.Y(n_5390)
);

INVx2_ASAP7_75t_SL g5391 ( 
.A(n_4769),
.Y(n_5391)
);

AOI22xp33_ASAP7_75t_L g5392 ( 
.A1(n_4920),
.A2(n_2460),
.B1(n_2455),
.B2(n_2471),
.Y(n_5392)
);

NAND2xp5_ASAP7_75t_SL g5393 ( 
.A(n_4672),
.B(n_4469),
.Y(n_5393)
);

OAI21xp5_ASAP7_75t_L g5394 ( 
.A1(n_4838),
.A2(n_4416),
.B(n_2605),
.Y(n_5394)
);

AO21x2_ASAP7_75t_L g5395 ( 
.A1(n_4936),
.A2(n_2463),
.B(n_2458),
.Y(n_5395)
);

AOI21xp5_ASAP7_75t_L g5396 ( 
.A1(n_5063),
.A2(n_4572),
.B(n_4038),
.Y(n_5396)
);

AOI21xp5_ASAP7_75t_L g5397 ( 
.A1(n_5078),
.A2(n_4572),
.B(n_4038),
.Y(n_5397)
);

INVx1_ASAP7_75t_L g5398 ( 
.A(n_4743),
.Y(n_5398)
);

AOI21xp5_ASAP7_75t_L g5399 ( 
.A1(n_4855),
.A2(n_4572),
.B(n_4038),
.Y(n_5399)
);

OR2x2_ASAP7_75t_L g5400 ( 
.A(n_4855),
.B(n_4355),
.Y(n_5400)
);

AOI211xp5_ASAP7_75t_L g5401 ( 
.A1(n_4672),
.A2(n_4727),
.B(n_4583),
.C(n_4589),
.Y(n_5401)
);

AO31x2_ASAP7_75t_L g5402 ( 
.A1(n_4663),
.A2(n_2458),
.A3(n_2454),
.B(n_2452),
.Y(n_5402)
);

AND2x2_ASAP7_75t_L g5403 ( 
.A(n_4814),
.B(n_4818),
.Y(n_5403)
);

OAI21x1_ASAP7_75t_L g5404 ( 
.A1(n_5014),
.A2(n_2748),
.B(n_2661),
.Y(n_5404)
);

HB1xp67_ASAP7_75t_L g5405 ( 
.A(n_4687),
.Y(n_5405)
);

AOI22xp33_ASAP7_75t_L g5406 ( 
.A1(n_4920),
.A2(n_2452),
.B1(n_2444),
.B2(n_2441),
.Y(n_5406)
);

OA21x2_ASAP7_75t_L g5407 ( 
.A1(n_4787),
.A2(n_4503),
.B(n_4507),
.Y(n_5407)
);

AND2x4_ASAP7_75t_L g5408 ( 
.A(n_4790),
.B(n_4355),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_4743),
.Y(n_5409)
);

AOI21xp5_ASAP7_75t_L g5410 ( 
.A1(n_4699),
.A2(n_4572),
.B(n_4384),
.Y(n_5410)
);

OAI21x1_ASAP7_75t_L g5411 ( 
.A1(n_5014),
.A2(n_2756),
.B(n_2797),
.Y(n_5411)
);

AOI21xp5_ASAP7_75t_L g5412 ( 
.A1(n_4699),
.A2(n_4563),
.B(n_4384),
.Y(n_5412)
);

NAND2xp5_ASAP7_75t_L g5413 ( 
.A(n_4771),
.B(n_4013),
.Y(n_5413)
);

NAND2x1p5_ASAP7_75t_L g5414 ( 
.A(n_5056),
.B(n_4994),
.Y(n_5414)
);

OA21x2_ASAP7_75t_L g5415 ( 
.A1(n_4798),
.A2(n_4503),
.B(n_4507),
.Y(n_5415)
);

AO31x2_ASAP7_75t_L g5416 ( 
.A1(n_4663),
.A2(n_2441),
.A3(n_2607),
.B(n_2611),
.Y(n_5416)
);

OAI21x1_ASAP7_75t_L g5417 ( 
.A1(n_5015),
.A2(n_2675),
.B(n_2797),
.Y(n_5417)
);

NAND2xp5_ASAP7_75t_L g5418 ( 
.A(n_4684),
.B(n_4013),
.Y(n_5418)
);

NAND2x1_ASAP7_75t_L g5419 ( 
.A(n_4966),
.B(n_4038),
.Y(n_5419)
);

AOI22xp33_ASAP7_75t_L g5420 ( 
.A1(n_4920),
.A2(n_2576),
.B1(n_2416),
.B2(n_2431),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_4625),
.Y(n_5421)
);

OAI22xp5_ASAP7_75t_L g5422 ( 
.A1(n_4998),
.A2(n_4384),
.B1(n_4293),
.B2(n_4179),
.Y(n_5422)
);

NAND2xp5_ASAP7_75t_L g5423 ( 
.A(n_4684),
.B(n_4013),
.Y(n_5423)
);

INVx2_ASAP7_75t_L g5424 ( 
.A(n_4936),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_4625),
.Y(n_5425)
);

OAI21x1_ASAP7_75t_L g5426 ( 
.A1(n_5015),
.A2(n_2661),
.B(n_2795),
.Y(n_5426)
);

OR2x2_ASAP7_75t_L g5427 ( 
.A(n_4632),
.B(n_4355),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_4625),
.Y(n_5428)
);

INVx2_ASAP7_75t_L g5429 ( 
.A(n_4940),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_4629),
.Y(n_5430)
);

AOI21xp5_ASAP7_75t_L g5431 ( 
.A1(n_4699),
.A2(n_4972),
.B(n_4822),
.Y(n_5431)
);

AO31x2_ASAP7_75t_L g5432 ( 
.A1(n_4663),
.A2(n_2656),
.A3(n_2820),
.B(n_2819),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_4629),
.Y(n_5433)
);

AND2x2_ASAP7_75t_L g5434 ( 
.A(n_4814),
.B(n_4188),
.Y(n_5434)
);

NAND2xp5_ASAP7_75t_L g5435 ( 
.A(n_4623),
.B(n_4013),
.Y(n_5435)
);

INVx4_ASAP7_75t_L g5436 ( 
.A(n_5075),
.Y(n_5436)
);

INVx1_ASAP7_75t_SL g5437 ( 
.A(n_4813),
.Y(n_5437)
);

NAND2xp5_ASAP7_75t_L g5438 ( 
.A(n_4623),
.B(n_4125),
.Y(n_5438)
);

BUFx3_ASAP7_75t_L g5439 ( 
.A(n_4980),
.Y(n_5439)
);

A2O1A1Ixp33_ASAP7_75t_L g5440 ( 
.A1(n_5039),
.A2(n_4136),
.B(n_4125),
.C(n_4324),
.Y(n_5440)
);

NAND2xp5_ASAP7_75t_L g5441 ( 
.A(n_4642),
.B(n_4125),
.Y(n_5441)
);

NOR2x1_ASAP7_75t_SL g5442 ( 
.A(n_4671),
.B(n_4063),
.Y(n_5442)
);

HB1xp67_ASAP7_75t_L g5443 ( 
.A(n_4582),
.Y(n_5443)
);

OA21x2_ASAP7_75t_L g5444 ( 
.A1(n_5015),
.A2(n_4503),
.B(n_4507),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_4629),
.Y(n_5445)
);

OR2x6_ASAP7_75t_L g5446 ( 
.A(n_4671),
.B(n_4063),
.Y(n_5446)
);

AND2x2_ASAP7_75t_L g5447 ( 
.A(n_4818),
.B(n_4188),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_4678),
.Y(n_5448)
);

AOI21xp5_ASAP7_75t_L g5449 ( 
.A1(n_4972),
.A2(n_4563),
.B(n_4384),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_4678),
.Y(n_5450)
);

AOI22xp33_ASAP7_75t_L g5451 ( 
.A1(n_4920),
.A2(n_2576),
.B1(n_2416),
.B2(n_2431),
.Y(n_5451)
);

NAND2xp5_ASAP7_75t_L g5452 ( 
.A(n_4642),
.B(n_4125),
.Y(n_5452)
);

A2O1A1Ixp33_ASAP7_75t_L g5453 ( 
.A1(n_5039),
.A2(n_4136),
.B(n_4328),
.C(n_4324),
.Y(n_5453)
);

BUFx3_ASAP7_75t_L g5454 ( 
.A(n_5075),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_4678),
.Y(n_5455)
);

INVx1_ASAP7_75t_L g5456 ( 
.A(n_4702),
.Y(n_5456)
);

INVx1_ASAP7_75t_L g5457 ( 
.A(n_4702),
.Y(n_5457)
);

AOI22xp33_ASAP7_75t_L g5458 ( 
.A1(n_5033),
.A2(n_2576),
.B1(n_2416),
.B2(n_2431),
.Y(n_5458)
);

OAI211xp5_ASAP7_75t_L g5459 ( 
.A1(n_4727),
.A2(n_4563),
.B(n_4116),
.C(n_4071),
.Y(n_5459)
);

INVx2_ASAP7_75t_L g5460 ( 
.A(n_4940),
.Y(n_5460)
);

OAI22xp5_ASAP7_75t_L g5461 ( 
.A1(n_4998),
.A2(n_4071),
.B1(n_4113),
.B2(n_4116),
.Y(n_5461)
);

INVx2_ASAP7_75t_SL g5462 ( 
.A(n_4769),
.Y(n_5462)
);

NOR2xp67_ASAP7_75t_L g5463 ( 
.A(n_5006),
.B(n_4063),
.Y(n_5463)
);

INVx2_ASAP7_75t_L g5464 ( 
.A(n_4940),
.Y(n_5464)
);

NAND2xp5_ASAP7_75t_L g5465 ( 
.A(n_4923),
.B(n_4296),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_4702),
.Y(n_5466)
);

OAI22xp5_ASAP7_75t_L g5467 ( 
.A1(n_4902),
.A2(n_4563),
.B1(n_4069),
.B2(n_4071),
.Y(n_5467)
);

AOI21xp5_ASAP7_75t_L g5468 ( 
.A1(n_4822),
.A2(n_4563),
.B(n_4069),
.Y(n_5468)
);

NAND2xp5_ASAP7_75t_L g5469 ( 
.A(n_4923),
.B(n_4296),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_4705),
.Y(n_5470)
);

AND2x2_ASAP7_75t_L g5471 ( 
.A(n_4818),
.B(n_4188),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_4746),
.Y(n_5472)
);

OA21x2_ASAP7_75t_L g5473 ( 
.A1(n_5022),
.A2(n_4503),
.B(n_4532),
.Y(n_5473)
);

AOI21xp5_ASAP7_75t_L g5474 ( 
.A1(n_4877),
.A2(n_4113),
.B(n_4384),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_4746),
.Y(n_5475)
);

OAI21xp5_ASAP7_75t_L g5476 ( 
.A1(n_5025),
.A2(n_4416),
.B(n_2605),
.Y(n_5476)
);

INVx2_ASAP7_75t_L g5477 ( 
.A(n_4940),
.Y(n_5477)
);

INVx1_ASAP7_75t_L g5478 ( 
.A(n_4749),
.Y(n_5478)
);

AOI21xp5_ASAP7_75t_L g5479 ( 
.A1(n_4877),
.A2(n_4113),
.B(n_4430),
.Y(n_5479)
);

AOI21xp5_ASAP7_75t_L g5480 ( 
.A1(n_4583),
.A2(n_4113),
.B(n_4430),
.Y(n_5480)
);

OAI22xp33_ASAP7_75t_L g5481 ( 
.A1(n_4727),
.A2(n_4116),
.B1(n_4069),
.B2(n_4071),
.Y(n_5481)
);

AOI21xp5_ASAP7_75t_L g5482 ( 
.A1(n_4589),
.A2(n_4113),
.B(n_4430),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_4749),
.Y(n_5483)
);

INVx4_ASAP7_75t_L g5484 ( 
.A(n_5031),
.Y(n_5484)
);

AOI22xp33_ASAP7_75t_L g5485 ( 
.A1(n_5033),
.A2(n_2565),
.B1(n_2416),
.B2(n_2431),
.Y(n_5485)
);

AOI21xp5_ASAP7_75t_L g5486 ( 
.A1(n_4851),
.A2(n_4293),
.B(n_4509),
.Y(n_5486)
);

OAI22xp33_ASAP7_75t_L g5487 ( 
.A1(n_4727),
.A2(n_4116),
.B1(n_4069),
.B2(n_4071),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_4753),
.Y(n_5488)
);

BUFx6f_ASAP7_75t_L g5489 ( 
.A(n_4762),
.Y(n_5489)
);

NAND2xp5_ASAP7_75t_L g5490 ( 
.A(n_4889),
.B(n_4296),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_4753),
.Y(n_5491)
);

BUFx2_ASAP7_75t_L g5492 ( 
.A(n_4741),
.Y(n_5492)
);

INVx1_ASAP7_75t_L g5493 ( 
.A(n_4785),
.Y(n_5493)
);

AND2x2_ASAP7_75t_L g5494 ( 
.A(n_4639),
.B(n_4069),
.Y(n_5494)
);

INVx5_ASAP7_75t_L g5495 ( 
.A(n_4762),
.Y(n_5495)
);

INVx2_ASAP7_75t_L g5496 ( 
.A(n_4947),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_4785),
.Y(n_5497)
);

AND2x4_ASAP7_75t_L g5498 ( 
.A(n_4741),
.B(n_4324),
.Y(n_5498)
);

AOI221xp5_ASAP7_75t_L g5499 ( 
.A1(n_4727),
.A2(n_4503),
.B1(n_4532),
.B2(n_4507),
.C(n_4324),
.Y(n_5499)
);

BUFx8_ASAP7_75t_L g5500 ( 
.A(n_5050),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_4889),
.B(n_4296),
.Y(n_5501)
);

OAI21xp5_ASAP7_75t_L g5502 ( 
.A1(n_4943),
.A2(n_4416),
.B(n_4136),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_4808),
.Y(n_5503)
);

CKINVDCx5p33_ASAP7_75t_R g5504 ( 
.A(n_4996),
.Y(n_5504)
);

INVx4_ASAP7_75t_SL g5505 ( 
.A(n_5031),
.Y(n_5505)
);

AOI22xp5_ASAP7_75t_L g5506 ( 
.A1(n_5033),
.A2(n_4509),
.B1(n_4116),
.B2(n_4167),
.Y(n_5506)
);

AOI21xp5_ASAP7_75t_L g5507 ( 
.A1(n_4851),
.A2(n_4167),
.B(n_4179),
.Y(n_5507)
);

HB1xp67_ASAP7_75t_L g5508 ( 
.A(n_4582),
.Y(n_5508)
);

CKINVDCx6p67_ASAP7_75t_R g5509 ( 
.A(n_5031),
.Y(n_5509)
);

AOI21xp5_ASAP7_75t_L g5510 ( 
.A1(n_4851),
.A2(n_4167),
.B(n_4179),
.Y(n_5510)
);

NOR2xp33_ASAP7_75t_L g5511 ( 
.A(n_5031),
.B(n_4167),
.Y(n_5511)
);

INVx2_ASAP7_75t_L g5512 ( 
.A(n_4947),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_4808),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_4811),
.Y(n_5514)
);

AOI21xp5_ASAP7_75t_L g5515 ( 
.A1(n_4744),
.A2(n_4943),
.B(n_4674),
.Y(n_5515)
);

AO31x2_ASAP7_75t_L g5516 ( 
.A1(n_4947),
.A2(n_4963),
.A3(n_4999),
.B(n_4956),
.Y(n_5516)
);

INVx2_ASAP7_75t_L g5517 ( 
.A(n_4947),
.Y(n_5517)
);

AND2x4_ASAP7_75t_L g5518 ( 
.A(n_4741),
.B(n_4803),
.Y(n_5518)
);

INVx2_ASAP7_75t_L g5519 ( 
.A(n_4956),
.Y(n_5519)
);

AOI21xp5_ASAP7_75t_L g5520 ( 
.A1(n_4744),
.A2(n_4167),
.B(n_4179),
.Y(n_5520)
);

AOI21xp5_ASAP7_75t_L g5521 ( 
.A1(n_4943),
.A2(n_4509),
.B(n_4179),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_4811),
.Y(n_5522)
);

AOI21xp5_ASAP7_75t_L g5523 ( 
.A1(n_4674),
.A2(n_4293),
.B(n_4430),
.Y(n_5523)
);

AOI21xp5_ASAP7_75t_L g5524 ( 
.A1(n_4674),
.A2(n_4293),
.B(n_4430),
.Y(n_5524)
);

AOI21x1_ASAP7_75t_L g5525 ( 
.A1(n_4765),
.A2(n_4507),
.B(n_4532),
.Y(n_5525)
);

NAND2xp5_ASAP7_75t_L g5526 ( 
.A(n_4900),
.B(n_4296),
.Y(n_5526)
);

OAI221xp5_ASAP7_75t_L g5527 ( 
.A1(n_4727),
.A2(n_4509),
.B1(n_4546),
.B2(n_4293),
.C(n_4324),
.Y(n_5527)
);

OA21x2_ASAP7_75t_L g5528 ( 
.A1(n_5022),
.A2(n_4532),
.B(n_4147),
.Y(n_5528)
);

AOI221xp5_ASAP7_75t_L g5529 ( 
.A1(n_4598),
.A2(n_4328),
.B1(n_4546),
.B2(n_4509),
.C(n_4551),
.Y(n_5529)
);

NAND2xp5_ASAP7_75t_L g5530 ( 
.A(n_4900),
.B(n_3841),
.Y(n_5530)
);

AND2x2_ASAP7_75t_L g5531 ( 
.A(n_4639),
.B(n_4546),
.Y(n_5531)
);

OR2x6_ASAP7_75t_L g5532 ( 
.A(n_4671),
.B(n_4546),
.Y(n_5532)
);

NAND2xp5_ASAP7_75t_L g5533 ( 
.A(n_4632),
.B(n_3841),
.Y(n_5533)
);

AOI22xp5_ASAP7_75t_L g5534 ( 
.A1(n_5033),
.A2(n_3538),
.B1(n_3734),
.B2(n_3759),
.Y(n_5534)
);

NOR2xp33_ASAP7_75t_L g5535 ( 
.A(n_5050),
.B(n_4965),
.Y(n_5535)
);

AOI22xp5_ASAP7_75t_SL g5536 ( 
.A1(n_4965),
.A2(n_3538),
.B1(n_3759),
.B2(n_3887),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_4852),
.Y(n_5537)
);

OA21x2_ASAP7_75t_L g5538 ( 
.A1(n_5022),
.A2(n_4616),
.B(n_4690),
.Y(n_5538)
);

NAND2xp5_ASAP7_75t_L g5539 ( 
.A(n_4643),
.B(n_3841),
.Y(n_5539)
);

A2O1A1Ixp33_ASAP7_75t_L g5540 ( 
.A1(n_4902),
.A2(n_4328),
.B(n_4036),
.C(n_4056),
.Y(n_5540)
);

AOI21xp5_ASAP7_75t_L g5541 ( 
.A1(n_4674),
.A2(n_3759),
.B(n_3887),
.Y(n_5541)
);

AOI22xp33_ASAP7_75t_L g5542 ( 
.A1(n_5033),
.A2(n_2604),
.B1(n_2416),
.B2(n_2431),
.Y(n_5542)
);

INVx2_ASAP7_75t_L g5543 ( 
.A(n_4956),
.Y(n_5543)
);

AND2x2_ASAP7_75t_L g5544 ( 
.A(n_4639),
.B(n_4416),
.Y(n_5544)
);

AOI22xp33_ASAP7_75t_L g5545 ( 
.A1(n_5018),
.A2(n_2604),
.B1(n_2431),
.B2(n_2435),
.Y(n_5545)
);

AND2x2_ASAP7_75t_L g5546 ( 
.A(n_4639),
.B(n_4416),
.Y(n_5546)
);

INVx2_ASAP7_75t_L g5547 ( 
.A(n_4963),
.Y(n_5547)
);

AOI211xp5_ASAP7_75t_SL g5548 ( 
.A1(n_5024),
.A2(n_4562),
.B(n_4313),
.C(n_4304),
.Y(n_5548)
);

AOI21xp5_ASAP7_75t_L g5549 ( 
.A1(n_4674),
.A2(n_3887),
.B(n_3903),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_4705),
.Y(n_5550)
);

INVx4_ASAP7_75t_L g5551 ( 
.A(n_5050),
.Y(n_5551)
);

OA21x2_ASAP7_75t_L g5552 ( 
.A1(n_4616),
.A2(n_4147),
.B(n_4148),
.Y(n_5552)
);

AOI22xp33_ASAP7_75t_L g5553 ( 
.A1(n_5018),
.A2(n_2598),
.B1(n_2435),
.B2(n_2448),
.Y(n_5553)
);

AOI22xp33_ASAP7_75t_L g5554 ( 
.A1(n_5018),
.A2(n_2591),
.B1(n_2435),
.B2(n_2448),
.Y(n_5554)
);

INVx1_ASAP7_75t_L g5555 ( 
.A(n_4852),
.Y(n_5555)
);

NAND2xp5_ASAP7_75t_L g5556 ( 
.A(n_4643),
.B(n_3841),
.Y(n_5556)
);

OAI21x1_ASAP7_75t_SL g5557 ( 
.A1(n_4966),
.A2(n_4562),
.B(n_3953),
.Y(n_5557)
);

NAND2x1p5_ASAP7_75t_L g5558 ( 
.A(n_5056),
.B(n_3538),
.Y(n_5558)
);

INVx2_ASAP7_75t_L g5559 ( 
.A(n_4963),
.Y(n_5559)
);

AND2x4_ASAP7_75t_L g5560 ( 
.A(n_4803),
.B(n_4960),
.Y(n_5560)
);

NAND3xp33_ASAP7_75t_L g5561 ( 
.A(n_4979),
.B(n_3734),
.C(n_3759),
.Y(n_5561)
);

AOI22xp33_ASAP7_75t_L g5562 ( 
.A1(n_5018),
.A2(n_2591),
.B1(n_2435),
.B2(n_2448),
.Y(n_5562)
);

AOI22xp33_ASAP7_75t_L g5563 ( 
.A1(n_5018),
.A2(n_2591),
.B1(n_2435),
.B2(n_2448),
.Y(n_5563)
);

OR2x2_ASAP7_75t_L g5564 ( 
.A(n_4870),
.B(n_4328),
.Y(n_5564)
);

AND2x2_ASAP7_75t_L g5565 ( 
.A(n_4639),
.B(n_4328),
.Y(n_5565)
);

NAND2xp5_ASAP7_75t_L g5566 ( 
.A(n_4997),
.B(n_3564),
.Y(n_5566)
);

AOI21xp5_ASAP7_75t_L g5567 ( 
.A1(n_5016),
.A2(n_3759),
.B(n_3887),
.Y(n_5567)
);

CKINVDCx12_ASAP7_75t_R g5568 ( 
.A(n_4682),
.Y(n_5568)
);

INVx8_ASAP7_75t_L g5569 ( 
.A(n_5049),
.Y(n_5569)
);

INVx3_ASAP7_75t_L g5570 ( 
.A(n_4580),
.Y(n_5570)
);

AND2x2_ASAP7_75t_L g5571 ( 
.A(n_4673),
.B(n_4277),
.Y(n_5571)
);

HB1xp67_ASAP7_75t_L g5572 ( 
.A(n_4774),
.Y(n_5572)
);

OR2x6_ASAP7_75t_L g5573 ( 
.A(n_4605),
.B(n_4666),
.Y(n_5573)
);

NAND2xp5_ASAP7_75t_L g5574 ( 
.A(n_4997),
.B(n_3564),
.Y(n_5574)
);

NAND3xp33_ASAP7_75t_L g5575 ( 
.A(n_4979),
.B(n_3734),
.C(n_3759),
.Y(n_5575)
);

NAND2xp5_ASAP7_75t_L g5576 ( 
.A(n_4577),
.B(n_3564),
.Y(n_5576)
);

NAND2xp5_ASAP7_75t_L g5577 ( 
.A(n_4577),
.B(n_3564),
.Y(n_5577)
);

OAI22xp33_ASAP7_75t_L g5578 ( 
.A1(n_4578),
.A2(n_3903),
.B1(n_3887),
.B2(n_3734),
.Y(n_5578)
);

BUFx12f_ASAP7_75t_L g5579 ( 
.A(n_4700),
.Y(n_5579)
);

INVx2_ASAP7_75t_L g5580 ( 
.A(n_4963),
.Y(n_5580)
);

AOI21xp5_ASAP7_75t_L g5581 ( 
.A1(n_5016),
.A2(n_3734),
.B(n_3903),
.Y(n_5581)
);

NAND2xp5_ASAP7_75t_L g5582 ( 
.A(n_4903),
.B(n_3564),
.Y(n_5582)
);

AOI21xp5_ASAP7_75t_L g5583 ( 
.A1(n_4949),
.A2(n_3734),
.B(n_3903),
.Y(n_5583)
);

AND2x2_ASAP7_75t_L g5584 ( 
.A(n_4673),
.B(n_4277),
.Y(n_5584)
);

OAI21xp5_ASAP7_75t_L g5585 ( 
.A1(n_4774),
.A2(n_4036),
.B(n_4056),
.Y(n_5585)
);

INVx1_ASAP7_75t_L g5586 ( 
.A(n_4862),
.Y(n_5586)
);

NOR2x1_ASAP7_75t_SL g5587 ( 
.A(n_4961),
.B(n_3903),
.Y(n_5587)
);

OAI21x1_ASAP7_75t_L g5588 ( 
.A1(n_4988),
.A2(n_4616),
.B(n_4865),
.Y(n_5588)
);

AOI21xp5_ASAP7_75t_L g5589 ( 
.A1(n_4949),
.A2(n_2612),
.B(n_2722),
.Y(n_5589)
);

AOI22xp33_ASAP7_75t_SL g5590 ( 
.A1(n_4747),
.A2(n_3696),
.B1(n_3710),
.B2(n_4036),
.Y(n_5590)
);

OAI22xp33_ASAP7_75t_L g5591 ( 
.A1(n_4578),
.A2(n_2576),
.B1(n_2435),
.B2(n_2448),
.Y(n_5591)
);

OAI222xp33_ASAP7_75t_L g5592 ( 
.A1(n_4598),
.A2(n_4670),
.B1(n_4599),
.B2(n_4649),
.C1(n_4645),
.C2(n_4690),
.Y(n_5592)
);

OR2x6_ASAP7_75t_L g5593 ( 
.A(n_4605),
.B(n_2435),
.Y(n_5593)
);

NOR2x1_ASAP7_75t_R g5594 ( 
.A(n_4996),
.B(n_2612),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_4862),
.Y(n_5595)
);

HB1xp67_ASAP7_75t_L g5596 ( 
.A(n_4895),
.Y(n_5596)
);

NOR2xp33_ASAP7_75t_L g5597 ( 
.A(n_4682),
.B(n_4715),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_4864),
.Y(n_5598)
);

AOI21xp5_ASAP7_75t_L g5599 ( 
.A1(n_4961),
.A2(n_2612),
.B(n_2647),
.Y(n_5599)
);

AOI21xp5_ASAP7_75t_L g5600 ( 
.A1(n_4961),
.A2(n_2612),
.B(n_2647),
.Y(n_5600)
);

AND2x4_ASAP7_75t_L g5601 ( 
.A(n_4803),
.B(n_4056),
.Y(n_5601)
);

NAND2xp5_ASAP7_75t_L g5602 ( 
.A(n_4903),
.B(n_3564),
.Y(n_5602)
);

INVx4_ASAP7_75t_L g5603 ( 
.A(n_4700),
.Y(n_5603)
);

CKINVDCx5p33_ASAP7_75t_R g5604 ( 
.A(n_4800),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_4705),
.Y(n_5605)
);

NAND2xp5_ASAP7_75t_L g5606 ( 
.A(n_4860),
.B(n_4830),
.Y(n_5606)
);

OAI22xp5_ASAP7_75t_L g5607 ( 
.A1(n_4578),
.A2(n_4661),
.B1(n_4721),
.B2(n_4657),
.Y(n_5607)
);

INVx2_ASAP7_75t_L g5608 ( 
.A(n_5028),
.Y(n_5608)
);

AOI21xp5_ASAP7_75t_L g5609 ( 
.A1(n_4961),
.A2(n_2647),
.B(n_2696),
.Y(n_5609)
);

INVx2_ASAP7_75t_L g5610 ( 
.A(n_5028),
.Y(n_5610)
);

NOR2xp33_ASAP7_75t_L g5611 ( 
.A(n_4715),
.B(n_4905),
.Y(n_5611)
);

AND2x2_ASAP7_75t_L g5612 ( 
.A(n_4673),
.B(n_4277),
.Y(n_5612)
);

NAND2xp5_ASAP7_75t_L g5613 ( 
.A(n_4860),
.B(n_3596),
.Y(n_5613)
);

AOI22xp33_ASAP7_75t_SL g5614 ( 
.A1(n_4747),
.A2(n_3710),
.B1(n_3696),
.B2(n_4056),
.Y(n_5614)
);

NAND2xp5_ASAP7_75t_L g5615 ( 
.A(n_4830),
.B(n_3596),
.Y(n_5615)
);

AOI22xp33_ASAP7_75t_L g5616 ( 
.A1(n_5018),
.A2(n_5044),
.B1(n_5038),
.B2(n_4991),
.Y(n_5616)
);

AOI21xp5_ASAP7_75t_L g5617 ( 
.A1(n_4961),
.A2(n_2647),
.B(n_2696),
.Y(n_5617)
);

AND2x4_ASAP7_75t_L g5618 ( 
.A(n_4803),
.B(n_4056),
.Y(n_5618)
);

NOR2xp67_ASAP7_75t_L g5619 ( 
.A(n_5006),
.B(n_2647),
.Y(n_5619)
);

OA21x2_ASAP7_75t_L g5620 ( 
.A1(n_4690),
.A2(n_4147),
.B(n_4148),
.Y(n_5620)
);

AOI21xp5_ASAP7_75t_L g5621 ( 
.A1(n_4961),
.A2(n_2647),
.B(n_2696),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_4864),
.Y(n_5622)
);

INVx2_ASAP7_75t_L g5623 ( 
.A(n_5037),
.Y(n_5623)
);

AOI21x1_ASAP7_75t_L g5624 ( 
.A1(n_4698),
.A2(n_2780),
.B(n_2661),
.Y(n_5624)
);

INVx2_ASAP7_75t_L g5625 ( 
.A(n_5037),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_4875),
.Y(n_5626)
);

AOI21xp5_ASAP7_75t_L g5627 ( 
.A1(n_4961),
.A2(n_2696),
.B(n_2722),
.Y(n_5627)
);

NAND2xp5_ASAP7_75t_L g5628 ( 
.A(n_4654),
.B(n_3596),
.Y(n_5628)
);

AOI21xp5_ASAP7_75t_L g5629 ( 
.A1(n_4955),
.A2(n_5070),
.B(n_4919),
.Y(n_5629)
);

AND2x2_ASAP7_75t_L g5630 ( 
.A(n_4673),
.B(n_4313),
.Y(n_5630)
);

AOI22xp33_ASAP7_75t_L g5631 ( 
.A1(n_5038),
.A2(n_2591),
.B1(n_2435),
.B2(n_2448),
.Y(n_5631)
);

NAND2xp5_ASAP7_75t_L g5632 ( 
.A(n_4654),
.B(n_3596),
.Y(n_5632)
);

HB1xp67_ASAP7_75t_L g5633 ( 
.A(n_4895),
.Y(n_5633)
);

A2O1A1Ixp33_ASAP7_75t_L g5634 ( 
.A1(n_4578),
.A2(n_4661),
.B(n_5040),
.C(n_4910),
.Y(n_5634)
);

AOI22xp33_ASAP7_75t_L g5635 ( 
.A1(n_5038),
.A2(n_2591),
.B1(n_2457),
.B2(n_2474),
.Y(n_5635)
);

AOI21xp5_ASAP7_75t_SL g5636 ( 
.A1(n_4989),
.A2(n_2722),
.B(n_2696),
.Y(n_5636)
);

INVx2_ASAP7_75t_SL g5637 ( 
.A(n_5049),
.Y(n_5637)
);

NOR2xp33_ASAP7_75t_L g5638 ( 
.A(n_4905),
.B(n_3791),
.Y(n_5638)
);

AND2x4_ASAP7_75t_L g5639 ( 
.A(n_4803),
.B(n_4147),
.Y(n_5639)
);

AOI22xp33_ASAP7_75t_L g5640 ( 
.A1(n_5038),
.A2(n_2565),
.B1(n_2457),
.B2(n_2474),
.Y(n_5640)
);

AOI22xp33_ASAP7_75t_L g5641 ( 
.A1(n_5091),
.A2(n_4867),
.B1(n_4882),
.B2(n_4648),
.Y(n_5641)
);

CKINVDCx5p33_ASAP7_75t_R g5642 ( 
.A(n_5219),
.Y(n_5642)
);

BUFx3_ASAP7_75t_L g5643 ( 
.A(n_5210),
.Y(n_5643)
);

NOR2xp33_ASAP7_75t_R g5644 ( 
.A(n_5326),
.B(n_4775),
.Y(n_5644)
);

NAND2xp5_ASAP7_75t_L g5645 ( 
.A(n_5106),
.B(n_4693),
.Y(n_5645)
);

NAND2xp5_ASAP7_75t_L g5646 ( 
.A(n_5606),
.B(n_4693),
.Y(n_5646)
);

INVx2_ASAP7_75t_L g5647 ( 
.A(n_5223),
.Y(n_5647)
);

INVx2_ASAP7_75t_L g5648 ( 
.A(n_5223),
.Y(n_5648)
);

OAI21x1_ASAP7_75t_L g5649 ( 
.A1(n_5227),
.A2(n_4994),
.B(n_4948),
.Y(n_5649)
);

NAND2xp5_ASAP7_75t_L g5650 ( 
.A(n_5382),
.B(n_4955),
.Y(n_5650)
);

OAI21xp5_ASAP7_75t_SL g5651 ( 
.A1(n_5431),
.A2(n_5228),
.B(n_5083),
.Y(n_5651)
);

CKINVDCx16_ASAP7_75t_R g5652 ( 
.A(n_5210),
.Y(n_5652)
);

NOR3xp33_ASAP7_75t_SL g5653 ( 
.A(n_5125),
.B(n_4775),
.C(n_4800),
.Y(n_5653)
);

OR2x6_ASAP7_75t_L g5654 ( 
.A(n_5207),
.B(n_5049),
.Y(n_5654)
);

NAND2xp5_ASAP7_75t_L g5655 ( 
.A(n_5348),
.B(n_4803),
.Y(n_5655)
);

OAI22xp5_ASAP7_75t_L g5656 ( 
.A1(n_5222),
.A2(n_4661),
.B1(n_4721),
.B2(n_4657),
.Y(n_5656)
);

NOR2xp33_ASAP7_75t_SL g5657 ( 
.A(n_5238),
.B(n_5125),
.Y(n_5657)
);

INVx2_ASAP7_75t_SL g5658 ( 
.A(n_5238),
.Y(n_5658)
);

OR2x2_ASAP7_75t_L g5659 ( 
.A(n_5183),
.B(n_4870),
.Y(n_5659)
);

OAI22xp5_ASAP7_75t_L g5660 ( 
.A1(n_5220),
.A2(n_4661),
.B1(n_4721),
.B2(n_4657),
.Y(n_5660)
);

AO31x2_ASAP7_75t_L g5661 ( 
.A1(n_5189),
.A2(n_4717),
.A3(n_4719),
.B(n_4698),
.Y(n_5661)
);

NAND2xp5_ASAP7_75t_L g5662 ( 
.A(n_5126),
.B(n_4803),
.Y(n_5662)
);

NAND2xp5_ASAP7_75t_SL g5663 ( 
.A(n_5257),
.B(n_5056),
.Y(n_5663)
);

INVx3_ASAP7_75t_L g5664 ( 
.A(n_5323),
.Y(n_5664)
);

CKINVDCx16_ASAP7_75t_R g5665 ( 
.A(n_5218),
.Y(n_5665)
);

INVx2_ASAP7_75t_L g5666 ( 
.A(n_5223),
.Y(n_5666)
);

NOR2xp33_ASAP7_75t_L g5667 ( 
.A(n_5568),
.B(n_4926),
.Y(n_5667)
);

NAND2xp33_ASAP7_75t_R g5668 ( 
.A(n_5367),
.B(n_4979),
.Y(n_5668)
);

NAND2xp5_ASAP7_75t_SL g5669 ( 
.A(n_5257),
.B(n_5056),
.Y(n_5669)
);

OR2x6_ASAP7_75t_L g5670 ( 
.A(n_5207),
.B(n_5049),
.Y(n_5670)
);

OR2x6_ASAP7_75t_L g5671 ( 
.A(n_5270),
.B(n_5049),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_5572),
.Y(n_5672)
);

NOR2xp33_ASAP7_75t_R g5673 ( 
.A(n_5326),
.B(n_4946),
.Y(n_5673)
);

AOI22xp33_ASAP7_75t_L g5674 ( 
.A1(n_5225),
.A2(n_4867),
.B1(n_4882),
.B2(n_4648),
.Y(n_5674)
);

INVx2_ASAP7_75t_L g5675 ( 
.A(n_5402),
.Y(n_5675)
);

HB1xp67_ASAP7_75t_L g5676 ( 
.A(n_5233),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_5596),
.Y(n_5677)
);

AOI22xp33_ASAP7_75t_SL g5678 ( 
.A1(n_5380),
.A2(n_5030),
.B1(n_4747),
.B2(n_4599),
.Y(n_5678)
);

NAND3xp33_ASAP7_75t_SL g5679 ( 
.A(n_5401),
.B(n_4813),
.C(n_4881),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5633),
.Y(n_5680)
);

OR2x6_ASAP7_75t_L g5681 ( 
.A(n_5270),
.B(n_5049),
.Y(n_5681)
);

HB1xp67_ASAP7_75t_L g5682 ( 
.A(n_5233),
.Y(n_5682)
);

NOR2xp33_ASAP7_75t_R g5683 ( 
.A(n_5568),
.B(n_4946),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_5099),
.Y(n_5684)
);

OAI22xp5_ASAP7_75t_L g5685 ( 
.A1(n_5209),
.A2(n_4960),
.B1(n_4944),
.B2(n_4817),
.Y(n_5685)
);

INVx4_ASAP7_75t_L g5686 ( 
.A(n_5579),
.Y(n_5686)
);

BUFx6f_ASAP7_75t_L g5687 ( 
.A(n_5082),
.Y(n_5687)
);

CKINVDCx16_ASAP7_75t_R g5688 ( 
.A(n_5287),
.Y(n_5688)
);

NOR2xp33_ASAP7_75t_R g5689 ( 
.A(n_5158),
.B(n_5049),
.Y(n_5689)
);

OR2x2_ASAP7_75t_L g5690 ( 
.A(n_5184),
.B(n_4880),
.Y(n_5690)
);

INVx3_ASAP7_75t_L g5691 ( 
.A(n_5323),
.Y(n_5691)
);

NOR2xp33_ASAP7_75t_R g5692 ( 
.A(n_5158),
.B(n_4622),
.Y(n_5692)
);

AND2x2_ASAP7_75t_L g5693 ( 
.A(n_5145),
.B(n_4622),
.Y(n_5693)
);

NAND2xp5_ASAP7_75t_L g5694 ( 
.A(n_5150),
.B(n_4803),
.Y(n_5694)
);

AOI22xp33_ASAP7_75t_L g5695 ( 
.A1(n_5110),
.A2(n_4867),
.B1(n_4882),
.B2(n_4648),
.Y(n_5695)
);

AO31x2_ASAP7_75t_L g5696 ( 
.A1(n_5293),
.A2(n_4717),
.A3(n_4719),
.B(n_4698),
.Y(n_5696)
);

INVxp67_ASAP7_75t_SL g5697 ( 
.A(n_5181),
.Y(n_5697)
);

AO31x2_ASAP7_75t_L g5698 ( 
.A1(n_5293),
.A2(n_4717),
.A3(n_4719),
.B(n_4698),
.Y(n_5698)
);

AOI22xp33_ASAP7_75t_SL g5699 ( 
.A1(n_5434),
.A2(n_5030),
.B1(n_4747),
.B2(n_4599),
.Y(n_5699)
);

HB1xp67_ASAP7_75t_L g5700 ( 
.A(n_5237),
.Y(n_5700)
);

OAI21xp5_ASAP7_75t_L g5701 ( 
.A1(n_5515),
.A2(n_4719),
.B(n_4717),
.Y(n_5701)
);

INVx2_ASAP7_75t_L g5702 ( 
.A(n_5402),
.Y(n_5702)
);

BUFx8_ASAP7_75t_L g5703 ( 
.A(n_5579),
.Y(n_5703)
);

CKINVDCx16_ASAP7_75t_R g5704 ( 
.A(n_5258),
.Y(n_5704)
);

OR2x6_ASAP7_75t_L g5705 ( 
.A(n_5270),
.B(n_5569),
.Y(n_5705)
);

OR2x6_ASAP7_75t_L g5706 ( 
.A(n_5270),
.B(n_5569),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5100),
.Y(n_5707)
);

AO31x2_ASAP7_75t_L g5708 ( 
.A1(n_5098),
.A2(n_4729),
.A3(n_5037),
.B(n_5077),
.Y(n_5708)
);

BUFx2_ASAP7_75t_L g5709 ( 
.A(n_5314),
.Y(n_5709)
);

BUFx6f_ASAP7_75t_L g5710 ( 
.A(n_5082),
.Y(n_5710)
);

NOR2xp33_ASAP7_75t_R g5711 ( 
.A(n_5158),
.B(n_4622),
.Y(n_5711)
);

INVx2_ASAP7_75t_L g5712 ( 
.A(n_5402),
.Y(n_5712)
);

BUFx4f_ASAP7_75t_SL g5713 ( 
.A(n_5258),
.Y(n_5713)
);

OAI22xp33_ASAP7_75t_L g5714 ( 
.A1(n_5121),
.A2(n_4989),
.B1(n_4979),
.B2(n_4944),
.Y(n_5714)
);

NOR2xp33_ASAP7_75t_R g5715 ( 
.A(n_5219),
.B(n_5367),
.Y(n_5715)
);

NAND2xp33_ASAP7_75t_R g5716 ( 
.A(n_5264),
.B(n_4979),
.Y(n_5716)
);

HB1xp67_ASAP7_75t_L g5717 ( 
.A(n_5237),
.Y(n_5717)
);

BUFx10_ASAP7_75t_L g5718 ( 
.A(n_5265),
.Y(n_5718)
);

BUFx2_ASAP7_75t_L g5719 ( 
.A(n_5314),
.Y(n_5719)
);

NAND2xp33_ASAP7_75t_SL g5720 ( 
.A(n_5129),
.B(n_4622),
.Y(n_5720)
);

CKINVDCx5p33_ASAP7_75t_R g5721 ( 
.A(n_5504),
.Y(n_5721)
);

AOI22xp33_ASAP7_75t_L g5722 ( 
.A1(n_5244),
.A2(n_4867),
.B1(n_4882),
.B2(n_4648),
.Y(n_5722)
);

BUFx2_ASAP7_75t_L g5723 ( 
.A(n_5314),
.Y(n_5723)
);

INVx3_ASAP7_75t_L g5724 ( 
.A(n_5323),
.Y(n_5724)
);

INVx1_ASAP7_75t_L g5725 ( 
.A(n_5107),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_5113),
.Y(n_5726)
);

AND2x4_ASAP7_75t_L g5727 ( 
.A(n_5215),
.B(n_4686),
.Y(n_5727)
);

NAND2xp5_ASAP7_75t_SL g5728 ( 
.A(n_5214),
.B(n_5056),
.Y(n_5728)
);

AND2x4_ASAP7_75t_L g5729 ( 
.A(n_5215),
.B(n_4686),
.Y(n_5729)
);

AOI22xp33_ASAP7_75t_L g5730 ( 
.A1(n_5369),
.A2(n_4867),
.B1(n_4882),
.B2(n_4648),
.Y(n_5730)
);

INVx2_ASAP7_75t_L g5731 ( 
.A(n_5223),
.Y(n_5731)
);

INVx2_ASAP7_75t_L g5732 ( 
.A(n_5223),
.Y(n_5732)
);

INVx2_ASAP7_75t_L g5733 ( 
.A(n_5246),
.Y(n_5733)
);

AO31x2_ASAP7_75t_L g5734 ( 
.A1(n_5098),
.A2(n_4729),
.A3(n_5080),
.B(n_5077),
.Y(n_5734)
);

INVxp67_ASAP7_75t_L g5735 ( 
.A(n_5597),
.Y(n_5735)
);

NOR3xp33_ASAP7_75t_SL g5736 ( 
.A(n_5504),
.B(n_5011),
.C(n_4926),
.Y(n_5736)
);

CKINVDCx20_ASAP7_75t_R g5737 ( 
.A(n_5346),
.Y(n_5737)
);

OAI22xp5_ASAP7_75t_L g5738 ( 
.A1(n_5209),
.A2(n_4960),
.B1(n_4817),
.B2(n_5011),
.Y(n_5738)
);

OR2x6_ASAP7_75t_L g5739 ( 
.A(n_5569),
.B(n_5064),
.Y(n_5739)
);

CKINVDCx5p33_ASAP7_75t_R g5740 ( 
.A(n_5604),
.Y(n_5740)
);

AO31x2_ASAP7_75t_L g5741 ( 
.A1(n_5102),
.A2(n_4729),
.A3(n_5080),
.B(n_5077),
.Y(n_5741)
);

INVx2_ASAP7_75t_L g5742 ( 
.A(n_5246),
.Y(n_5742)
);

CKINVDCx5p33_ASAP7_75t_R g5743 ( 
.A(n_5604),
.Y(n_5743)
);

NOR3xp33_ASAP7_75t_SL g5744 ( 
.A(n_5131),
.B(n_4842),
.C(n_4857),
.Y(n_5744)
);

NOR2xp33_ASAP7_75t_R g5745 ( 
.A(n_5500),
.B(n_4622),
.Y(n_5745)
);

NAND3xp33_ASAP7_75t_L g5746 ( 
.A(n_5360),
.B(n_5634),
.C(n_5339),
.Y(n_5746)
);

A2O1A1Ixp33_ASAP7_75t_L g5747 ( 
.A1(n_5119),
.A2(n_5040),
.B(n_4598),
.C(n_4645),
.Y(n_5747)
);

CKINVDCx5p33_ASAP7_75t_R g5748 ( 
.A(n_5387),
.Y(n_5748)
);

NAND2xp33_ASAP7_75t_R g5749 ( 
.A(n_5611),
.B(n_4979),
.Y(n_5749)
);

NAND2xp5_ASAP7_75t_SL g5750 ( 
.A(n_5104),
.B(n_5056),
.Y(n_5750)
);

CKINVDCx16_ASAP7_75t_R g5751 ( 
.A(n_5350),
.Y(n_5751)
);

NAND2xp5_ASAP7_75t_L g5752 ( 
.A(n_5092),
.B(n_4760),
.Y(n_5752)
);

INVx3_ASAP7_75t_L g5753 ( 
.A(n_5419),
.Y(n_5753)
);

INVx2_ASAP7_75t_L g5754 ( 
.A(n_5246),
.Y(n_5754)
);

NOR3xp33_ASAP7_75t_SL g5755 ( 
.A(n_5090),
.B(n_4842),
.C(n_4857),
.Y(n_5755)
);

OR2x6_ASAP7_75t_L g5756 ( 
.A(n_5569),
.B(n_5064),
.Y(n_5756)
);

AND2x4_ASAP7_75t_L g5757 ( 
.A(n_5215),
.B(n_4686),
.Y(n_5757)
);

INVxp33_ASAP7_75t_SL g5758 ( 
.A(n_5535),
.Y(n_5758)
);

INVx1_ASAP7_75t_L g5759 ( 
.A(n_5162),
.Y(n_5759)
);

AND2x2_ASAP7_75t_L g5760 ( 
.A(n_5145),
.B(n_4681),
.Y(n_5760)
);

NAND3xp33_ASAP7_75t_L g5761 ( 
.A(n_5634),
.B(n_5030),
.C(n_4747),
.Y(n_5761)
);

AND2x2_ASAP7_75t_L g5762 ( 
.A(n_5299),
.B(n_4681),
.Y(n_5762)
);

NOR3xp33_ASAP7_75t_SL g5763 ( 
.A(n_5213),
.B(n_5012),
.C(n_5059),
.Y(n_5763)
);

INVx2_ASAP7_75t_L g5764 ( 
.A(n_5246),
.Y(n_5764)
);

AND2x4_ASAP7_75t_L g5765 ( 
.A(n_5215),
.B(n_4686),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_5171),
.Y(n_5766)
);

INVx1_ASAP7_75t_SL g5767 ( 
.A(n_5350),
.Y(n_5767)
);

CKINVDCx5p33_ASAP7_75t_R g5768 ( 
.A(n_5387),
.Y(n_5768)
);

INVx2_ASAP7_75t_L g5769 ( 
.A(n_5246),
.Y(n_5769)
);

CKINVDCx20_ASAP7_75t_R g5770 ( 
.A(n_5500),
.Y(n_5770)
);

NAND2xp5_ASAP7_75t_L g5771 ( 
.A(n_5103),
.B(n_5316),
.Y(n_5771)
);

AND2x2_ASAP7_75t_L g5772 ( 
.A(n_5299),
.B(n_4681),
.Y(n_5772)
);

NAND2xp5_ASAP7_75t_L g5773 ( 
.A(n_5383),
.B(n_4760),
.Y(n_5773)
);

AO31x2_ASAP7_75t_L g5774 ( 
.A1(n_5102),
.A2(n_4729),
.A3(n_5080),
.B(n_5077),
.Y(n_5774)
);

INVx3_ASAP7_75t_L g5775 ( 
.A(n_5419),
.Y(n_5775)
);

HB1xp67_ASAP7_75t_L g5776 ( 
.A(n_5250),
.Y(n_5776)
);

AND2x2_ASAP7_75t_L g5777 ( 
.A(n_5302),
.B(n_4681),
.Y(n_5777)
);

NOR3xp33_ASAP7_75t_SL g5778 ( 
.A(n_5341),
.B(n_5012),
.C(n_5059),
.Y(n_5778)
);

INVx2_ASAP7_75t_L g5779 ( 
.A(n_5402),
.Y(n_5779)
);

BUFx2_ASAP7_75t_L g5780 ( 
.A(n_5500),
.Y(n_5780)
);

NOR3xp33_ASAP7_75t_SL g5781 ( 
.A(n_5393),
.B(n_4890),
.C(n_4919),
.Y(n_5781)
);

INVx2_ASAP7_75t_L g5782 ( 
.A(n_5402),
.Y(n_5782)
);

NOR2xp33_ASAP7_75t_R g5783 ( 
.A(n_5135),
.B(n_4681),
.Y(n_5783)
);

INVxp67_ASAP7_75t_SL g5784 ( 
.A(n_5086),
.Y(n_5784)
);

BUFx2_ASAP7_75t_L g5785 ( 
.A(n_5135),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5172),
.Y(n_5786)
);

OA21x2_ASAP7_75t_L g5787 ( 
.A1(n_5588),
.A2(n_4740),
.B(n_4733),
.Y(n_5787)
);

INVx2_ASAP7_75t_L g5788 ( 
.A(n_5167),
.Y(n_5788)
);

AOI22xp33_ASAP7_75t_L g5789 ( 
.A1(n_5182),
.A2(n_4867),
.B1(n_4882),
.B2(n_4819),
.Y(n_5789)
);

NAND2xp33_ASAP7_75t_R g5790 ( 
.A(n_5148),
.B(n_5163),
.Y(n_5790)
);

NAND2xp5_ASAP7_75t_L g5791 ( 
.A(n_5122),
.B(n_4766),
.Y(n_5791)
);

BUFx3_ASAP7_75t_L g5792 ( 
.A(n_5439),
.Y(n_5792)
);

AND2x4_ASAP7_75t_L g5793 ( 
.A(n_5252),
.B(n_4686),
.Y(n_5793)
);

NAND2xp5_ASAP7_75t_L g5794 ( 
.A(n_5124),
.B(n_4766),
.Y(n_5794)
);

BUFx5_ASAP7_75t_L g5795 ( 
.A(n_5454),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5186),
.Y(n_5796)
);

NOR2xp33_ASAP7_75t_R g5797 ( 
.A(n_5235),
.B(n_4707),
.Y(n_5797)
);

NOR3xp33_ASAP7_75t_SL g5798 ( 
.A(n_5393),
.B(n_4890),
.C(n_4707),
.Y(n_5798)
);

NAND2xp33_ASAP7_75t_R g5799 ( 
.A(n_5148),
.B(n_4989),
.Y(n_5799)
);

NOR2x1_ASAP7_75t_SL g5800 ( 
.A(n_5197),
.B(n_4960),
.Y(n_5800)
);

INVx3_ASAP7_75t_L g5801 ( 
.A(n_5089),
.Y(n_5801)
);

INVx3_ASAP7_75t_L g5802 ( 
.A(n_5089),
.Y(n_5802)
);

NAND2xp33_ASAP7_75t_R g5803 ( 
.A(n_5148),
.B(n_4989),
.Y(n_5803)
);

INVx1_ASAP7_75t_SL g5804 ( 
.A(n_5437),
.Y(n_5804)
);

CKINVDCx16_ASAP7_75t_R g5805 ( 
.A(n_5439),
.Y(n_5805)
);

INVxp67_ASAP7_75t_L g5806 ( 
.A(n_5087),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5263),
.Y(n_5807)
);

INVxp67_ASAP7_75t_L g5808 ( 
.A(n_5081),
.Y(n_5808)
);

NOR2xp33_ASAP7_75t_R g5809 ( 
.A(n_5235),
.B(n_4707),
.Y(n_5809)
);

AO31x2_ASAP7_75t_L g5810 ( 
.A1(n_5267),
.A2(n_5080),
.A3(n_4598),
.B(n_4645),
.Y(n_5810)
);

NOR2xp33_ASAP7_75t_L g5811 ( 
.A(n_5603),
.B(n_4707),
.Y(n_5811)
);

AND2x2_ASAP7_75t_L g5812 ( 
.A(n_5302),
.B(n_4707),
.Y(n_5812)
);

BUFx2_ASAP7_75t_L g5813 ( 
.A(n_5385),
.Y(n_5813)
);

AND2x2_ASAP7_75t_L g5814 ( 
.A(n_5356),
.B(n_5005),
.Y(n_5814)
);

HB1xp67_ASAP7_75t_L g5815 ( 
.A(n_5250),
.Y(n_5815)
);

AOI21xp5_ASAP7_75t_L g5816 ( 
.A1(n_5108),
.A2(n_4819),
.B(n_4951),
.Y(n_5816)
);

NAND2xp5_ASAP7_75t_L g5817 ( 
.A(n_5157),
.B(n_4898),
.Y(n_5817)
);

AND2x4_ASAP7_75t_L g5818 ( 
.A(n_5252),
.B(n_4712),
.Y(n_5818)
);

INVx4_ASAP7_75t_L g5819 ( 
.A(n_5265),
.Y(n_5819)
);

NOR3xp33_ASAP7_75t_SL g5820 ( 
.A(n_5459),
.B(n_5240),
.C(n_5311),
.Y(n_5820)
);

AOI22xp33_ASAP7_75t_L g5821 ( 
.A1(n_5182),
.A2(n_4819),
.B1(n_4591),
.B2(n_4602),
.Y(n_5821)
);

INVx2_ASAP7_75t_L g5822 ( 
.A(n_5306),
.Y(n_5822)
);

OAI21x1_ASAP7_75t_SL g5823 ( 
.A1(n_5587),
.A2(n_4966),
.B(n_5070),
.Y(n_5823)
);

CKINVDCx16_ASAP7_75t_R g5824 ( 
.A(n_5454),
.Y(n_5824)
);

NAND2xp5_ASAP7_75t_L g5825 ( 
.A(n_5180),
.B(n_4898),
.Y(n_5825)
);

NAND2xp5_ASAP7_75t_L g5826 ( 
.A(n_5190),
.B(n_4945),
.Y(n_5826)
);

OR2x2_ASAP7_75t_L g5827 ( 
.A(n_5190),
.B(n_4880),
.Y(n_5827)
);

INVx1_ASAP7_75t_L g5828 ( 
.A(n_5284),
.Y(n_5828)
);

BUFx2_ASAP7_75t_L g5829 ( 
.A(n_5385),
.Y(n_5829)
);

INVx2_ASAP7_75t_L g5830 ( 
.A(n_5306),
.Y(n_5830)
);

CKINVDCx5p33_ASAP7_75t_R g5831 ( 
.A(n_5509),
.Y(n_5831)
);

HB1xp67_ASAP7_75t_L g5832 ( 
.A(n_5342),
.Y(n_5832)
);

OR2x6_ASAP7_75t_L g5833 ( 
.A(n_5436),
.B(n_5064),
.Y(n_5833)
);

AND2x2_ASAP7_75t_L g5834 ( 
.A(n_5356),
.B(n_5005),
.Y(n_5834)
);

HB1xp67_ASAP7_75t_L g5835 ( 
.A(n_5342),
.Y(n_5835)
);

NOR2xp33_ASAP7_75t_R g5836 ( 
.A(n_5509),
.B(n_5005),
.Y(n_5836)
);

CKINVDCx16_ASAP7_75t_R g5837 ( 
.A(n_5436),
.Y(n_5837)
);

INVx2_ASAP7_75t_L g5838 ( 
.A(n_5306),
.Y(n_5838)
);

AND2x4_ASAP7_75t_L g5839 ( 
.A(n_5252),
.B(n_4712),
.Y(n_5839)
);

OAI22xp5_ASAP7_75t_L g5840 ( 
.A1(n_5200),
.A2(n_4960),
.B1(n_4673),
.B2(n_4987),
.Y(n_5840)
);

HB1xp67_ASAP7_75t_L g5841 ( 
.A(n_5347),
.Y(n_5841)
);

AND2x2_ASAP7_75t_L g5842 ( 
.A(n_5391),
.B(n_5005),
.Y(n_5842)
);

OAI21xp5_ASAP7_75t_L g5843 ( 
.A1(n_5196),
.A2(n_4910),
.B(n_4645),
.Y(n_5843)
);

NOR3xp33_ASAP7_75t_SL g5844 ( 
.A(n_5311),
.B(n_5005),
.C(n_5009),
.Y(n_5844)
);

AOI22xp33_ASAP7_75t_L g5845 ( 
.A1(n_5182),
.A2(n_4819),
.B1(n_4591),
.B2(n_4602),
.Y(n_5845)
);

INVx1_ASAP7_75t_L g5846 ( 
.A(n_5290),
.Y(n_5846)
);

INVx3_ASAP7_75t_L g5847 ( 
.A(n_5089),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_5292),
.Y(n_5848)
);

OAI22xp5_ASAP7_75t_L g5849 ( 
.A1(n_5156),
.A2(n_5212),
.B1(n_5151),
.B2(n_5388),
.Y(n_5849)
);

OR2x6_ASAP7_75t_L g5850 ( 
.A(n_5436),
.B(n_5064),
.Y(n_5850)
);

NOR3xp33_ASAP7_75t_SL g5851 ( 
.A(n_5132),
.B(n_5283),
.C(n_5261),
.Y(n_5851)
);

AOI22xp33_ASAP7_75t_L g5852 ( 
.A1(n_5201),
.A2(n_4819),
.B1(n_4591),
.B2(n_4602),
.Y(n_5852)
);

AND2x2_ASAP7_75t_L g5853 ( 
.A(n_5391),
.B(n_4914),
.Y(n_5853)
);

HB1xp67_ASAP7_75t_L g5854 ( 
.A(n_5347),
.Y(n_5854)
);

NAND2xp33_ASAP7_75t_R g5855 ( 
.A(n_5163),
.B(n_4989),
.Y(n_5855)
);

OR2x2_ASAP7_75t_L g5856 ( 
.A(n_5236),
.B(n_5170),
.Y(n_5856)
);

NOR2xp33_ASAP7_75t_L g5857 ( 
.A(n_5603),
.B(n_4945),
.Y(n_5857)
);

INVxp67_ASAP7_75t_L g5858 ( 
.A(n_5133),
.Y(n_5858)
);

NAND3xp33_ASAP7_75t_SL g5859 ( 
.A(n_5153),
.B(n_4823),
.C(n_4897),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_5295),
.Y(n_5860)
);

INVx2_ASAP7_75t_L g5861 ( 
.A(n_5167),
.Y(n_5861)
);

NAND2xp33_ASAP7_75t_R g5862 ( 
.A(n_5163),
.B(n_4989),
.Y(n_5862)
);

CKINVDCx11_ASAP7_75t_R g5863 ( 
.A(n_5603),
.Y(n_5863)
);

NAND3xp33_ASAP7_75t_SL g5864 ( 
.A(n_5205),
.B(n_5629),
.C(n_5156),
.Y(n_5864)
);

CKINVDCx5p33_ASAP7_75t_R g5865 ( 
.A(n_5551),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5298),
.Y(n_5866)
);

NOR2xp33_ASAP7_75t_R g5867 ( 
.A(n_5265),
.B(n_5045),
.Y(n_5867)
);

CKINVDCx16_ASAP7_75t_R g5868 ( 
.A(n_5265),
.Y(n_5868)
);

INVx3_ASAP7_75t_L g5869 ( 
.A(n_5111),
.Y(n_5869)
);

OAI21xp5_ASAP7_75t_L g5870 ( 
.A1(n_5108),
.A2(n_4910),
.B(n_4649),
.Y(n_5870)
);

NOR2xp33_ASAP7_75t_L g5871 ( 
.A(n_5551),
.B(n_4712),
.Y(n_5871)
);

INVx2_ASAP7_75t_L g5872 ( 
.A(n_5249),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5307),
.Y(n_5873)
);

OR2x6_ASAP7_75t_L g5874 ( 
.A(n_5636),
.B(n_4666),
.Y(n_5874)
);

NAND2xp5_ASAP7_75t_L g5875 ( 
.A(n_5236),
.B(n_4688),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_5309),
.Y(n_5876)
);

OR2x2_ASAP7_75t_L g5877 ( 
.A(n_5170),
.B(n_4909),
.Y(n_5877)
);

NAND3xp33_ASAP7_75t_SL g5878 ( 
.A(n_5188),
.B(n_4823),
.C(n_4897),
.Y(n_5878)
);

CKINVDCx5p33_ASAP7_75t_R g5879 ( 
.A(n_5551),
.Y(n_5879)
);

AND2x2_ASAP7_75t_L g5880 ( 
.A(n_5462),
.B(n_4914),
.Y(n_5880)
);

CKINVDCx5p33_ASAP7_75t_R g5881 ( 
.A(n_5484),
.Y(n_5881)
);

AO31x2_ASAP7_75t_L g5882 ( 
.A1(n_5267),
.A2(n_4599),
.A3(n_4670),
.B(n_4649),
.Y(n_5882)
);

BUFx3_ASAP7_75t_L g5883 ( 
.A(n_5265),
.Y(n_5883)
);

O2A1O1Ixp33_ASAP7_75t_SL g5884 ( 
.A1(n_5548),
.A2(n_4689),
.B(n_4732),
.C(n_4688),
.Y(n_5884)
);

NOR3xp33_ASAP7_75t_SL g5885 ( 
.A(n_5275),
.B(n_5254),
.C(n_5101),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5313),
.Y(n_5886)
);

CKINVDCx5p33_ASAP7_75t_R g5887 ( 
.A(n_5484),
.Y(n_5887)
);

NOR3xp33_ASAP7_75t_SL g5888 ( 
.A(n_5481),
.B(n_5027),
.C(n_5009),
.Y(n_5888)
);

INVx2_ASAP7_75t_L g5889 ( 
.A(n_5249),
.Y(n_5889)
);

AND2x2_ASAP7_75t_L g5890 ( 
.A(n_5462),
.B(n_4914),
.Y(n_5890)
);

NAND2xp5_ASAP7_75t_L g5891 ( 
.A(n_5232),
.B(n_4689),
.Y(n_5891)
);

NAND2xp5_ASAP7_75t_L g5892 ( 
.A(n_5234),
.B(n_4732),
.Y(n_5892)
);

AND2x2_ASAP7_75t_L g5893 ( 
.A(n_5252),
.B(n_4873),
.Y(n_5893)
);

INVx2_ASAP7_75t_L g5894 ( 
.A(n_5324),
.Y(n_5894)
);

CKINVDCx5p33_ASAP7_75t_R g5895 ( 
.A(n_5484),
.Y(n_5895)
);

AND2x4_ASAP7_75t_L g5896 ( 
.A(n_5259),
.B(n_4712),
.Y(n_5896)
);

AOI22xp33_ASAP7_75t_SL g5897 ( 
.A1(n_5434),
.A2(n_5030),
.B1(n_4670),
.B2(n_4649),
.Y(n_5897)
);

AOI22xp33_ASAP7_75t_L g5898 ( 
.A1(n_5201),
.A2(n_4591),
.B1(n_4602),
.B2(n_4670),
.Y(n_5898)
);

HB1xp67_ASAP7_75t_L g5899 ( 
.A(n_5351),
.Y(n_5899)
);

NOR2xp33_ASAP7_75t_R g5900 ( 
.A(n_5105),
.B(n_5045),
.Y(n_5900)
);

AND2x2_ASAP7_75t_L g5901 ( 
.A(n_5259),
.B(n_4873),
.Y(n_5901)
);

AO31x2_ASAP7_75t_L g5902 ( 
.A1(n_5321),
.A2(n_5492),
.A3(n_5374),
.B(n_5469),
.Y(n_5902)
);

INVx2_ASAP7_75t_L g5903 ( 
.A(n_5324),
.Y(n_5903)
);

AOI22xp33_ASAP7_75t_L g5904 ( 
.A1(n_5201),
.A2(n_4591),
.B1(n_4602),
.B2(n_4621),
.Y(n_5904)
);

NAND2xp5_ASAP7_75t_L g5905 ( 
.A(n_5114),
.B(n_4750),
.Y(n_5905)
);

AO31x2_ASAP7_75t_L g5906 ( 
.A1(n_5321),
.A2(n_5054),
.A3(n_5057),
.B(n_5046),
.Y(n_5906)
);

OAI22xp5_ASAP7_75t_L g5907 ( 
.A1(n_5192),
.A2(n_4960),
.B1(n_4987),
.B2(n_5062),
.Y(n_5907)
);

BUFx8_ASAP7_75t_SL g5908 ( 
.A(n_5373),
.Y(n_5908)
);

OR2x6_ASAP7_75t_L g5909 ( 
.A(n_5636),
.B(n_4666),
.Y(n_5909)
);

AND2x2_ASAP7_75t_L g5910 ( 
.A(n_5259),
.B(n_4873),
.Y(n_5910)
);

BUFx6f_ASAP7_75t_L g5911 ( 
.A(n_5489),
.Y(n_5911)
);

AND2x2_ASAP7_75t_L g5912 ( 
.A(n_5259),
.B(n_4856),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_5320),
.Y(n_5913)
);

INVx2_ASAP7_75t_L g5914 ( 
.A(n_5286),
.Y(n_5914)
);

AND2x2_ASAP7_75t_L g5915 ( 
.A(n_5637),
.B(n_4856),
.Y(n_5915)
);

INVx2_ASAP7_75t_L g5916 ( 
.A(n_5286),
.Y(n_5916)
);

AND2x2_ASAP7_75t_L g5917 ( 
.A(n_5637),
.B(n_4856),
.Y(n_5917)
);

AOI22xp33_ASAP7_75t_SL g5918 ( 
.A1(n_5447),
.A2(n_5471),
.B1(n_5518),
.B2(n_5030),
.Y(n_5918)
);

CKINVDCx16_ASAP7_75t_R g5919 ( 
.A(n_5105),
.Y(n_5919)
);

INVx1_ASAP7_75t_L g5920 ( 
.A(n_5325),
.Y(n_5920)
);

AND2x2_ASAP7_75t_L g5921 ( 
.A(n_5105),
.B(n_4930),
.Y(n_5921)
);

OAI21xp5_ASAP7_75t_SL g5922 ( 
.A1(n_5136),
.A2(n_5062),
.B(n_4987),
.Y(n_5922)
);

NOR2xp33_ASAP7_75t_L g5923 ( 
.A(n_5115),
.B(n_4712),
.Y(n_5923)
);

INVx2_ASAP7_75t_L g5924 ( 
.A(n_5286),
.Y(n_5924)
);

NOR3xp33_ASAP7_75t_SL g5925 ( 
.A(n_5487),
.B(n_5042),
.C(n_5027),
.Y(n_5925)
);

NOR2xp33_ASAP7_75t_L g5926 ( 
.A(n_5638),
.B(n_4745),
.Y(n_5926)
);

AND2x2_ASAP7_75t_L g5927 ( 
.A(n_5280),
.B(n_4930),
.Y(n_5927)
);

CKINVDCx5p33_ASAP7_75t_R g5928 ( 
.A(n_5505),
.Y(n_5928)
);

BUFx6f_ASAP7_75t_L g5929 ( 
.A(n_5489),
.Y(n_5929)
);

AO31x2_ASAP7_75t_L g5930 ( 
.A1(n_5374),
.A2(n_5054),
.A3(n_5057),
.B(n_5046),
.Y(n_5930)
);

AND2x6_ASAP7_75t_L g5931 ( 
.A(n_5489),
.B(n_4762),
.Y(n_5931)
);

OR2x6_ASAP7_75t_L g5932 ( 
.A(n_5303),
.B(n_4666),
.Y(n_5932)
);

HB1xp67_ASAP7_75t_L g5933 ( 
.A(n_5351),
.Y(n_5933)
);

AND2x2_ASAP7_75t_L g5934 ( 
.A(n_5280),
.B(n_5319),
.Y(n_5934)
);

AO31x2_ASAP7_75t_L g5935 ( 
.A1(n_5492),
.A2(n_5054),
.A3(n_5057),
.B(n_5046),
.Y(n_5935)
);

OR2x2_ASAP7_75t_L g5936 ( 
.A(n_5085),
.B(n_4909),
.Y(n_5936)
);

OR2x2_ASAP7_75t_L g5937 ( 
.A(n_5085),
.B(n_4921),
.Y(n_5937)
);

INVx1_ASAP7_75t_SL g5938 ( 
.A(n_5505),
.Y(n_5938)
);

INVx2_ASAP7_75t_L g5939 ( 
.A(n_5286),
.Y(n_5939)
);

NOR2xp33_ASAP7_75t_L g5940 ( 
.A(n_5129),
.B(n_4745),
.Y(n_5940)
);

NOR2xp33_ASAP7_75t_L g5941 ( 
.A(n_5247),
.B(n_4745),
.Y(n_5941)
);

AND2x2_ASAP7_75t_L g5942 ( 
.A(n_5280),
.B(n_4930),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_5329),
.Y(n_5943)
);

INVx1_ASAP7_75t_L g5944 ( 
.A(n_5330),
.Y(n_5944)
);

NAND2xp5_ASAP7_75t_L g5945 ( 
.A(n_5357),
.B(n_4750),
.Y(n_5945)
);

NOR2xp67_ASAP7_75t_L g5946 ( 
.A(n_5211),
.B(n_4825),
.Y(n_5946)
);

NOR3xp33_ASAP7_75t_SL g5947 ( 
.A(n_5229),
.B(n_5042),
.C(n_4916),
.Y(n_5947)
);

CKINVDCx5p33_ASAP7_75t_R g5948 ( 
.A(n_5505),
.Y(n_5948)
);

AND2x2_ASAP7_75t_L g5949 ( 
.A(n_5319),
.B(n_4930),
.Y(n_5949)
);

AND2x2_ASAP7_75t_L g5950 ( 
.A(n_5319),
.B(n_4930),
.Y(n_5950)
);

NOR2xp33_ASAP7_75t_R g5951 ( 
.A(n_5505),
.B(n_5045),
.Y(n_5951)
);

AND2x2_ASAP7_75t_L g5952 ( 
.A(n_5111),
.B(n_4975),
.Y(n_5952)
);

NOR2x1p5_ASAP7_75t_L g5953 ( 
.A(n_5111),
.B(n_5143),
.Y(n_5953)
);

INVx3_ASAP7_75t_L g5954 ( 
.A(n_5143),
.Y(n_5954)
);

AOI22xp33_ASAP7_75t_L g5955 ( 
.A1(n_5202),
.A2(n_4621),
.B1(n_4758),
.B2(n_4610),
.Y(n_5955)
);

NAND3xp33_ASAP7_75t_SL g5956 ( 
.A(n_5188),
.B(n_4897),
.C(n_4885),
.Y(n_5956)
);

INVx2_ASAP7_75t_L g5957 ( 
.A(n_5269),
.Y(n_5957)
);

AND2x2_ASAP7_75t_L g5958 ( 
.A(n_5143),
.B(n_4975),
.Y(n_5958)
);

AO31x2_ASAP7_75t_L g5959 ( 
.A1(n_5465),
.A2(n_5054),
.A3(n_5057),
.B(n_5046),
.Y(n_5959)
);

CKINVDCx5p33_ASAP7_75t_R g5960 ( 
.A(n_5511),
.Y(n_5960)
);

INVx1_ASAP7_75t_L g5961 ( 
.A(n_5332),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5335),
.Y(n_5962)
);

OR2x6_ASAP7_75t_L g5963 ( 
.A(n_5303),
.B(n_4666),
.Y(n_5963)
);

CKINVDCx5p33_ASAP7_75t_R g5964 ( 
.A(n_5607),
.Y(n_5964)
);

CKINVDCx12_ASAP7_75t_R g5965 ( 
.A(n_5373),
.Y(n_5965)
);

INVx1_ASAP7_75t_L g5966 ( 
.A(n_5336),
.Y(n_5966)
);

AND2x2_ASAP7_75t_L g5967 ( 
.A(n_5179),
.B(n_4975),
.Y(n_5967)
);

INVx3_ASAP7_75t_L g5968 ( 
.A(n_5179),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_5358),
.Y(n_5969)
);

AND2x2_ASAP7_75t_L g5970 ( 
.A(n_5179),
.B(n_4975),
.Y(n_5970)
);

AOI22xp33_ASAP7_75t_L g5971 ( 
.A1(n_5202),
.A2(n_4621),
.B1(n_4758),
.B2(n_4610),
.Y(n_5971)
);

OR2x6_ASAP7_75t_L g5972 ( 
.A(n_5303),
.B(n_4666),
.Y(n_5972)
);

OR2x6_ASAP7_75t_L g5973 ( 
.A(n_5414),
.B(n_4666),
.Y(n_5973)
);

HB1xp67_ASAP7_75t_L g5974 ( 
.A(n_5421),
.Y(n_5974)
);

BUFx3_ASAP7_75t_L g5975 ( 
.A(n_5489),
.Y(n_5975)
);

OAI21xp5_ASAP7_75t_L g5976 ( 
.A1(n_5191),
.A2(n_4885),
.B(n_4951),
.Y(n_5976)
);

AND2x4_ASAP7_75t_L g5977 ( 
.A(n_5273),
.B(n_4745),
.Y(n_5977)
);

INVx1_ASAP7_75t_SL g5978 ( 
.A(n_5217),
.Y(n_5978)
);

BUFx2_ASAP7_75t_L g5979 ( 
.A(n_5139),
.Y(n_5979)
);

CKINVDCx5p33_ASAP7_75t_R g5980 ( 
.A(n_5146),
.Y(n_5980)
);

INVx1_ASAP7_75t_L g5981 ( 
.A(n_5370),
.Y(n_5981)
);

INVxp67_ASAP7_75t_L g5982 ( 
.A(n_5149),
.Y(n_5982)
);

AND2x4_ASAP7_75t_L g5983 ( 
.A(n_5273),
.B(n_4745),
.Y(n_5983)
);

CKINVDCx16_ASAP7_75t_R g5984 ( 
.A(n_5373),
.Y(n_5984)
);

AND2x2_ASAP7_75t_L g5985 ( 
.A(n_5273),
.B(n_4975),
.Y(n_5985)
);

INVx2_ASAP7_75t_L g5986 ( 
.A(n_5269),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5371),
.Y(n_5987)
);

OAI21xp5_ASAP7_75t_L g5988 ( 
.A1(n_5191),
.A2(n_4885),
.B(n_4844),
.Y(n_5988)
);

AND2x4_ASAP7_75t_L g5989 ( 
.A(n_5587),
.B(n_4763),
.Y(n_5989)
);

NOR2x1_ASAP7_75t_L g5990 ( 
.A(n_5199),
.B(n_5045),
.Y(n_5990)
);

AO21x2_ASAP7_75t_L g5991 ( 
.A1(n_5526),
.A2(n_4626),
.B(n_4621),
.Y(n_5991)
);

NOR2xp33_ASAP7_75t_L g5992 ( 
.A(n_5331),
.B(n_4763),
.Y(n_5992)
);

NOR2xp33_ASAP7_75t_R g5993 ( 
.A(n_5495),
.B(n_5045),
.Y(n_5993)
);

AND2x2_ASAP7_75t_L g5994 ( 
.A(n_5571),
.B(n_5035),
.Y(n_5994)
);

AND2x4_ASAP7_75t_L g5995 ( 
.A(n_5495),
.B(n_4763),
.Y(n_5995)
);

OR2x2_ASAP7_75t_L g5996 ( 
.A(n_5159),
.B(n_4921),
.Y(n_5996)
);

INVx1_ASAP7_75t_L g5997 ( 
.A(n_5379),
.Y(n_5997)
);

AND2x2_ASAP7_75t_L g5998 ( 
.A(n_5571),
.B(n_5035),
.Y(n_5998)
);

OR2x6_ASAP7_75t_L g5999 ( 
.A(n_5414),
.B(n_4677),
.Y(n_5999)
);

NOR2xp33_ASAP7_75t_R g6000 ( 
.A(n_5495),
.B(n_5024),
.Y(n_6000)
);

NAND2xp5_ASAP7_75t_L g6001 ( 
.A(n_5243),
.B(n_4754),
.Y(n_6001)
);

OAI21xp5_ASAP7_75t_SL g6002 ( 
.A1(n_5239),
.A2(n_5062),
.B(n_4987),
.Y(n_6002)
);

AO31x2_ASAP7_75t_L g6003 ( 
.A1(n_5440),
.A2(n_5069),
.A3(n_5066),
.B(n_4757),
.Y(n_6003)
);

OR2x2_ASAP7_75t_L g6004 ( 
.A(n_5159),
.B(n_4777),
.Y(n_6004)
);

OR2x2_ASAP7_75t_L g6005 ( 
.A(n_5221),
.B(n_4777),
.Y(n_6005)
);

OR2x2_ASAP7_75t_L g6006 ( 
.A(n_5242),
.B(n_4777),
.Y(n_6006)
);

CKINVDCx16_ASAP7_75t_R g6007 ( 
.A(n_5373),
.Y(n_6007)
);

CKINVDCx5p33_ASAP7_75t_R g6008 ( 
.A(n_5168),
.Y(n_6008)
);

BUFx3_ASAP7_75t_L g6009 ( 
.A(n_5489),
.Y(n_6009)
);

BUFx3_ASAP7_75t_L g6010 ( 
.A(n_5495),
.Y(n_6010)
);

AND2x2_ASAP7_75t_L g6011 ( 
.A(n_5584),
.B(n_5035),
.Y(n_6011)
);

INVx2_ASAP7_75t_L g6012 ( 
.A(n_5096),
.Y(n_6012)
);

INVx1_ASAP7_75t_L g6013 ( 
.A(n_5398),
.Y(n_6013)
);

CKINVDCx11_ASAP7_75t_R g6014 ( 
.A(n_5573),
.Y(n_6014)
);

NOR2x1_ASAP7_75t_SL g6015 ( 
.A(n_5197),
.B(n_4960),
.Y(n_6015)
);

AND2x4_ASAP7_75t_L g6016 ( 
.A(n_5495),
.B(n_4763),
.Y(n_6016)
);

AND2x2_ASAP7_75t_L g6017 ( 
.A(n_5584),
.B(n_5035),
.Y(n_6017)
);

AND2x2_ASAP7_75t_L g6018 ( 
.A(n_5612),
.B(n_5630),
.Y(n_6018)
);

AND2x4_ASAP7_75t_L g6019 ( 
.A(n_5560),
.B(n_4763),
.Y(n_6019)
);

BUFx3_ASAP7_75t_L g6020 ( 
.A(n_5208),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5409),
.Y(n_6021)
);

AND2x4_ASAP7_75t_L g6022 ( 
.A(n_5560),
.B(n_4806),
.Y(n_6022)
);

NAND2xp5_ASAP7_75t_L g6023 ( 
.A(n_5274),
.B(n_4754),
.Y(n_6023)
);

NAND2xp5_ASAP7_75t_L g6024 ( 
.A(n_5331),
.B(n_4761),
.Y(n_6024)
);

AND2x2_ASAP7_75t_L g6025 ( 
.A(n_5612),
.B(n_5035),
.Y(n_6025)
);

NAND3x1_ASAP7_75t_L g6026 ( 
.A(n_5147),
.B(n_4659),
.C(n_4588),
.Y(n_6026)
);

CKINVDCx20_ASAP7_75t_R g6027 ( 
.A(n_5294),
.Y(n_6027)
);

INVx1_ASAP7_75t_L g6028 ( 
.A(n_5472),
.Y(n_6028)
);

CKINVDCx5p33_ASAP7_75t_R g6029 ( 
.A(n_5224),
.Y(n_6029)
);

AND2x2_ASAP7_75t_L g6030 ( 
.A(n_5630),
.B(n_4806),
.Y(n_6030)
);

CKINVDCx20_ASAP7_75t_R g6031 ( 
.A(n_5127),
.Y(n_6031)
);

AOI22xp33_ASAP7_75t_L g6032 ( 
.A1(n_5202),
.A2(n_4621),
.B1(n_4758),
.B2(n_4610),
.Y(n_6032)
);

AND2x2_ASAP7_75t_L g6033 ( 
.A(n_5494),
.B(n_4806),
.Y(n_6033)
);

AOI22xp33_ASAP7_75t_L g6034 ( 
.A1(n_5174),
.A2(n_4758),
.B1(n_4610),
.B2(n_4611),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5475),
.Y(n_6035)
);

INVx2_ASAP7_75t_L g6036 ( 
.A(n_5096),
.Y(n_6036)
);

NAND2x1p5_ASAP7_75t_L g6037 ( 
.A(n_5536),
.B(n_5056),
.Y(n_6037)
);

AOI22xp33_ASAP7_75t_SL g6038 ( 
.A1(n_5447),
.A2(n_4991),
.B1(n_5044),
.B2(n_5038),
.Y(n_6038)
);

INVx1_ASAP7_75t_L g6039 ( 
.A(n_5478),
.Y(n_6039)
);

CKINVDCx16_ASAP7_75t_R g6040 ( 
.A(n_5308),
.Y(n_6040)
);

AND2x2_ASAP7_75t_L g6041 ( 
.A(n_5494),
.B(n_4806),
.Y(n_6041)
);

NAND2xp5_ASAP7_75t_L g6042 ( 
.A(n_5242),
.B(n_4761),
.Y(n_6042)
);

INVx1_ASAP7_75t_L g6043 ( 
.A(n_5483),
.Y(n_6043)
);

CKINVDCx16_ASAP7_75t_R g6044 ( 
.A(n_5333),
.Y(n_6044)
);

INVx2_ASAP7_75t_L g6045 ( 
.A(n_5096),
.Y(n_6045)
);

OAI21xp5_ASAP7_75t_L g6046 ( 
.A1(n_5440),
.A2(n_4844),
.B(n_4631),
.Y(n_6046)
);

NAND2xp5_ASAP7_75t_SL g6047 ( 
.A(n_5463),
.B(n_5414),
.Y(n_6047)
);

INVx2_ASAP7_75t_L g6048 ( 
.A(n_5206),
.Y(n_6048)
);

AND2x2_ASAP7_75t_L g6049 ( 
.A(n_5531),
.B(n_4806),
.Y(n_6049)
);

BUFx8_ASAP7_75t_L g6050 ( 
.A(n_5531),
.Y(n_6050)
);

INVx2_ASAP7_75t_L g6051 ( 
.A(n_5518),
.Y(n_6051)
);

NAND2xp5_ASAP7_75t_L g6052 ( 
.A(n_5245),
.B(n_4797),
.Y(n_6052)
);

AOI22xp5_ASAP7_75t_L g6053 ( 
.A1(n_5093),
.A2(n_4991),
.B1(n_4934),
.B2(n_5038),
.Y(n_6053)
);

NOR3xp33_ASAP7_75t_SL g6054 ( 
.A(n_5389),
.B(n_4916),
.C(n_4718),
.Y(n_6054)
);

AND2x2_ASAP7_75t_SL g6055 ( 
.A(n_5518),
.B(n_4762),
.Y(n_6055)
);

NOR2xp33_ASAP7_75t_L g6056 ( 
.A(n_5245),
.B(n_4846),
.Y(n_6056)
);

AND2x4_ASAP7_75t_L g6057 ( 
.A(n_5560),
.B(n_4846),
.Y(n_6057)
);

AND2x2_ASAP7_75t_L g6058 ( 
.A(n_5349),
.B(n_4846),
.Y(n_6058)
);

AND2x2_ASAP7_75t_L g6059 ( 
.A(n_5349),
.B(n_4846),
.Y(n_6059)
);

AND2x6_ASAP7_75t_L g6060 ( 
.A(n_5601),
.B(n_4762),
.Y(n_6060)
);

CKINVDCx16_ASAP7_75t_R g6061 ( 
.A(n_5333),
.Y(n_6061)
);

A2O1A1Ixp33_ASAP7_75t_L g6062 ( 
.A1(n_5453),
.A2(n_4580),
.B(n_4884),
.C(n_4827),
.Y(n_6062)
);

AO31x2_ASAP7_75t_L g6063 ( 
.A1(n_5453),
.A2(n_5069),
.A3(n_5066),
.B(n_4757),
.Y(n_6063)
);

INVx2_ASAP7_75t_L g6064 ( 
.A(n_5206),
.Y(n_6064)
);

AND2x4_ASAP7_75t_L g6065 ( 
.A(n_5279),
.B(n_4846),
.Y(n_6065)
);

INVx3_ASAP7_75t_L g6066 ( 
.A(n_5416),
.Y(n_6066)
);

NAND2xp5_ASAP7_75t_L g6067 ( 
.A(n_5615),
.B(n_4797),
.Y(n_6067)
);

AND2x2_ASAP7_75t_L g6068 ( 
.A(n_5353),
.B(n_5021),
.Y(n_6068)
);

BUFx2_ASAP7_75t_L g6069 ( 
.A(n_5197),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_5206),
.Y(n_6070)
);

CKINVDCx16_ASAP7_75t_R g6071 ( 
.A(n_5333),
.Y(n_6071)
);

CKINVDCx5p33_ASAP7_75t_R g6072 ( 
.A(n_5226),
.Y(n_6072)
);

NAND2xp33_ASAP7_75t_R g6073 ( 
.A(n_5174),
.B(n_4986),
.Y(n_6073)
);

INVx2_ASAP7_75t_L g6074 ( 
.A(n_5206),
.Y(n_6074)
);

BUFx6f_ASAP7_75t_L g6075 ( 
.A(n_5446),
.Y(n_6075)
);

OAI22xp33_ASAP7_75t_L g6076 ( 
.A1(n_5628),
.A2(n_5632),
.B1(n_5413),
.B2(n_5266),
.Y(n_6076)
);

AND2x2_ASAP7_75t_L g6077 ( 
.A(n_5353),
.B(n_5021),
.Y(n_6077)
);

XNOR2x1_ASAP7_75t_L g6078 ( 
.A(n_5403),
.B(n_4825),
.Y(n_6078)
);

NAND2xp33_ASAP7_75t_SL g6079 ( 
.A(n_5097),
.B(n_4812),
.Y(n_6079)
);

AOI22xp5_ASAP7_75t_L g6080 ( 
.A1(n_5590),
.A2(n_4991),
.B1(n_4934),
.B2(n_5044),
.Y(n_6080)
);

NAND2xp5_ASAP7_75t_L g6081 ( 
.A(n_5288),
.B(n_4812),
.Y(n_6081)
);

INVx2_ASAP7_75t_SL g6082 ( 
.A(n_5405),
.Y(n_6082)
);

NAND3xp33_ASAP7_75t_SL g6083 ( 
.A(n_5094),
.B(n_5062),
.C(n_4974),
.Y(n_6083)
);

NOR2xp33_ASAP7_75t_R g6084 ( 
.A(n_5372),
.B(n_5056),
.Y(n_6084)
);

NAND2xp5_ASAP7_75t_L g6085 ( 
.A(n_5359),
.B(n_4829),
.Y(n_6085)
);

AND2x2_ASAP7_75t_L g6086 ( 
.A(n_5368),
.B(n_5021),
.Y(n_6086)
);

NAND2xp5_ASAP7_75t_L g6087 ( 
.A(n_5364),
.B(n_4829),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_5488),
.Y(n_6088)
);

NOR2xp33_ASAP7_75t_R g6089 ( 
.A(n_5372),
.B(n_4762),
.Y(n_6089)
);

NOR2x1p5_ASAP7_75t_L g6090 ( 
.A(n_5570),
.B(n_4827),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_5491),
.Y(n_6091)
);

AND2x4_ASAP7_75t_L g6092 ( 
.A(n_5279),
.B(n_4825),
.Y(n_6092)
);

NOR3xp33_ASAP7_75t_SL g6093 ( 
.A(n_5268),
.B(n_4718),
.C(n_4706),
.Y(n_6093)
);

NAND2xp5_ASAP7_75t_L g6094 ( 
.A(n_5318),
.B(n_4871),
.Y(n_6094)
);

BUFx2_ASAP7_75t_L g6095 ( 
.A(n_5197),
.Y(n_6095)
);

CKINVDCx16_ASAP7_75t_R g6096 ( 
.A(n_5333),
.Y(n_6096)
);

AND2x2_ASAP7_75t_L g6097 ( 
.A(n_5368),
.B(n_5021),
.Y(n_6097)
);

INVx3_ASAP7_75t_L g6098 ( 
.A(n_5416),
.Y(n_6098)
);

BUFx3_ASAP7_75t_L g6099 ( 
.A(n_5443),
.Y(n_6099)
);

BUFx2_ASAP7_75t_L g6100 ( 
.A(n_5508),
.Y(n_6100)
);

AO31x2_ASAP7_75t_L g6101 ( 
.A1(n_5540),
.A2(n_5069),
.A3(n_5066),
.B(n_4757),
.Y(n_6101)
);

OAI21xp5_ASAP7_75t_L g6102 ( 
.A1(n_5272),
.A2(n_4844),
.B(n_4631),
.Y(n_6102)
);

INVx1_ASAP7_75t_SL g6103 ( 
.A(n_5318),
.Y(n_6103)
);

NOR2xp33_ASAP7_75t_L g6104 ( 
.A(n_5400),
.B(n_4871),
.Y(n_6104)
);

HB1xp67_ASAP7_75t_L g6105 ( 
.A(n_5421),
.Y(n_6105)
);

BUFx3_ASAP7_75t_L g6106 ( 
.A(n_5446),
.Y(n_6106)
);

NAND2xp5_ASAP7_75t_L g6107 ( 
.A(n_5343),
.B(n_4911),
.Y(n_6107)
);

NAND2xp5_ASAP7_75t_L g6108 ( 
.A(n_5530),
.B(n_4911),
.Y(n_6108)
);

INVx3_ASAP7_75t_L g6109 ( 
.A(n_5416),
.Y(n_6109)
);

AND2x2_ASAP7_75t_L g6110 ( 
.A(n_5544),
.B(n_5021),
.Y(n_6110)
);

BUFx2_ASAP7_75t_L g6111 ( 
.A(n_5416),
.Y(n_6111)
);

CKINVDCx5p33_ASAP7_75t_R g6112 ( 
.A(n_5446),
.Y(n_6112)
);

CKINVDCx5p33_ASAP7_75t_R g6113 ( 
.A(n_5446),
.Y(n_6113)
);

NOR2x1_ASAP7_75t_SL g6114 ( 
.A(n_5279),
.B(n_5305),
.Y(n_6114)
);

AO31x2_ASAP7_75t_L g6115 ( 
.A1(n_5540),
.A2(n_5069),
.A3(n_5066),
.B(n_4757),
.Y(n_6115)
);

NAND3xp33_ASAP7_75t_SL g6116 ( 
.A(n_5345),
.B(n_4974),
.C(n_4993),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5493),
.Y(n_6117)
);

INVx1_ASAP7_75t_L g6118 ( 
.A(n_5676),
.Y(n_6118)
);

AND2x4_ASAP7_75t_L g6119 ( 
.A(n_5953),
.B(n_5416),
.Y(n_6119)
);

OA21x2_ASAP7_75t_L g6120 ( 
.A1(n_5904),
.A2(n_5971),
.B(n_5955),
.Y(n_6120)
);

AND2x2_ASAP7_75t_L g6121 ( 
.A(n_5727),
.B(n_5185),
.Y(n_6121)
);

NAND2xp5_ASAP7_75t_L g6122 ( 
.A(n_5697),
.B(n_5471),
.Y(n_6122)
);

OR2x2_ASAP7_75t_L g6123 ( 
.A(n_5856),
.B(n_6103),
.Y(n_6123)
);

OR2x6_ASAP7_75t_L g6124 ( 
.A(n_5671),
.B(n_5573),
.Y(n_6124)
);

AND2x2_ASAP7_75t_L g6125 ( 
.A(n_5727),
.B(n_5185),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5676),
.Y(n_6126)
);

BUFx3_ASAP7_75t_L g6127 ( 
.A(n_5703),
.Y(n_6127)
);

AO21x2_ASAP7_75t_L g6128 ( 
.A1(n_5864),
.A2(n_5592),
.B(n_5501),
.Y(n_6128)
);

AND2x4_ASAP7_75t_L g6129 ( 
.A(n_5729),
.B(n_5432),
.Y(n_6129)
);

OAI21x1_ASAP7_75t_L g6130 ( 
.A1(n_5816),
.A2(n_5142),
.B(n_5130),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_5682),
.Y(n_6131)
);

AOI21xp5_ASAP7_75t_SL g6132 ( 
.A1(n_5849),
.A2(n_5381),
.B(n_5442),
.Y(n_6132)
);

INVx2_ASAP7_75t_L g6133 ( 
.A(n_6101),
.Y(n_6133)
);

OR2x6_ASAP7_75t_L g6134 ( 
.A(n_5671),
.B(n_5681),
.Y(n_6134)
);

AO21x2_ASAP7_75t_L g6135 ( 
.A1(n_5746),
.A2(n_5490),
.B(n_5585),
.Y(n_6135)
);

INVx2_ASAP7_75t_L g6136 ( 
.A(n_6101),
.Y(n_6136)
);

AO21x2_ASAP7_75t_L g6137 ( 
.A1(n_5655),
.A2(n_5588),
.B(n_5142),
.Y(n_6137)
);

OR2x2_ASAP7_75t_L g6138 ( 
.A(n_5771),
.B(n_5400),
.Y(n_6138)
);

INVx2_ASAP7_75t_L g6139 ( 
.A(n_6101),
.Y(n_6139)
);

OA21x2_ASAP7_75t_L g6140 ( 
.A1(n_5904),
.A2(n_5499),
.B(n_5616),
.Y(n_6140)
);

AO21x2_ASAP7_75t_L g6141 ( 
.A1(n_5747),
.A2(n_5130),
.B(n_5095),
.Y(n_6141)
);

INVx1_ASAP7_75t_L g6142 ( 
.A(n_5682),
.Y(n_6142)
);

INVx2_ASAP7_75t_SL g6143 ( 
.A(n_5751),
.Y(n_6143)
);

NOR2xp33_ASAP7_75t_L g6144 ( 
.A(n_5652),
.B(n_5312),
.Y(n_6144)
);

AOI22xp33_ASAP7_75t_L g6145 ( 
.A1(n_6083),
.A2(n_5614),
.B1(n_5174),
.B2(n_5498),
.Y(n_6145)
);

AOI22xp33_ASAP7_75t_L g6146 ( 
.A1(n_5674),
.A2(n_5498),
.B1(n_4991),
.B2(n_5140),
.Y(n_6146)
);

AND2x2_ASAP7_75t_L g6147 ( 
.A(n_5729),
.B(n_5338),
.Y(n_6147)
);

AND2x2_ASAP7_75t_L g6148 ( 
.A(n_5757),
.B(n_5338),
.Y(n_6148)
);

NAND2xp5_ASAP7_75t_L g6149 ( 
.A(n_5645),
.B(n_5204),
.Y(n_6149)
);

AO21x2_ASAP7_75t_L g6150 ( 
.A1(n_5747),
.A2(n_5095),
.B(n_5084),
.Y(n_6150)
);

INVx2_ASAP7_75t_L g6151 ( 
.A(n_6101),
.Y(n_6151)
);

AND2x2_ASAP7_75t_L g6152 ( 
.A(n_5757),
.B(n_5544),
.Y(n_6152)
);

INVx1_ASAP7_75t_L g6153 ( 
.A(n_5700),
.Y(n_6153)
);

AND2x2_ASAP7_75t_L g6154 ( 
.A(n_5765),
.B(n_5793),
.Y(n_6154)
);

AND2x2_ASAP7_75t_L g6155 ( 
.A(n_5765),
.B(n_5546),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_5700),
.Y(n_6156)
);

OR2x2_ASAP7_75t_L g6157 ( 
.A(n_5827),
.B(n_5134),
.Y(n_6157)
);

INVx2_ASAP7_75t_L g6158 ( 
.A(n_6115),
.Y(n_6158)
);

HB1xp67_ASAP7_75t_L g6159 ( 
.A(n_5980),
.Y(n_6159)
);

OR2x6_ASAP7_75t_L g6160 ( 
.A(n_5671),
.B(n_5573),
.Y(n_6160)
);

INVx2_ASAP7_75t_L g6161 ( 
.A(n_6115),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_5717),
.Y(n_6162)
);

OAI21xp5_ASAP7_75t_L g6163 ( 
.A1(n_5651),
.A2(n_5381),
.B(n_5376),
.Y(n_6163)
);

INVx1_ASAP7_75t_L g6164 ( 
.A(n_5717),
.Y(n_6164)
);

AND2x2_ASAP7_75t_L g6165 ( 
.A(n_5793),
.B(n_5546),
.Y(n_6165)
);

AND2x2_ASAP7_75t_L g6166 ( 
.A(n_5818),
.B(n_5403),
.Y(n_6166)
);

CKINVDCx5p33_ASAP7_75t_R g6167 ( 
.A(n_5715),
.Y(n_6167)
);

INVx2_ASAP7_75t_L g6168 ( 
.A(n_6115),
.Y(n_6168)
);

AND2x2_ASAP7_75t_L g6169 ( 
.A(n_5818),
.B(n_5097),
.Y(n_6169)
);

OA21x2_ASAP7_75t_L g6170 ( 
.A1(n_5955),
.A2(n_5529),
.B(n_5502),
.Y(n_6170)
);

INVx2_ASAP7_75t_L g6171 ( 
.A(n_6115),
.Y(n_6171)
);

AND2x4_ASAP7_75t_L g6172 ( 
.A(n_5839),
.B(n_5432),
.Y(n_6172)
);

AOI21xp5_ASAP7_75t_SL g6173 ( 
.A1(n_5667),
.A2(n_5442),
.B(n_5384),
.Y(n_6173)
);

INVx4_ASAP7_75t_L g6174 ( 
.A(n_5643),
.Y(n_6174)
);

INVx2_ASAP7_75t_L g6175 ( 
.A(n_5647),
.Y(n_6175)
);

INVxp67_ASAP7_75t_L g6176 ( 
.A(n_5667),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_5776),
.Y(n_6177)
);

AOI22xp33_ASAP7_75t_L g6178 ( 
.A1(n_5674),
.A2(n_5498),
.B1(n_4991),
.B2(n_5140),
.Y(n_6178)
);

INVx2_ASAP7_75t_L g6179 ( 
.A(n_5647),
.Y(n_6179)
);

OR2x2_ASAP7_75t_L g6180 ( 
.A(n_5877),
.B(n_5134),
.Y(n_6180)
);

OR2x6_ASAP7_75t_L g6181 ( 
.A(n_5681),
.B(n_5573),
.Y(n_6181)
);

INVx2_ASAP7_75t_L g6182 ( 
.A(n_5648),
.Y(n_6182)
);

OR2x2_ASAP7_75t_L g6183 ( 
.A(n_5659),
.B(n_5160),
.Y(n_6183)
);

AOI22xp33_ASAP7_75t_L g6184 ( 
.A1(n_5956),
.A2(n_5140),
.B1(n_5118),
.B2(n_5601),
.Y(n_6184)
);

OA21x2_ASAP7_75t_L g6185 ( 
.A1(n_5971),
.A2(n_5340),
.B(n_5112),
.Y(n_6185)
);

INVx3_ASAP7_75t_L g6186 ( 
.A(n_5787),
.Y(n_6186)
);

INVx1_ASAP7_75t_L g6187 ( 
.A(n_5776),
.Y(n_6187)
);

OR2x2_ASAP7_75t_L g6188 ( 
.A(n_5690),
.B(n_5160),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_5815),
.Y(n_6189)
);

INVxp33_ASAP7_75t_L g6190 ( 
.A(n_5715),
.Y(n_6190)
);

INVxp67_ASAP7_75t_SL g6191 ( 
.A(n_5735),
.Y(n_6191)
);

AND2x2_ASAP7_75t_L g6192 ( 
.A(n_5839),
.B(n_5193),
.Y(n_6192)
);

AO21x2_ASAP7_75t_L g6193 ( 
.A1(n_5843),
.A2(n_5095),
.B(n_5084),
.Y(n_6193)
);

AND2x4_ASAP7_75t_L g6194 ( 
.A(n_5896),
.B(n_5432),
.Y(n_6194)
);

INVx1_ASAP7_75t_L g6195 ( 
.A(n_5815),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_5832),
.Y(n_6196)
);

INVx1_ASAP7_75t_L g6197 ( 
.A(n_5832),
.Y(n_6197)
);

AND2x2_ASAP7_75t_L g6198 ( 
.A(n_5896),
.B(n_5193),
.Y(n_6198)
);

BUFx2_ASAP7_75t_L g6199 ( 
.A(n_5683),
.Y(n_6199)
);

OAI33xp33_ASAP7_75t_L g6200 ( 
.A1(n_6076),
.A2(n_5435),
.A3(n_5418),
.B1(n_5423),
.B2(n_5427),
.B3(n_5438),
.Y(n_6200)
);

BUFx2_ASAP7_75t_L g6201 ( 
.A(n_5683),
.Y(n_6201)
);

AND2x2_ASAP7_75t_L g6202 ( 
.A(n_6093),
.B(n_5277),
.Y(n_6202)
);

OA21x2_ASAP7_75t_L g6203 ( 
.A1(n_6032),
.A2(n_5340),
.B(n_5112),
.Y(n_6203)
);

INVx2_ASAP7_75t_L g6204 ( 
.A(n_5648),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_5835),
.Y(n_6205)
);

OAI221xp5_ASAP7_75t_L g6206 ( 
.A1(n_6038),
.A2(n_5322),
.B1(n_5476),
.B2(n_5352),
.C(n_5394),
.Y(n_6206)
);

OR2x6_ASAP7_75t_L g6207 ( 
.A(n_5681),
.B(n_5137),
.Y(n_6207)
);

INVx2_ASAP7_75t_L g6208 ( 
.A(n_5666),
.Y(n_6208)
);

OAI22xp5_ASAP7_75t_L g6209 ( 
.A1(n_5744),
.A2(n_5128),
.B1(n_5304),
.B2(n_5300),
.Y(n_6209)
);

INVx1_ASAP7_75t_SL g6210 ( 
.A(n_5737),
.Y(n_6210)
);

INVx2_ASAP7_75t_L g6211 ( 
.A(n_5666),
.Y(n_6211)
);

INVx2_ASAP7_75t_L g6212 ( 
.A(n_5731),
.Y(n_6212)
);

AND2x2_ASAP7_75t_L g6213 ( 
.A(n_6093),
.B(n_5277),
.Y(n_6213)
);

INVx2_ASAP7_75t_L g6214 ( 
.A(n_5731),
.Y(n_6214)
);

AOI221xp5_ASAP7_75t_L g6215 ( 
.A1(n_6076),
.A2(n_5714),
.B1(n_5730),
.B2(n_5988),
.C(n_5852),
.Y(n_6215)
);

INVx1_ASAP7_75t_L g6216 ( 
.A(n_5835),
.Y(n_6216)
);

NOR2xp33_ASAP7_75t_L g6217 ( 
.A(n_5657),
.B(n_5665),
.Y(n_6217)
);

INVx3_ASAP7_75t_L g6218 ( 
.A(n_5787),
.Y(n_6218)
);

BUFx3_ASAP7_75t_L g6219 ( 
.A(n_5703),
.Y(n_6219)
);

AND2x4_ASAP7_75t_L g6220 ( 
.A(n_5977),
.B(n_5432),
.Y(n_6220)
);

INVx5_ASAP7_75t_L g6221 ( 
.A(n_5686),
.Y(n_6221)
);

INVx2_ASAP7_75t_L g6222 ( 
.A(n_5732),
.Y(n_6222)
);

BUFx6f_ASAP7_75t_L g6223 ( 
.A(n_5643),
.Y(n_6223)
);

AND2x2_ASAP7_75t_L g6224 ( 
.A(n_5844),
.B(n_5315),
.Y(n_6224)
);

AND2x2_ASAP7_75t_L g6225 ( 
.A(n_5844),
.B(n_5315),
.Y(n_6225)
);

INVx2_ASAP7_75t_L g6226 ( 
.A(n_5732),
.Y(n_6226)
);

OAI221xp5_ASAP7_75t_L g6227 ( 
.A1(n_5749),
.A2(n_5203),
.B1(n_5451),
.B2(n_5420),
.C(n_5545),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_L g6228 ( 
.A(n_5784),
.B(n_5361),
.Y(n_6228)
);

BUFx2_ASAP7_75t_L g6229 ( 
.A(n_5673),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_5841),
.Y(n_6230)
);

INVx1_ASAP7_75t_L g6231 ( 
.A(n_5841),
.Y(n_6231)
);

OAI21xp5_ASAP7_75t_L g6232 ( 
.A1(n_5755),
.A2(n_5524),
.B(n_5523),
.Y(n_6232)
);

BUFx3_ASAP7_75t_L g6233 ( 
.A(n_5642),
.Y(n_6233)
);

AND2x2_ASAP7_75t_L g6234 ( 
.A(n_5912),
.B(n_5334),
.Y(n_6234)
);

OR2x6_ASAP7_75t_L g6235 ( 
.A(n_5705),
.B(n_5137),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_5854),
.Y(n_6236)
);

HB1xp67_ASAP7_75t_L g6237 ( 
.A(n_6008),
.Y(n_6237)
);

AND2x2_ASAP7_75t_L g6238 ( 
.A(n_6054),
.B(n_5334),
.Y(n_6238)
);

OR2x2_ASAP7_75t_L g6239 ( 
.A(n_5936),
.B(n_5173),
.Y(n_6239)
);

INVxp67_ASAP7_75t_SL g6240 ( 
.A(n_5792),
.Y(n_6240)
);

INVx2_ASAP7_75t_L g6241 ( 
.A(n_5733),
.Y(n_6241)
);

INVx2_ASAP7_75t_L g6242 ( 
.A(n_5733),
.Y(n_6242)
);

AO21x2_ASAP7_75t_L g6243 ( 
.A1(n_6046),
.A2(n_5123),
.B(n_5084),
.Y(n_6243)
);

INVx3_ASAP7_75t_L g6244 ( 
.A(n_5787),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_5854),
.Y(n_6245)
);

OAI321xp33_ASAP7_75t_L g6246 ( 
.A1(n_5714),
.A2(n_5527),
.A3(n_5562),
.B1(n_5553),
.B2(n_5563),
.C(n_5554),
.Y(n_6246)
);

HB1xp67_ASAP7_75t_L g6247 ( 
.A(n_6029),
.Y(n_6247)
);

BUFx2_ASAP7_75t_SL g6248 ( 
.A(n_5770),
.Y(n_6248)
);

HB1xp67_ASAP7_75t_L g6249 ( 
.A(n_6072),
.Y(n_6249)
);

HB1xp67_ASAP7_75t_L g6250 ( 
.A(n_5767),
.Y(n_6250)
);

INVx2_ASAP7_75t_L g6251 ( 
.A(n_5742),
.Y(n_6251)
);

OR2x2_ASAP7_75t_L g6252 ( 
.A(n_5937),
.B(n_5173),
.Y(n_6252)
);

OA21x2_ASAP7_75t_L g6253 ( 
.A1(n_6032),
.A2(n_5852),
.B(n_5845),
.Y(n_6253)
);

HB1xp67_ASAP7_75t_L g6254 ( 
.A(n_6020),
.Y(n_6254)
);

INVx3_ASAP7_75t_L g6255 ( 
.A(n_6037),
.Y(n_6255)
);

AO21x2_ASAP7_75t_L g6256 ( 
.A1(n_6102),
.A2(n_5123),
.B(n_5116),
.Y(n_6256)
);

BUFx6f_ASAP7_75t_L g6257 ( 
.A(n_5863),
.Y(n_6257)
);

AO21x2_ASAP7_75t_L g6258 ( 
.A1(n_5728),
.A2(n_5123),
.B(n_5116),
.Y(n_6258)
);

AO21x2_ASAP7_75t_L g6259 ( 
.A1(n_5728),
.A2(n_5120),
.B(n_5088),
.Y(n_6259)
);

HB1xp67_ASAP7_75t_L g6260 ( 
.A(n_6020),
.Y(n_6260)
);

NAND2xp5_ASAP7_75t_L g6261 ( 
.A(n_5646),
.B(n_5650),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_5899),
.Y(n_6262)
);

OAI21xp5_ASAP7_75t_L g6263 ( 
.A1(n_5755),
.A2(n_5744),
.B(n_5763),
.Y(n_6263)
);

INVx1_ASAP7_75t_L g6264 ( 
.A(n_5899),
.Y(n_6264)
);

HB1xp67_ASAP7_75t_L g6265 ( 
.A(n_6099),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_5933),
.Y(n_6266)
);

HB1xp67_ASAP7_75t_L g6267 ( 
.A(n_6099),
.Y(n_6267)
);

NAND4xp25_ASAP7_75t_L g6268 ( 
.A(n_5884),
.B(n_5857),
.C(n_5785),
.D(n_5679),
.Y(n_6268)
);

HB1xp67_ASAP7_75t_L g6269 ( 
.A(n_5804),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_5933),
.Y(n_6270)
);

INVx2_ASAP7_75t_L g6271 ( 
.A(n_5742),
.Y(n_6271)
);

INVx2_ASAP7_75t_L g6272 ( 
.A(n_5754),
.Y(n_6272)
);

AND2x2_ASAP7_75t_L g6273 ( 
.A(n_6054),
.B(n_5337),
.Y(n_6273)
);

INVx2_ASAP7_75t_SL g6274 ( 
.A(n_5704),
.Y(n_6274)
);

AND2x2_ASAP7_75t_L g6275 ( 
.A(n_5654),
.B(n_5337),
.Y(n_6275)
);

INVx2_ASAP7_75t_SL g6276 ( 
.A(n_5658),
.Y(n_6276)
);

INVx2_ASAP7_75t_L g6277 ( 
.A(n_5754),
.Y(n_6277)
);

OA21x2_ASAP7_75t_L g6278 ( 
.A1(n_5821),
.A2(n_5120),
.B(n_5088),
.Y(n_6278)
);

AO21x2_ASAP7_75t_L g6279 ( 
.A1(n_5701),
.A2(n_5155),
.B(n_5141),
.Y(n_6279)
);

OR2x2_ASAP7_75t_L g6280 ( 
.A(n_5996),
.B(n_5230),
.Y(n_6280)
);

INVx2_ASAP7_75t_L g6281 ( 
.A(n_5764),
.Y(n_6281)
);

INVx1_ASAP7_75t_L g6282 ( 
.A(n_5974),
.Y(n_6282)
);

OR2x2_ASAP7_75t_L g6283 ( 
.A(n_6004),
.B(n_5230),
.Y(n_6283)
);

AND2x2_ASAP7_75t_L g6284 ( 
.A(n_5654),
.B(n_5532),
.Y(n_6284)
);

OA21x2_ASAP7_75t_L g6285 ( 
.A1(n_5821),
.A2(n_5155),
.B(n_5141),
.Y(n_6285)
);

OR2x2_ASAP7_75t_L g6286 ( 
.A(n_5957),
.B(n_5361),
.Y(n_6286)
);

OAI21xp5_ASAP7_75t_L g6287 ( 
.A1(n_5763),
.A2(n_5253),
.B(n_5601),
.Y(n_6287)
);

AO21x2_ASAP7_75t_L g6288 ( 
.A1(n_5764),
.A2(n_5769),
.B(n_5822),
.Y(n_6288)
);

INVx2_ASAP7_75t_L g6289 ( 
.A(n_5769),
.Y(n_6289)
);

AND2x2_ASAP7_75t_L g6290 ( 
.A(n_5654),
.B(n_5670),
.Y(n_6290)
);

INVx2_ASAP7_75t_L g6291 ( 
.A(n_6048),
.Y(n_6291)
);

NOR2xp33_ASAP7_75t_L g6292 ( 
.A(n_5688),
.B(n_5251),
.Y(n_6292)
);

AND2x2_ASAP7_75t_L g6293 ( 
.A(n_5670),
.B(n_5532),
.Y(n_6293)
);

INVx3_ASAP7_75t_L g6294 ( 
.A(n_6037),
.Y(n_6294)
);

AND2x2_ASAP7_75t_L g6295 ( 
.A(n_5670),
.B(n_5532),
.Y(n_6295)
);

HB1xp67_ASAP7_75t_L g6296 ( 
.A(n_6100),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_5974),
.Y(n_6297)
);

OR2x2_ASAP7_75t_L g6298 ( 
.A(n_5986),
.B(n_5361),
.Y(n_6298)
);

AO21x1_ASAP7_75t_SL g6299 ( 
.A1(n_5672),
.A2(n_5363),
.B(n_4973),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_6105),
.Y(n_6300)
);

INVx2_ASAP7_75t_L g6301 ( 
.A(n_6048),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_6105),
.Y(n_6302)
);

INVx2_ASAP7_75t_L g6303 ( 
.A(n_6064),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_5684),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_5707),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_5725),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_5726),
.Y(n_6307)
);

NOR2xp33_ASAP7_75t_L g6308 ( 
.A(n_5713),
.B(n_5176),
.Y(n_6308)
);

AND2x4_ASAP7_75t_L g6309 ( 
.A(n_5977),
.B(n_5432),
.Y(n_6309)
);

AND2x2_ASAP7_75t_L g6310 ( 
.A(n_5781),
.B(n_5532),
.Y(n_6310)
);

BUFx6f_ASAP7_75t_L g6311 ( 
.A(n_5686),
.Y(n_6311)
);

OA21x2_ASAP7_75t_L g6312 ( 
.A1(n_5845),
.A2(n_5282),
.B(n_5169),
.Y(n_6312)
);

NAND3xp33_ASAP7_75t_L g6313 ( 
.A(n_5947),
.B(n_5344),
.C(n_5458),
.Y(n_6313)
);

OAI21xp5_ASAP7_75t_L g6314 ( 
.A1(n_5947),
.A2(n_5618),
.B(n_5549),
.Y(n_6314)
);

AND2x2_ASAP7_75t_L g6315 ( 
.A(n_5781),
.B(n_5355),
.Y(n_6315)
);

INVx2_ASAP7_75t_L g6316 ( 
.A(n_6064),
.Y(n_6316)
);

AO21x2_ASAP7_75t_L g6317 ( 
.A1(n_5822),
.A2(n_5618),
.B(n_5452),
.Y(n_6317)
);

INVx3_ASAP7_75t_L g6318 ( 
.A(n_6026),
.Y(n_6318)
);

INVx1_ASAP7_75t_L g6319 ( 
.A(n_5759),
.Y(n_6319)
);

AND2x2_ASAP7_75t_L g6320 ( 
.A(n_5893),
.B(n_5216),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_5766),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_5786),
.Y(n_6322)
);

OAI21x1_ASAP7_75t_L g6323 ( 
.A1(n_5641),
.A2(n_5187),
.B(n_5154),
.Y(n_6323)
);

INVx2_ASAP7_75t_L g6324 ( 
.A(n_6070),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_5796),
.Y(n_6325)
);

INVx1_ASAP7_75t_L g6326 ( 
.A(n_5807),
.Y(n_6326)
);

OA21x2_ASAP7_75t_L g6327 ( 
.A1(n_6034),
.A2(n_5898),
.B(n_5641),
.Y(n_6327)
);

OAI21x1_ASAP7_75t_L g6328 ( 
.A1(n_5898),
.A2(n_6034),
.B(n_5789),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_5828),
.Y(n_6329)
);

AOI22xp5_ASAP7_75t_L g6330 ( 
.A1(n_6031),
.A2(n_5194),
.B1(n_5161),
.B2(n_5618),
.Y(n_6330)
);

BUFx2_ASAP7_75t_L g6331 ( 
.A(n_5673),
.Y(n_6331)
);

NAND2xp5_ASAP7_75t_L g6332 ( 
.A(n_5806),
.B(n_5361),
.Y(n_6332)
);

BUFx6f_ASAP7_75t_SL g6333 ( 
.A(n_5687),
.Y(n_6333)
);

OR2x2_ASAP7_75t_L g6334 ( 
.A(n_6005),
.B(n_5361),
.Y(n_6334)
);

OA21x2_ASAP7_75t_L g6335 ( 
.A1(n_5789),
.A2(n_5695),
.B(n_6070),
.Y(n_6335)
);

OAI21xp5_ASAP7_75t_L g6336 ( 
.A1(n_5820),
.A2(n_5541),
.B(n_5241),
.Y(n_6336)
);

OA21x2_ASAP7_75t_L g6337 ( 
.A1(n_5695),
.A2(n_5282),
.B(n_5169),
.Y(n_6337)
);

BUFx2_ASAP7_75t_L g6338 ( 
.A(n_5644),
.Y(n_6338)
);

INVx1_ASAP7_75t_L g6339 ( 
.A(n_5846),
.Y(n_6339)
);

NAND3xp33_ASAP7_75t_L g6340 ( 
.A(n_5749),
.B(n_5344),
.C(n_5485),
.Y(n_6340)
);

OA21x2_ASAP7_75t_L g6341 ( 
.A1(n_6074),
.A2(n_5730),
.B(n_5722),
.Y(n_6341)
);

BUFx3_ASAP7_75t_L g6342 ( 
.A(n_5713),
.Y(n_6342)
);

NAND2xp33_ASAP7_75t_R g6343 ( 
.A(n_5644),
.B(n_5164),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_5848),
.Y(n_6344)
);

INVx2_ASAP7_75t_SL g6345 ( 
.A(n_6050),
.Y(n_6345)
);

AO21x2_ASAP7_75t_L g6346 ( 
.A1(n_5830),
.A2(n_5441),
.B(n_5639),
.Y(n_6346)
);

INVx2_ASAP7_75t_L g6347 ( 
.A(n_6074),
.Y(n_6347)
);

INVx2_ASAP7_75t_L g6348 ( 
.A(n_6063),
.Y(n_6348)
);

AND2x2_ASAP7_75t_L g6349 ( 
.A(n_5901),
.B(n_5216),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_5860),
.Y(n_6350)
);

OAI221xp5_ASAP7_75t_L g6351 ( 
.A1(n_5722),
.A2(n_5276),
.B1(n_5640),
.B2(n_5635),
.C(n_5631),
.Y(n_6351)
);

INVx2_ASAP7_75t_SL g6352 ( 
.A(n_6050),
.Y(n_6352)
);

INVx2_ASAP7_75t_L g6353 ( 
.A(n_6063),
.Y(n_6353)
);

OA21x2_ASAP7_75t_L g6354 ( 
.A1(n_5830),
.A2(n_5144),
.B(n_5117),
.Y(n_6354)
);

INVx2_ASAP7_75t_L g6355 ( 
.A(n_6063),
.Y(n_6355)
);

AND2x2_ASAP7_75t_L g6356 ( 
.A(n_5910),
.B(n_5241),
.Y(n_6356)
);

INVx2_ASAP7_75t_L g6357 ( 
.A(n_6063),
.Y(n_6357)
);

NAND2xp5_ASAP7_75t_L g6358 ( 
.A(n_5978),
.B(n_5362),
.Y(n_6358)
);

OR2x6_ASAP7_75t_L g6359 ( 
.A(n_5705),
.B(n_5706),
.Y(n_6359)
);

AND2x2_ASAP7_75t_L g6360 ( 
.A(n_5739),
.B(n_5570),
.Y(n_6360)
);

INVx1_ASAP7_75t_L g6361 ( 
.A(n_5866),
.Y(n_6361)
);

INVx1_ASAP7_75t_L g6362 ( 
.A(n_5873),
.Y(n_6362)
);

HB1xp67_ASAP7_75t_L g6363 ( 
.A(n_6082),
.Y(n_6363)
);

INVx1_ASAP7_75t_L g6364 ( 
.A(n_5876),
.Y(n_6364)
);

AO21x2_ASAP7_75t_L g6365 ( 
.A1(n_5838),
.A2(n_5639),
.B(n_5577),
.Y(n_6365)
);

AND2x2_ASAP7_75t_L g6366 ( 
.A(n_5739),
.B(n_5570),
.Y(n_6366)
);

AO21x2_ASAP7_75t_L g6367 ( 
.A1(n_5838),
.A2(n_5639),
.B(n_5576),
.Y(n_6367)
);

INVx2_ASAP7_75t_L g6368 ( 
.A(n_6003),
.Y(n_6368)
);

OA21x2_ASAP7_75t_L g6369 ( 
.A1(n_5976),
.A2(n_5144),
.B(n_5117),
.Y(n_6369)
);

NAND2xp5_ASAP7_75t_SL g6370 ( 
.A(n_5984),
.B(n_5410),
.Y(n_6370)
);

INVx1_ASAP7_75t_L g6371 ( 
.A(n_5886),
.Y(n_6371)
);

BUFx2_ASAP7_75t_L g6372 ( 
.A(n_5692),
.Y(n_6372)
);

AND2x2_ASAP7_75t_L g6373 ( 
.A(n_5739),
.B(n_4603),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_5913),
.Y(n_6374)
);

INVxp67_ASAP7_75t_L g6375 ( 
.A(n_5792),
.Y(n_6375)
);

INVx4_ASAP7_75t_L g6376 ( 
.A(n_5687),
.Y(n_6376)
);

INVxp67_ASAP7_75t_L g6377 ( 
.A(n_5857),
.Y(n_6377)
);

NAND2x1_ASAP7_75t_L g6378 ( 
.A(n_5820),
.B(n_5557),
.Y(n_6378)
);

INVx1_ASAP7_75t_L g6379 ( 
.A(n_5920),
.Y(n_6379)
);

NAND3xp33_ASAP7_75t_L g6380 ( 
.A(n_5851),
.B(n_5668),
.C(n_5888),
.Y(n_6380)
);

INVx3_ASAP7_75t_L g6381 ( 
.A(n_5989),
.Y(n_6381)
);

AND2x2_ASAP7_75t_L g6382 ( 
.A(n_5756),
.B(n_4603),
.Y(n_6382)
);

OR2x2_ASAP7_75t_L g6383 ( 
.A(n_6006),
.B(n_5362),
.Y(n_6383)
);

BUFx3_ASAP7_75t_L g6384 ( 
.A(n_5709),
.Y(n_6384)
);

INVx4_ASAP7_75t_L g6385 ( 
.A(n_5687),
.Y(n_6385)
);

OR2x6_ASAP7_75t_L g6386 ( 
.A(n_5705),
.B(n_5137),
.Y(n_6386)
);

AND2x4_ASAP7_75t_L g6387 ( 
.A(n_5983),
.B(n_5279),
.Y(n_6387)
);

HB1xp67_ASAP7_75t_L g6388 ( 
.A(n_5677),
.Y(n_6388)
);

AND2x2_ASAP7_75t_L g6389 ( 
.A(n_5756),
.B(n_4603),
.Y(n_6389)
);

AOI222xp33_ASAP7_75t_L g6390 ( 
.A1(n_5878),
.A2(n_5406),
.B1(n_5392),
.B2(n_5556),
.C1(n_5539),
.C2(n_5533),
.Y(n_6390)
);

INVx1_ASAP7_75t_L g6391 ( 
.A(n_5943),
.Y(n_6391)
);

AND2x4_ASAP7_75t_L g6392 ( 
.A(n_5983),
.B(n_5305),
.Y(n_6392)
);

BUFx2_ASAP7_75t_L g6393 ( 
.A(n_5692),
.Y(n_6393)
);

INVx2_ASAP7_75t_SL g6394 ( 
.A(n_5805),
.Y(n_6394)
);

INVx2_ASAP7_75t_L g6395 ( 
.A(n_6003),
.Y(n_6395)
);

AO21x2_ASAP7_75t_L g6396 ( 
.A1(n_5870),
.A2(n_5166),
.B(n_5165),
.Y(n_6396)
);

AOI22xp33_ASAP7_75t_L g6397 ( 
.A1(n_6053),
.A2(n_5118),
.B1(n_5248),
.B2(n_5044),
.Y(n_6397)
);

OA21x2_ASAP7_75t_L g6398 ( 
.A1(n_6062),
.A2(n_4740),
.B(n_4733),
.Y(n_6398)
);

BUFx2_ASAP7_75t_L g6399 ( 
.A(n_5711),
.Y(n_6399)
);

AOI21xp33_ASAP7_75t_L g6400 ( 
.A1(n_5668),
.A2(n_4626),
.B(n_5344),
.Y(n_6400)
);

INVx1_ASAP7_75t_L g6401 ( 
.A(n_5944),
.Y(n_6401)
);

AO21x2_ASAP7_75t_L g6402 ( 
.A1(n_5991),
.A2(n_5166),
.B(n_5165),
.Y(n_6402)
);

HB1xp67_ASAP7_75t_L g6403 ( 
.A(n_5680),
.Y(n_6403)
);

AOI22xp33_ASAP7_75t_L g6404 ( 
.A1(n_5859),
.A2(n_5118),
.B1(n_5248),
.B2(n_5044),
.Y(n_6404)
);

AND2x2_ASAP7_75t_L g6405 ( 
.A(n_5756),
.B(n_4603),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_5961),
.Y(n_6406)
);

OAI21xp5_ASAP7_75t_L g6407 ( 
.A1(n_5851),
.A2(n_5542),
.B(n_5399),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_5962),
.Y(n_6408)
);

AND2x2_ASAP7_75t_L g6409 ( 
.A(n_5833),
.B(n_4603),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_5966),
.Y(n_6410)
);

AOI21xp5_ASAP7_75t_SL g6411 ( 
.A1(n_5750),
.A2(n_5231),
.B(n_5305),
.Y(n_6411)
);

INVx1_ASAP7_75t_L g6412 ( 
.A(n_5969),
.Y(n_6412)
);

OA21x2_ASAP7_75t_L g6413 ( 
.A1(n_6062),
.A2(n_4740),
.B(n_4733),
.Y(n_6413)
);

OAI21x1_ASAP7_75t_L g6414 ( 
.A1(n_5753),
.A2(n_5775),
.B(n_5649),
.Y(n_6414)
);

INVxp67_ASAP7_75t_L g6415 ( 
.A(n_5687),
.Y(n_6415)
);

AOI22xp33_ASAP7_75t_L g6416 ( 
.A1(n_6080),
.A2(n_5248),
.B1(n_5044),
.B2(n_4934),
.Y(n_6416)
);

INVx2_ASAP7_75t_L g6417 ( 
.A(n_6003),
.Y(n_6417)
);

INVx2_ASAP7_75t_L g6418 ( 
.A(n_6003),
.Y(n_6418)
);

OA21x2_ASAP7_75t_L g6419 ( 
.A1(n_6012),
.A2(n_4740),
.B(n_4733),
.Y(n_6419)
);

HB1xp67_ASAP7_75t_L g6420 ( 
.A(n_5808),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_5981),
.Y(n_6421)
);

OR2x2_ASAP7_75t_L g6422 ( 
.A(n_5875),
.B(n_5362),
.Y(n_6422)
);

INVxp33_ASAP7_75t_L g6423 ( 
.A(n_5736),
.Y(n_6423)
);

AND2x2_ASAP7_75t_L g6424 ( 
.A(n_5833),
.B(n_5154),
.Y(n_6424)
);

INVx1_ASAP7_75t_L g6425 ( 
.A(n_5987),
.Y(n_6425)
);

AND2x2_ASAP7_75t_L g6426 ( 
.A(n_5833),
.B(n_5154),
.Y(n_6426)
);

AND2x4_ASAP7_75t_L g6427 ( 
.A(n_6092),
.B(n_5305),
.Y(n_6427)
);

OR2x2_ASAP7_75t_L g6428 ( 
.A(n_6024),
.B(n_5362),
.Y(n_6428)
);

BUFx2_ASAP7_75t_L g6429 ( 
.A(n_5711),
.Y(n_6429)
);

AND2x2_ASAP7_75t_L g6430 ( 
.A(n_5850),
.B(n_5798),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_5997),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_6013),
.Y(n_6432)
);

AOI21x1_ASAP7_75t_L g6433 ( 
.A1(n_5780),
.A2(n_4973),
.B(n_4912),
.Y(n_6433)
);

INVx1_ASAP7_75t_L g6434 ( 
.A(n_6021),
.Y(n_6434)
);

AO21x2_ASAP7_75t_L g6435 ( 
.A1(n_5991),
.A2(n_5178),
.B(n_5177),
.Y(n_6435)
);

INVx1_ASAP7_75t_L g6436 ( 
.A(n_6028),
.Y(n_6436)
);

OA21x2_ASAP7_75t_L g6437 ( 
.A1(n_6012),
.A2(n_5109),
.B(n_5177),
.Y(n_6437)
);

INVx3_ASAP7_75t_L g6438 ( 
.A(n_5989),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6035),
.Y(n_6439)
);

OA21x2_ASAP7_75t_L g6440 ( 
.A1(n_6036),
.A2(n_5109),
.B(n_5178),
.Y(n_6440)
);

INVx2_ASAP7_75t_L g6441 ( 
.A(n_6036),
.Y(n_6441)
);

AOI22xp33_ASAP7_75t_L g6442 ( 
.A1(n_6116),
.A2(n_5761),
.B1(n_5738),
.B2(n_5678),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_6039),
.Y(n_6443)
);

INVx1_ASAP7_75t_L g6444 ( 
.A(n_6043),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_6088),
.Y(n_6445)
);

AND2x2_ASAP7_75t_L g6446 ( 
.A(n_5850),
.B(n_5798),
.Y(n_6446)
);

AND2x2_ASAP7_75t_L g6447 ( 
.A(n_5850),
.B(n_5187),
.Y(n_6447)
);

OA21x2_ASAP7_75t_L g6448 ( 
.A1(n_6045),
.A2(n_5916),
.B(n_5914),
.Y(n_6448)
);

BUFx3_ASAP7_75t_L g6449 ( 
.A(n_5719),
.Y(n_6449)
);

HB1xp67_ASAP7_75t_L g6450 ( 
.A(n_5858),
.Y(n_6450)
);

AND2x4_ASAP7_75t_L g6451 ( 
.A(n_6092),
.B(n_5362),
.Y(n_6451)
);

BUFx3_ASAP7_75t_L g6452 ( 
.A(n_5723),
.Y(n_6452)
);

AND2x2_ASAP7_75t_L g6453 ( 
.A(n_5736),
.B(n_5187),
.Y(n_6453)
);

CKINVDCx14_ASAP7_75t_R g6454 ( 
.A(n_5689),
.Y(n_6454)
);

AND2x4_ASAP7_75t_L g6455 ( 
.A(n_6019),
.B(n_5366),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_6091),
.Y(n_6456)
);

AND2x2_ASAP7_75t_L g6457 ( 
.A(n_5934),
.B(n_5919),
.Y(n_6457)
);

AND2x4_ASAP7_75t_L g6458 ( 
.A(n_6019),
.B(n_5366),
.Y(n_6458)
);

AO31x2_ASAP7_75t_L g6459 ( 
.A1(n_5914),
.A2(n_5289),
.A3(n_5317),
.B(n_5260),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_6117),
.Y(n_6460)
);

AOI22xp33_ASAP7_75t_SL g6461 ( 
.A1(n_6040),
.A2(n_5407),
.B1(n_5415),
.B2(n_5231),
.Y(n_6461)
);

INVx1_ASAP7_75t_L g6462 ( 
.A(n_5882),
.Y(n_6462)
);

INVx2_ASAP7_75t_L g6463 ( 
.A(n_6045),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_5882),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_5882),
.Y(n_6465)
);

HB1xp67_ASAP7_75t_L g6466 ( 
.A(n_5982),
.Y(n_6466)
);

BUFx3_ASAP7_75t_L g6467 ( 
.A(n_5721),
.Y(n_6467)
);

AND2x2_ASAP7_75t_L g6468 ( 
.A(n_5941),
.B(n_5693),
.Y(n_6468)
);

INVx2_ASAP7_75t_L g6469 ( 
.A(n_5696),
.Y(n_6469)
);

INVx1_ASAP7_75t_L g6470 ( 
.A(n_5882),
.Y(n_6470)
);

AND2x2_ASAP7_75t_L g6471 ( 
.A(n_5941),
.B(n_5365),
.Y(n_6471)
);

NOR3xp33_ASAP7_75t_L g6472 ( 
.A(n_5824),
.B(n_5837),
.C(n_5938),
.Y(n_6472)
);

AOI22xp33_ASAP7_75t_L g6473 ( 
.A1(n_5897),
.A2(n_4934),
.B1(n_4896),
.B2(n_4758),
.Y(n_6473)
);

OAI21xp5_ASAP7_75t_L g6474 ( 
.A1(n_5888),
.A2(n_5575),
.B(n_5561),
.Y(n_6474)
);

AND2x4_ASAP7_75t_L g6475 ( 
.A(n_6022),
.B(n_5366),
.Y(n_6475)
);

OAI33xp33_ASAP7_75t_L g6476 ( 
.A1(n_5656),
.A2(n_5427),
.A3(n_5613),
.B1(n_5602),
.B2(n_5582),
.B3(n_5566),
.Y(n_6476)
);

OR2x6_ASAP7_75t_L g6477 ( 
.A(n_5706),
.B(n_5137),
.Y(n_6477)
);

INVx1_ASAP7_75t_L g6478 ( 
.A(n_5810),
.Y(n_6478)
);

AO21x2_ASAP7_75t_L g6479 ( 
.A1(n_5884),
.A2(n_5289),
.B(n_5260),
.Y(n_6479)
);

INVx2_ASAP7_75t_L g6480 ( 
.A(n_5696),
.Y(n_6480)
);

INVx2_ASAP7_75t_L g6481 ( 
.A(n_5696),
.Y(n_6481)
);

BUFx6f_ASAP7_75t_L g6482 ( 
.A(n_5710),
.Y(n_6482)
);

AO21x2_ASAP7_75t_L g6483 ( 
.A1(n_5872),
.A2(n_5894),
.B(n_5889),
.Y(n_6483)
);

NAND2xp5_ASAP7_75t_L g6484 ( 
.A(n_5752),
.B(n_5366),
.Y(n_6484)
);

INVx1_ASAP7_75t_L g6485 ( 
.A(n_5810),
.Y(n_6485)
);

INVx2_ASAP7_75t_L g6486 ( 
.A(n_5696),
.Y(n_6486)
);

AO21x2_ASAP7_75t_L g6487 ( 
.A1(n_5872),
.A2(n_5327),
.B(n_5317),
.Y(n_6487)
);

OA21x2_ASAP7_75t_L g6488 ( 
.A1(n_5916),
.A2(n_5390),
.B(n_5327),
.Y(n_6488)
);

AND2x2_ASAP7_75t_L g6489 ( 
.A(n_5760),
.B(n_5365),
.Y(n_6489)
);

OA21x2_ASAP7_75t_L g6490 ( 
.A1(n_5924),
.A2(n_5939),
.B(n_6111),
.Y(n_6490)
);

AOI21x1_ASAP7_75t_L g6491 ( 
.A1(n_5813),
.A2(n_5029),
.B(n_4912),
.Y(n_6491)
);

OA21x2_ASAP7_75t_L g6492 ( 
.A1(n_5924),
.A2(n_5424),
.B(n_5390),
.Y(n_6492)
);

AND2x2_ASAP7_75t_L g6493 ( 
.A(n_5762),
.B(n_5365),
.Y(n_6493)
);

INVx2_ASAP7_75t_L g6494 ( 
.A(n_5698),
.Y(n_6494)
);

BUFx3_ASAP7_75t_L g6495 ( 
.A(n_5748),
.Y(n_6495)
);

BUFx2_ASAP7_75t_L g6496 ( 
.A(n_5689),
.Y(n_6496)
);

INVx1_ASAP7_75t_L g6497 ( 
.A(n_5810),
.Y(n_6497)
);

INVx2_ASAP7_75t_SL g6498 ( 
.A(n_5718),
.Y(n_6498)
);

OA21x2_ASAP7_75t_L g6499 ( 
.A1(n_5939),
.A2(n_5429),
.B(n_5424),
.Y(n_6499)
);

OAI21xp5_ASAP7_75t_L g6500 ( 
.A1(n_5925),
.A2(n_5412),
.B(n_5468),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_5810),
.Y(n_6501)
);

AND2x2_ASAP7_75t_L g6502 ( 
.A(n_5772),
.B(n_5619),
.Y(n_6502)
);

INVx5_ASAP7_75t_SL g6503 ( 
.A(n_5710),
.Y(n_6503)
);

INVx2_ASAP7_75t_L g6504 ( 
.A(n_5698),
.Y(n_6504)
);

HB1xp67_ASAP7_75t_L g6505 ( 
.A(n_5826),
.Y(n_6505)
);

OR2x6_ASAP7_75t_L g6506 ( 
.A(n_5706),
.B(n_5593),
.Y(n_6506)
);

OAI21xp5_ASAP7_75t_L g6507 ( 
.A1(n_5925),
.A2(n_5262),
.B(n_5520),
.Y(n_6507)
);

INVx2_ASAP7_75t_L g6508 ( 
.A(n_5698),
.Y(n_6508)
);

INVx2_ASAP7_75t_L g6509 ( 
.A(n_5698),
.Y(n_6509)
);

AND2x2_ASAP7_75t_L g6510 ( 
.A(n_5777),
.B(n_5231),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_5902),
.Y(n_6511)
);

BUFx3_ASAP7_75t_L g6512 ( 
.A(n_5768),
.Y(n_6512)
);

INVx2_ASAP7_75t_L g6513 ( 
.A(n_5708),
.Y(n_6513)
);

AND2x4_ASAP7_75t_L g6514 ( 
.A(n_6022),
.B(n_5366),
.Y(n_6514)
);

AO21x2_ASAP7_75t_L g6515 ( 
.A1(n_5889),
.A2(n_5460),
.B(n_5429),
.Y(n_6515)
);

NOR2xp33_ASAP7_75t_L g6516 ( 
.A(n_6257),
.B(n_5758),
.Y(n_6516)
);

AND2x4_ASAP7_75t_L g6517 ( 
.A(n_6143),
.B(n_5829),
.Y(n_6517)
);

INVxp67_ASAP7_75t_SL g6518 ( 
.A(n_6217),
.Y(n_6518)
);

INVx2_ASAP7_75t_L g6519 ( 
.A(n_6150),
.Y(n_6519)
);

INVx1_ASAP7_75t_L g6520 ( 
.A(n_6269),
.Y(n_6520)
);

INVx2_ASAP7_75t_L g6521 ( 
.A(n_6150),
.Y(n_6521)
);

INVx1_ASAP7_75t_L g6522 ( 
.A(n_6250),
.Y(n_6522)
);

INVx1_ASAP7_75t_SL g6523 ( 
.A(n_6248),
.Y(n_6523)
);

INVx1_ASAP7_75t_L g6524 ( 
.A(n_6118),
.Y(n_6524)
);

INVx1_ASAP7_75t_L g6525 ( 
.A(n_6118),
.Y(n_6525)
);

INVx2_ASAP7_75t_L g6526 ( 
.A(n_6150),
.Y(n_6526)
);

INVx3_ASAP7_75t_L g6527 ( 
.A(n_6479),
.Y(n_6527)
);

AND2x4_ASAP7_75t_L g6528 ( 
.A(n_6143),
.B(n_5710),
.Y(n_6528)
);

NAND2xp5_ASAP7_75t_L g6529 ( 
.A(n_6191),
.B(n_5964),
.Y(n_6529)
);

NAND2xp5_ASAP7_75t_L g6530 ( 
.A(n_6261),
.B(n_6104),
.Y(n_6530)
);

AOI221xp5_ASAP7_75t_L g6531 ( 
.A1(n_6215),
.A2(n_5694),
.B1(n_5662),
.B2(n_6104),
.C(n_5685),
.Y(n_6531)
);

OR2x2_ASAP7_75t_L g6532 ( 
.A(n_6123),
.B(n_5773),
.Y(n_6532)
);

INVx2_ASAP7_75t_L g6533 ( 
.A(n_6141),
.Y(n_6533)
);

NOR2xp67_ASAP7_75t_L g6534 ( 
.A(n_6274),
.B(n_5922),
.Y(n_6534)
);

OR2x2_ASAP7_75t_L g6535 ( 
.A(n_6123),
.B(n_5891),
.Y(n_6535)
);

INVx1_ASAP7_75t_L g6536 ( 
.A(n_6126),
.Y(n_6536)
);

BUFx2_ASAP7_75t_L g6537 ( 
.A(n_6199),
.Y(n_6537)
);

AND2x2_ASAP7_75t_L g6538 ( 
.A(n_6121),
.B(n_6125),
.Y(n_6538)
);

INVx2_ASAP7_75t_L g6539 ( 
.A(n_6141),
.Y(n_6539)
);

AOI22xp33_ASAP7_75t_L g6540 ( 
.A1(n_6128),
.A2(n_5894),
.B1(n_5903),
.B2(n_5979),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_6126),
.Y(n_6541)
);

INVx1_ASAP7_75t_L g6542 ( 
.A(n_6142),
.Y(n_6542)
);

AND2x2_ASAP7_75t_L g6543 ( 
.A(n_6121),
.B(n_5868),
.Y(n_6543)
);

INVx2_ASAP7_75t_SL g6544 ( 
.A(n_6274),
.Y(n_6544)
);

AND2x2_ASAP7_75t_L g6545 ( 
.A(n_6125),
.B(n_5819),
.Y(n_6545)
);

BUFx2_ASAP7_75t_L g6546 ( 
.A(n_6199),
.Y(n_6546)
);

AND2x2_ASAP7_75t_L g6547 ( 
.A(n_6468),
.B(n_5819),
.Y(n_6547)
);

INVx2_ASAP7_75t_L g6548 ( 
.A(n_6141),
.Y(n_6548)
);

AND2x2_ASAP7_75t_L g6549 ( 
.A(n_6468),
.B(n_5883),
.Y(n_6549)
);

AND2x2_ASAP7_75t_L g6550 ( 
.A(n_6394),
.B(n_5653),
.Y(n_6550)
);

HB1xp67_ASAP7_75t_L g6551 ( 
.A(n_6186),
.Y(n_6551)
);

INVx4_ASAP7_75t_L g6552 ( 
.A(n_6127),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_6142),
.Y(n_6553)
);

INVx1_ASAP7_75t_L g6554 ( 
.A(n_6177),
.Y(n_6554)
);

INVxp67_ASAP7_75t_SL g6555 ( 
.A(n_6342),
.Y(n_6555)
);

HB1xp67_ASAP7_75t_L g6556 ( 
.A(n_6186),
.Y(n_6556)
);

HB1xp67_ASAP7_75t_L g6557 ( 
.A(n_6186),
.Y(n_6557)
);

NAND2xp5_ASAP7_75t_L g6558 ( 
.A(n_6128),
.B(n_5791),
.Y(n_6558)
);

AND2x2_ASAP7_75t_L g6559 ( 
.A(n_6166),
.B(n_5883),
.Y(n_6559)
);

INVx1_ASAP7_75t_SL g6560 ( 
.A(n_6248),
.Y(n_6560)
);

OR2x2_ASAP7_75t_L g6561 ( 
.A(n_6122),
.B(n_5892),
.Y(n_6561)
);

NAND2xp5_ASAP7_75t_L g6562 ( 
.A(n_6128),
.B(n_5794),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_6177),
.Y(n_6563)
);

AOI22xp33_ASAP7_75t_L g6564 ( 
.A1(n_6315),
.A2(n_6380),
.B1(n_6149),
.B2(n_6135),
.Y(n_6564)
);

HB1xp67_ASAP7_75t_L g6565 ( 
.A(n_6218),
.Y(n_6565)
);

INVx1_ASAP7_75t_L g6566 ( 
.A(n_6187),
.Y(n_6566)
);

INVx1_ASAP7_75t_L g6567 ( 
.A(n_6187),
.Y(n_6567)
);

BUFx6f_ASAP7_75t_L g6568 ( 
.A(n_6127),
.Y(n_6568)
);

BUFx2_ASAP7_75t_L g6569 ( 
.A(n_6201),
.Y(n_6569)
);

NAND2xp5_ASAP7_75t_L g6570 ( 
.A(n_6296),
.B(n_5710),
.Y(n_6570)
);

NAND2xp5_ASAP7_75t_L g6571 ( 
.A(n_6315),
.B(n_5817),
.Y(n_6571)
);

BUFx2_ASAP7_75t_L g6572 ( 
.A(n_6201),
.Y(n_6572)
);

BUFx2_ASAP7_75t_L g6573 ( 
.A(n_6176),
.Y(n_6573)
);

OAI22xp33_ASAP7_75t_L g6574 ( 
.A1(n_6163),
.A2(n_5716),
.B1(n_5803),
.B2(n_5799),
.Y(n_6574)
);

INVx1_ASAP7_75t_L g6575 ( 
.A(n_6189),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_6189),
.Y(n_6576)
);

INVx2_ASAP7_75t_L g6577 ( 
.A(n_6243),
.Y(n_6577)
);

INVx1_ASAP7_75t_L g6578 ( 
.A(n_6195),
.Y(n_6578)
);

OAI221xp5_ASAP7_75t_SL g6579 ( 
.A1(n_6132),
.A2(n_6002),
.B1(n_5918),
.B2(n_6095),
.C(n_6069),
.Y(n_6579)
);

AOI22xp33_ASAP7_75t_L g6580 ( 
.A1(n_6135),
.A2(n_5903),
.B1(n_4626),
.B2(n_5415),
.Y(n_6580)
);

INVx2_ASAP7_75t_L g6581 ( 
.A(n_6243),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_6195),
.Y(n_6582)
);

OR2x2_ASAP7_75t_L g6583 ( 
.A(n_6138),
.B(n_6042),
.Y(n_6583)
);

AND2x2_ASAP7_75t_L g6584 ( 
.A(n_6394),
.B(n_5653),
.Y(n_6584)
);

BUFx6f_ASAP7_75t_L g6585 ( 
.A(n_6219),
.Y(n_6585)
);

INVx1_ASAP7_75t_L g6586 ( 
.A(n_6196),
.Y(n_6586)
);

INVx1_ASAP7_75t_L g6587 ( 
.A(n_6196),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_6197),
.Y(n_6588)
);

AND2x2_ASAP7_75t_L g6589 ( 
.A(n_6345),
.B(n_6352),
.Y(n_6589)
);

AOI22xp33_ASAP7_75t_SL g6590 ( 
.A1(n_6292),
.A2(n_6015),
.B1(n_5800),
.B2(n_6055),
.Y(n_6590)
);

INVx2_ASAP7_75t_L g6591 ( 
.A(n_6243),
.Y(n_6591)
);

AND2x2_ASAP7_75t_SL g6592 ( 
.A(n_6229),
.B(n_6007),
.Y(n_6592)
);

AND2x2_ASAP7_75t_L g6593 ( 
.A(n_6345),
.B(n_5812),
.Y(n_6593)
);

NAND2x1p5_ASAP7_75t_L g6594 ( 
.A(n_6376),
.B(n_5663),
.Y(n_6594)
);

INVx1_ASAP7_75t_L g6595 ( 
.A(n_6197),
.Y(n_6595)
);

AND2x2_ASAP7_75t_L g6596 ( 
.A(n_6352),
.B(n_5814),
.Y(n_6596)
);

NAND2xp5_ASAP7_75t_L g6597 ( 
.A(n_6254),
.B(n_5905),
.Y(n_6597)
);

INVx1_ASAP7_75t_L g6598 ( 
.A(n_6205),
.Y(n_6598)
);

INVx1_ASAP7_75t_L g6599 ( 
.A(n_6205),
.Y(n_6599)
);

BUFx2_ASAP7_75t_L g6600 ( 
.A(n_6229),
.Y(n_6600)
);

NOR2xp33_ASAP7_75t_L g6601 ( 
.A(n_6257),
.B(n_5831),
.Y(n_6601)
);

NAND2xp5_ASAP7_75t_L g6602 ( 
.A(n_6260),
.B(n_5992),
.Y(n_6602)
);

AND2x2_ASAP7_75t_L g6603 ( 
.A(n_6154),
.B(n_5834),
.Y(n_6603)
);

INVx1_ASAP7_75t_L g6604 ( 
.A(n_6216),
.Y(n_6604)
);

INVx2_ASAP7_75t_L g6605 ( 
.A(n_6479),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_6216),
.Y(n_6606)
);

INVx1_ASAP7_75t_L g6607 ( 
.A(n_6230),
.Y(n_6607)
);

INVx2_ASAP7_75t_L g6608 ( 
.A(n_6479),
.Y(n_6608)
);

BUFx2_ASAP7_75t_L g6609 ( 
.A(n_6331),
.Y(n_6609)
);

NAND2xp5_ASAP7_75t_L g6610 ( 
.A(n_6265),
.B(n_5992),
.Y(n_6610)
);

INVxp67_ASAP7_75t_L g6611 ( 
.A(n_6338),
.Y(n_6611)
);

BUFx2_ASAP7_75t_L g6612 ( 
.A(n_6331),
.Y(n_6612)
);

INVx1_ASAP7_75t_L g6613 ( 
.A(n_6230),
.Y(n_6613)
);

OR2x2_ASAP7_75t_L g6614 ( 
.A(n_6138),
.B(n_6052),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_6231),
.Y(n_6615)
);

NOR2xp67_ASAP7_75t_L g6616 ( 
.A(n_6167),
.B(n_5664),
.Y(n_6616)
);

INVx2_ASAP7_75t_L g6617 ( 
.A(n_6193),
.Y(n_6617)
);

OR2x2_ASAP7_75t_L g6618 ( 
.A(n_6420),
.B(n_6450),
.Y(n_6618)
);

BUFx2_ASAP7_75t_L g6619 ( 
.A(n_6338),
.Y(n_6619)
);

HB1xp67_ASAP7_75t_L g6620 ( 
.A(n_6218),
.Y(n_6620)
);

AOI22xp33_ASAP7_75t_L g6621 ( 
.A1(n_6135),
.A2(n_4626),
.B1(n_5415),
.B2(n_5407),
.Y(n_6621)
);

INVx1_ASAP7_75t_L g6622 ( 
.A(n_6231),
.Y(n_6622)
);

AND2x2_ASAP7_75t_L g6623 ( 
.A(n_6166),
.B(n_5842),
.Y(n_6623)
);

INVx2_ASAP7_75t_L g6624 ( 
.A(n_6193),
.Y(n_6624)
);

INVxp67_ASAP7_75t_L g6625 ( 
.A(n_6342),
.Y(n_6625)
);

AND2x2_ASAP7_75t_L g6626 ( 
.A(n_6263),
.B(n_6310),
.Y(n_6626)
);

INVx1_ASAP7_75t_L g6627 ( 
.A(n_6236),
.Y(n_6627)
);

BUFx3_ASAP7_75t_L g6628 ( 
.A(n_6257),
.Y(n_6628)
);

AND2x4_ASAP7_75t_L g6629 ( 
.A(n_6240),
.B(n_6057),
.Y(n_6629)
);

INVx1_ASAP7_75t_L g6630 ( 
.A(n_6236),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_6310),
.B(n_5718),
.Y(n_6631)
);

INVx2_ASAP7_75t_L g6632 ( 
.A(n_6193),
.Y(n_6632)
);

NOR2xp33_ASAP7_75t_L g6633 ( 
.A(n_6257),
.B(n_5740),
.Y(n_6633)
);

NAND2xp5_ASAP7_75t_L g6634 ( 
.A(n_6267),
.B(n_6056),
.Y(n_6634)
);

INVx1_ASAP7_75t_L g6635 ( 
.A(n_6245),
.Y(n_6635)
);

INVx1_ASAP7_75t_L g6636 ( 
.A(n_6245),
.Y(n_6636)
);

AOI22xp33_ASAP7_75t_L g6637 ( 
.A1(n_6327),
.A2(n_4626),
.B1(n_5407),
.B2(n_4610),
.Y(n_6637)
);

NAND2xp5_ASAP7_75t_L g6638 ( 
.A(n_6505),
.B(n_6056),
.Y(n_6638)
);

AND2x4_ASAP7_75t_L g6639 ( 
.A(n_6154),
.B(n_6057),
.Y(n_6639)
);

NAND2xp5_ASAP7_75t_L g6640 ( 
.A(n_6377),
.B(n_6018),
.Y(n_6640)
);

INVx2_ASAP7_75t_L g6641 ( 
.A(n_6469),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_6262),
.Y(n_6642)
);

HB1xp67_ASAP7_75t_L g6643 ( 
.A(n_6218),
.Y(n_6643)
);

INVx2_ASAP7_75t_L g6644 ( 
.A(n_6469),
.Y(n_6644)
);

AND2x2_ASAP7_75t_L g6645 ( 
.A(n_6202),
.B(n_5940),
.Y(n_6645)
);

INVxp67_ASAP7_75t_SL g6646 ( 
.A(n_6257),
.Y(n_6646)
);

OR2x2_ASAP7_75t_L g6647 ( 
.A(n_6466),
.B(n_6094),
.Y(n_6647)
);

AND2x4_ASAP7_75t_L g6648 ( 
.A(n_6376),
.B(n_6065),
.Y(n_6648)
);

NAND2x1p5_ASAP7_75t_L g6649 ( 
.A(n_6376),
.B(n_5663),
.Y(n_6649)
);

AND2x2_ASAP7_75t_L g6650 ( 
.A(n_6202),
.B(n_5940),
.Y(n_6650)
);

INVx2_ASAP7_75t_L g6651 ( 
.A(n_6480),
.Y(n_6651)
);

AND2x2_ASAP7_75t_L g6652 ( 
.A(n_6213),
.B(n_5871),
.Y(n_6652)
);

AND2x2_ASAP7_75t_L g6653 ( 
.A(n_6213),
.B(n_5871),
.Y(n_6653)
);

NAND2xp5_ASAP7_75t_L g6654 ( 
.A(n_6363),
.B(n_5795),
.Y(n_6654)
);

OR2x2_ASAP7_75t_L g6655 ( 
.A(n_6183),
.B(n_5825),
.Y(n_6655)
);

INVx1_ASAP7_75t_L g6656 ( 
.A(n_6262),
.Y(n_6656)
);

INVx1_ASAP7_75t_L g6657 ( 
.A(n_6264),
.Y(n_6657)
);

AND2x2_ASAP7_75t_L g6658 ( 
.A(n_6169),
.B(n_5921),
.Y(n_6658)
);

AOI22xp33_ASAP7_75t_L g6659 ( 
.A1(n_6327),
.A2(n_6404),
.B1(n_6170),
.B2(n_6140),
.Y(n_6659)
);

INVx2_ASAP7_75t_L g6660 ( 
.A(n_6480),
.Y(n_6660)
);

AND2x2_ASAP7_75t_L g6661 ( 
.A(n_6169),
.B(n_5927),
.Y(n_6661)
);

OAI22xp5_ASAP7_75t_L g6662 ( 
.A1(n_6442),
.A2(n_5885),
.B1(n_5699),
.B2(n_5778),
.Y(n_6662)
);

AND2x2_ASAP7_75t_L g6663 ( 
.A(n_6147),
.B(n_5942),
.Y(n_6663)
);

BUFx2_ASAP7_75t_L g6664 ( 
.A(n_6384),
.Y(n_6664)
);

INVx1_ASAP7_75t_L g6665 ( 
.A(n_6264),
.Y(n_6665)
);

OR2x2_ASAP7_75t_L g6666 ( 
.A(n_6183),
.B(n_6001),
.Y(n_6666)
);

INVx2_ASAP7_75t_L g6667 ( 
.A(n_6481),
.Y(n_6667)
);

INVxp67_ASAP7_75t_L g6668 ( 
.A(n_6159),
.Y(n_6668)
);

NOR2xp67_ASAP7_75t_L g6669 ( 
.A(n_6167),
.B(n_5664),
.Y(n_6669)
);

AND2x2_ASAP7_75t_L g6670 ( 
.A(n_6457),
.B(n_5928),
.Y(n_6670)
);

AND2x2_ASAP7_75t_L g6671 ( 
.A(n_6457),
.B(n_5948),
.Y(n_6671)
);

INVx3_ASAP7_75t_L g6672 ( 
.A(n_6259),
.Y(n_6672)
);

AND2x2_ASAP7_75t_L g6673 ( 
.A(n_6496),
.B(n_5865),
.Y(n_6673)
);

INVx2_ASAP7_75t_L g6674 ( 
.A(n_6481),
.Y(n_6674)
);

AOI22xp5_ASAP7_75t_L g6675 ( 
.A1(n_6145),
.A2(n_5862),
.B1(n_5799),
.B2(n_5855),
.Y(n_6675)
);

AND2x2_ASAP7_75t_L g6676 ( 
.A(n_6496),
.B(n_5879),
.Y(n_6676)
);

NOR2xp33_ASAP7_75t_L g6677 ( 
.A(n_6190),
.B(n_5743),
.Y(n_6677)
);

AND2x2_ASAP7_75t_L g6678 ( 
.A(n_6384),
.B(n_6449),
.Y(n_6678)
);

INVx1_ASAP7_75t_L g6679 ( 
.A(n_6266),
.Y(n_6679)
);

OAI221xp5_ASAP7_75t_L g6680 ( 
.A1(n_6461),
.A2(n_5855),
.B1(n_5862),
.B2(n_5803),
.C(n_6073),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_6266),
.Y(n_6681)
);

INVxp33_ASAP7_75t_L g6682 ( 
.A(n_6308),
.Y(n_6682)
);

NAND2xp5_ASAP7_75t_SL g6683 ( 
.A(n_6482),
.B(n_5836),
.Y(n_6683)
);

NAND2xp5_ASAP7_75t_L g6684 ( 
.A(n_6388),
.B(n_6403),
.Y(n_6684)
);

NAND2xp5_ASAP7_75t_L g6685 ( 
.A(n_6375),
.B(n_5795),
.Y(n_6685)
);

INVx1_ASAP7_75t_L g6686 ( 
.A(n_6270),
.Y(n_6686)
);

NAND2xp5_ASAP7_75t_L g6687 ( 
.A(n_6237),
.B(n_5795),
.Y(n_6687)
);

NAND2xp5_ASAP7_75t_L g6688 ( 
.A(n_6247),
.B(n_5795),
.Y(n_6688)
);

BUFx3_ASAP7_75t_L g6689 ( 
.A(n_6219),
.Y(n_6689)
);

INVx1_ASAP7_75t_L g6690 ( 
.A(n_6270),
.Y(n_6690)
);

AND2x4_ASAP7_75t_L g6691 ( 
.A(n_6385),
.B(n_6065),
.Y(n_6691)
);

INVx1_ASAP7_75t_L g6692 ( 
.A(n_6282),
.Y(n_6692)
);

INVx2_ASAP7_75t_L g6693 ( 
.A(n_6486),
.Y(n_6693)
);

NAND2xp5_ASAP7_75t_L g6694 ( 
.A(n_6249),
.B(n_5795),
.Y(n_6694)
);

AND2x2_ASAP7_75t_L g6695 ( 
.A(n_6449),
.B(n_5811),
.Y(n_6695)
);

AND2x4_ASAP7_75t_L g6696 ( 
.A(n_6385),
.B(n_5691),
.Y(n_6696)
);

OR2x2_ASAP7_75t_L g6697 ( 
.A(n_6188),
.B(n_6023),
.Y(n_6697)
);

INVx2_ASAP7_75t_SL g6698 ( 
.A(n_6452),
.Y(n_6698)
);

NAND2xp5_ASAP7_75t_L g6699 ( 
.A(n_6415),
.B(n_5795),
.Y(n_6699)
);

NAND2xp5_ASAP7_75t_L g6700 ( 
.A(n_6452),
.B(n_6276),
.Y(n_6700)
);

INVx1_ASAP7_75t_L g6701 ( 
.A(n_6282),
.Y(n_6701)
);

INVx1_ASAP7_75t_L g6702 ( 
.A(n_6131),
.Y(n_6702)
);

OR2x2_ASAP7_75t_L g6703 ( 
.A(n_6188),
.B(n_5945),
.Y(n_6703)
);

NAND2xp5_ASAP7_75t_L g6704 ( 
.A(n_6276),
.B(n_5923),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_6153),
.Y(n_6705)
);

INVx2_ASAP7_75t_L g6706 ( 
.A(n_6486),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_6156),
.Y(n_6707)
);

AOI22xp33_ASAP7_75t_SL g6708 ( 
.A1(n_6340),
.A2(n_6055),
.B1(n_6114),
.B2(n_5840),
.Y(n_6708)
);

OR2x2_ASAP7_75t_L g6709 ( 
.A(n_6157),
.B(n_6081),
.Y(n_6709)
);

INVx2_ASAP7_75t_SL g6710 ( 
.A(n_6482),
.Y(n_6710)
);

BUFx6f_ASAP7_75t_L g6711 ( 
.A(n_6223),
.Y(n_6711)
);

INVx2_ASAP7_75t_L g6712 ( 
.A(n_6494),
.Y(n_6712)
);

INVxp67_ASAP7_75t_L g6713 ( 
.A(n_6343),
.Y(n_6713)
);

BUFx3_ASAP7_75t_L g6714 ( 
.A(n_6233),
.Y(n_6714)
);

INVx1_ASAP7_75t_L g6715 ( 
.A(n_6162),
.Y(n_6715)
);

BUFx2_ASAP7_75t_R g6716 ( 
.A(n_6233),
.Y(n_6716)
);

AND2x2_ASAP7_75t_L g6717 ( 
.A(n_6147),
.B(n_5949),
.Y(n_6717)
);

AND2x2_ASAP7_75t_L g6718 ( 
.A(n_6148),
.B(n_5950),
.Y(n_6718)
);

INVx2_ASAP7_75t_L g6719 ( 
.A(n_6494),
.Y(n_6719)
);

INVx2_ASAP7_75t_L g6720 ( 
.A(n_6504),
.Y(n_6720)
);

AND2x4_ASAP7_75t_SL g6721 ( 
.A(n_6359),
.B(n_5811),
.Y(n_6721)
);

INVx1_ASAP7_75t_SL g6722 ( 
.A(n_6210),
.Y(n_6722)
);

NAND2xp5_ASAP7_75t_L g6723 ( 
.A(n_6238),
.B(n_5923),
.Y(n_6723)
);

NAND2xp5_ASAP7_75t_L g6724 ( 
.A(n_6238),
.B(n_5885),
.Y(n_6724)
);

NAND2xp5_ASAP7_75t_L g6725 ( 
.A(n_6273),
.B(n_5902),
.Y(n_6725)
);

INVx1_ASAP7_75t_L g6726 ( 
.A(n_6164),
.Y(n_6726)
);

NAND2xp5_ASAP7_75t_L g6727 ( 
.A(n_6273),
.B(n_5902),
.Y(n_6727)
);

INVx1_ASAP7_75t_L g6728 ( 
.A(n_6297),
.Y(n_6728)
);

NAND2xp5_ASAP7_75t_L g6729 ( 
.A(n_6482),
.B(n_5902),
.Y(n_6729)
);

INVx4_ASAP7_75t_L g6730 ( 
.A(n_6223),
.Y(n_6730)
);

INVx2_ASAP7_75t_L g6731 ( 
.A(n_6504),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_6300),
.Y(n_6732)
);

AND4x1_ASAP7_75t_L g6733 ( 
.A(n_6472),
.B(n_6144),
.C(n_6453),
.D(n_6132),
.Y(n_6733)
);

HB1xp67_ASAP7_75t_L g6734 ( 
.A(n_6244),
.Y(n_6734)
);

INVx1_ASAP7_75t_L g6735 ( 
.A(n_6302),
.Y(n_6735)
);

INVx2_ASAP7_75t_L g6736 ( 
.A(n_6508),
.Y(n_6736)
);

NAND2xp5_ASAP7_75t_L g6737 ( 
.A(n_6482),
.B(n_5661),
.Y(n_6737)
);

INVx2_ASAP7_75t_L g6738 ( 
.A(n_6508),
.Y(n_6738)
);

AOI22xp5_ASAP7_75t_L g6739 ( 
.A1(n_6473),
.A2(n_6073),
.B1(n_5716),
.B2(n_5790),
.Y(n_6739)
);

INVx1_ASAP7_75t_L g6740 ( 
.A(n_6319),
.Y(n_6740)
);

AND2x2_ASAP7_75t_L g6741 ( 
.A(n_6148),
.B(n_5691),
.Y(n_6741)
);

AND2x2_ASAP7_75t_L g6742 ( 
.A(n_6503),
.B(n_5724),
.Y(n_6742)
);

AND2x2_ASAP7_75t_L g6743 ( 
.A(n_6503),
.B(n_6192),
.Y(n_6743)
);

AND2x2_ASAP7_75t_L g6744 ( 
.A(n_6503),
.B(n_5724),
.Y(n_6744)
);

INVx1_ASAP7_75t_L g6745 ( 
.A(n_6319),
.Y(n_6745)
);

INVx3_ASAP7_75t_L g6746 ( 
.A(n_6259),
.Y(n_6746)
);

HB1xp67_ASAP7_75t_L g6747 ( 
.A(n_6244),
.Y(n_6747)
);

INVx1_ASAP7_75t_L g6748 ( 
.A(n_6321),
.Y(n_6748)
);

AND2x2_ASAP7_75t_L g6749 ( 
.A(n_6503),
.B(n_5926),
.Y(n_6749)
);

AND2x2_ASAP7_75t_L g6750 ( 
.A(n_6192),
.B(n_5926),
.Y(n_6750)
);

BUFx2_ASAP7_75t_SL g6751 ( 
.A(n_6333),
.Y(n_6751)
);

INVx1_ASAP7_75t_L g6752 ( 
.A(n_6321),
.Y(n_6752)
);

INVx1_ASAP7_75t_L g6753 ( 
.A(n_6322),
.Y(n_6753)
);

INVx1_ASAP7_75t_L g6754 ( 
.A(n_6322),
.Y(n_6754)
);

INVx1_ASAP7_75t_L g6755 ( 
.A(n_6325),
.Y(n_6755)
);

NAND2xp5_ASAP7_75t_SL g6756 ( 
.A(n_6482),
.B(n_5836),
.Y(n_6756)
);

INVxp67_ASAP7_75t_SL g6757 ( 
.A(n_6495),
.Y(n_6757)
);

NAND2xp5_ASAP7_75t_L g6758 ( 
.A(n_6385),
.B(n_6304),
.Y(n_6758)
);

INVx1_ASAP7_75t_L g6759 ( 
.A(n_6325),
.Y(n_6759)
);

AND2x2_ASAP7_75t_L g6760 ( 
.A(n_6372),
.B(n_5915),
.Y(n_6760)
);

BUFx6f_ASAP7_75t_L g6761 ( 
.A(n_6223),
.Y(n_6761)
);

OR2x2_ASAP7_75t_L g6762 ( 
.A(n_6157),
.B(n_6085),
.Y(n_6762)
);

INVx2_ASAP7_75t_L g6763 ( 
.A(n_6509),
.Y(n_6763)
);

INVx1_ASAP7_75t_L g6764 ( 
.A(n_6326),
.Y(n_6764)
);

INVxp67_ASAP7_75t_SL g6765 ( 
.A(n_6495),
.Y(n_6765)
);

INVx2_ASAP7_75t_L g6766 ( 
.A(n_6509),
.Y(n_6766)
);

INVx1_ASAP7_75t_L g6767 ( 
.A(n_6326),
.Y(n_6767)
);

INVx2_ASAP7_75t_L g6768 ( 
.A(n_6402),
.Y(n_6768)
);

AND2x2_ASAP7_75t_L g6769 ( 
.A(n_6372),
.B(n_5917),
.Y(n_6769)
);

BUFx5_ASAP7_75t_L g6770 ( 
.A(n_6512),
.Y(n_6770)
);

NOR2x1_ASAP7_75t_SL g6771 ( 
.A(n_6359),
.B(n_5750),
.Y(n_6771)
);

INVx2_ASAP7_75t_L g6772 ( 
.A(n_6402),
.Y(n_6772)
);

OAI22xp5_ASAP7_75t_L g6773 ( 
.A1(n_6209),
.A2(n_6378),
.B1(n_6313),
.B2(n_5778),
.Y(n_6773)
);

INVx1_ASAP7_75t_L g6774 ( 
.A(n_6339),
.Y(n_6774)
);

OA21x2_ASAP7_75t_L g6775 ( 
.A1(n_6328),
.A2(n_5702),
.B(n_5675),
.Y(n_6775)
);

AND2x2_ASAP7_75t_L g6776 ( 
.A(n_6393),
.B(n_5745),
.Y(n_6776)
);

INVx1_ASAP7_75t_L g6777 ( 
.A(n_6339),
.Y(n_6777)
);

NOR2xp67_ASAP7_75t_L g6778 ( 
.A(n_6318),
.B(n_5801),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_6344),
.Y(n_6779)
);

INVx2_ASAP7_75t_L g6780 ( 
.A(n_6402),
.Y(n_6780)
);

AND2x2_ASAP7_75t_L g6781 ( 
.A(n_6393),
.B(n_5745),
.Y(n_6781)
);

OR2x2_ASAP7_75t_L g6782 ( 
.A(n_6180),
.B(n_6087),
.Y(n_6782)
);

AND2x2_ASAP7_75t_L g6783 ( 
.A(n_6399),
.B(n_5853),
.Y(n_6783)
);

BUFx2_ASAP7_75t_L g6784 ( 
.A(n_6454),
.Y(n_6784)
);

BUFx2_ASAP7_75t_L g6785 ( 
.A(n_6359),
.Y(n_6785)
);

AOI22xp33_ASAP7_75t_L g6786 ( 
.A1(n_6327),
.A2(n_4611),
.B1(n_4789),
.B2(n_5660),
.Y(n_6786)
);

AND2x2_ASAP7_75t_L g6787 ( 
.A(n_6198),
.B(n_5801),
.Y(n_6787)
);

BUFx12f_ASAP7_75t_L g6788 ( 
.A(n_6223),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_6344),
.Y(n_6789)
);

AND2x2_ASAP7_75t_L g6790 ( 
.A(n_6198),
.B(n_5802),
.Y(n_6790)
);

INVxp67_ASAP7_75t_L g6791 ( 
.A(n_6223),
.Y(n_6791)
);

NAND2xp5_ASAP7_75t_L g6792 ( 
.A(n_6305),
.B(n_5661),
.Y(n_6792)
);

INVx1_ASAP7_75t_L g6793 ( 
.A(n_6350),
.Y(n_6793)
);

AND2x2_ASAP7_75t_L g6794 ( 
.A(n_6453),
.B(n_5802),
.Y(n_6794)
);

AND2x2_ASAP7_75t_L g6795 ( 
.A(n_6152),
.B(n_5847),
.Y(n_6795)
);

HB1xp67_ASAP7_75t_L g6796 ( 
.A(n_6244),
.Y(n_6796)
);

OR2x2_ASAP7_75t_L g6797 ( 
.A(n_6180),
.B(n_6107),
.Y(n_6797)
);

AND2x2_ASAP7_75t_L g6798 ( 
.A(n_6152),
.B(n_5847),
.Y(n_6798)
);

AOI22xp5_ASAP7_75t_L g6799 ( 
.A1(n_6327),
.A2(n_6416),
.B1(n_6397),
.B2(n_6140),
.Y(n_6799)
);

AND2x4_ASAP7_75t_L g6800 ( 
.A(n_6359),
.B(n_5869),
.Y(n_6800)
);

OR2x2_ASAP7_75t_L g6801 ( 
.A(n_6239),
.B(n_6067),
.Y(n_6801)
);

NAND2xp5_ASAP7_75t_L g6802 ( 
.A(n_6306),
.B(n_5661),
.Y(n_6802)
);

AND2x2_ASAP7_75t_L g6803 ( 
.A(n_6155),
.B(n_5869),
.Y(n_6803)
);

AOI21xp33_ASAP7_75t_L g6804 ( 
.A1(n_6120),
.A2(n_5790),
.B(n_5911),
.Y(n_6804)
);

AND2x4_ASAP7_75t_L g6805 ( 
.A(n_6134),
.B(n_5954),
.Y(n_6805)
);

AND2x2_ASAP7_75t_L g6806 ( 
.A(n_6155),
.B(n_5954),
.Y(n_6806)
);

INVx2_ASAP7_75t_L g6807 ( 
.A(n_6435),
.Y(n_6807)
);

HB1xp67_ASAP7_75t_L g6808 ( 
.A(n_6483),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_6350),
.Y(n_6809)
);

AND2x2_ASAP7_75t_L g6810 ( 
.A(n_6399),
.B(n_5880),
.Y(n_6810)
);

INVx1_ASAP7_75t_L g6811 ( 
.A(n_6362),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_6362),
.Y(n_6812)
);

INVx1_ASAP7_75t_L g6813 ( 
.A(n_6364),
.Y(n_6813)
);

INVx1_ASAP7_75t_L g6814 ( 
.A(n_6364),
.Y(n_6814)
);

OR2x2_ASAP7_75t_L g6815 ( 
.A(n_6239),
.B(n_6108),
.Y(n_6815)
);

INVx2_ASAP7_75t_L g6816 ( 
.A(n_6435),
.Y(n_6816)
);

INVx1_ASAP7_75t_L g6817 ( 
.A(n_6391),
.Y(n_6817)
);

OR2x2_ASAP7_75t_L g6818 ( 
.A(n_6252),
.B(n_5788),
.Y(n_6818)
);

INVx2_ASAP7_75t_L g6819 ( 
.A(n_6435),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_6391),
.Y(n_6820)
);

NAND2xp5_ASAP7_75t_L g6821 ( 
.A(n_6307),
.B(n_5661),
.Y(n_6821)
);

AND2x2_ASAP7_75t_L g6822 ( 
.A(n_6429),
.B(n_5890),
.Y(n_6822)
);

INVx1_ASAP7_75t_L g6823 ( 
.A(n_6401),
.Y(n_6823)
);

OAI22xp5_ASAP7_75t_L g6824 ( 
.A1(n_6378),
.A2(n_6206),
.B1(n_6287),
.B2(n_6507),
.Y(n_6824)
);

INVx2_ASAP7_75t_SL g6825 ( 
.A(n_6512),
.Y(n_6825)
);

NOR2xp33_ASAP7_75t_L g6826 ( 
.A(n_6423),
.B(n_5881),
.Y(n_6826)
);

AND2x2_ASAP7_75t_L g6827 ( 
.A(n_6429),
.B(n_5960),
.Y(n_6827)
);

NAND2xp5_ASAP7_75t_L g6828 ( 
.A(n_6329),
.B(n_5861),
.Y(n_6828)
);

INVx2_ASAP7_75t_L g6829 ( 
.A(n_6279),
.Y(n_6829)
);

AOI22xp33_ASAP7_75t_L g6830 ( 
.A1(n_6170),
.A2(n_4611),
.B1(n_4789),
.B2(n_6027),
.Y(n_6830)
);

NOR2xp67_ASAP7_75t_L g6831 ( 
.A(n_6318),
.B(n_5968),
.Y(n_6831)
);

AND2x2_ASAP7_75t_L g6832 ( 
.A(n_6134),
.B(n_5887),
.Y(n_6832)
);

INVx2_ASAP7_75t_L g6833 ( 
.A(n_6279),
.Y(n_6833)
);

AND2x2_ASAP7_75t_L g6834 ( 
.A(n_6134),
.B(n_5895),
.Y(n_6834)
);

INVx1_ASAP7_75t_L g6835 ( 
.A(n_6401),
.Y(n_6835)
);

AND2x4_ASAP7_75t_L g6836 ( 
.A(n_6134),
.B(n_5968),
.Y(n_6836)
);

BUFx2_ASAP7_75t_L g6837 ( 
.A(n_6174),
.Y(n_6837)
);

AND2x2_ASAP7_75t_L g6838 ( 
.A(n_6165),
.B(n_5952),
.Y(n_6838)
);

NAND2xp5_ASAP7_75t_L g6839 ( 
.A(n_6361),
.B(n_6078),
.Y(n_6839)
);

BUFx3_ASAP7_75t_L g6840 ( 
.A(n_6467),
.Y(n_6840)
);

AND2x2_ASAP7_75t_L g6841 ( 
.A(n_6165),
.B(n_5958),
.Y(n_6841)
);

INVx1_ASAP7_75t_L g6842 ( 
.A(n_6406),
.Y(n_6842)
);

AND2x2_ASAP7_75t_L g6843 ( 
.A(n_6430),
.B(n_5967),
.Y(n_6843)
);

INVx2_ASAP7_75t_SL g6844 ( 
.A(n_6221),
.Y(n_6844)
);

AOI22xp33_ASAP7_75t_L g6845 ( 
.A1(n_6170),
.A2(n_4611),
.B1(n_4789),
.B2(n_6051),
.Y(n_6845)
);

AOI22xp33_ASAP7_75t_L g6846 ( 
.A1(n_6170),
.A2(n_4611),
.B1(n_4789),
.B2(n_5712),
.Y(n_6846)
);

INVxp67_ASAP7_75t_SL g6847 ( 
.A(n_6467),
.Y(n_6847)
);

NAND2xp5_ASAP7_75t_L g6848 ( 
.A(n_6371),
.B(n_6374),
.Y(n_6848)
);

AND2x2_ASAP7_75t_L g6849 ( 
.A(n_6430),
.B(n_5797),
.Y(n_6849)
);

HB1xp67_ASAP7_75t_L g6850 ( 
.A(n_6483),
.Y(n_6850)
);

NAND2x1_ASAP7_75t_L g6851 ( 
.A(n_6173),
.B(n_6060),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_6406),
.Y(n_6852)
);

AOI22xp33_ASAP7_75t_L g6853 ( 
.A1(n_6140),
.A2(n_4789),
.B1(n_5782),
.B2(n_5779),
.Y(n_6853)
);

INVx4_ASAP7_75t_L g6854 ( 
.A(n_6221),
.Y(n_6854)
);

NAND2x1p5_ASAP7_75t_L g6855 ( 
.A(n_6221),
.B(n_5669),
.Y(n_6855)
);

AND2x2_ASAP7_75t_L g6856 ( 
.A(n_6446),
.B(n_5970),
.Y(n_6856)
);

INVx1_ASAP7_75t_L g6857 ( 
.A(n_6408),
.Y(n_6857)
);

AND2x2_ASAP7_75t_L g6858 ( 
.A(n_6446),
.B(n_5985),
.Y(n_6858)
);

BUFx2_ASAP7_75t_L g6859 ( 
.A(n_6174),
.Y(n_6859)
);

AND2x2_ASAP7_75t_L g6860 ( 
.A(n_6234),
.B(n_6058),
.Y(n_6860)
);

INVx1_ASAP7_75t_L g6861 ( 
.A(n_6408),
.Y(n_6861)
);

NAND2xp5_ASAP7_75t_L g6862 ( 
.A(n_6379),
.B(n_5285),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_6410),
.Y(n_6863)
);

INVx1_ASAP7_75t_L g6864 ( 
.A(n_6410),
.Y(n_6864)
);

AOI22xp33_ASAP7_75t_L g6865 ( 
.A1(n_6140),
.A2(n_6014),
.B1(n_5538),
.B2(n_4801),
.Y(n_6865)
);

INVx1_ASAP7_75t_L g6866 ( 
.A(n_6412),
.Y(n_6866)
);

BUFx2_ASAP7_75t_L g6867 ( 
.A(n_6174),
.Y(n_6867)
);

OAI22xp5_ASAP7_75t_L g6868 ( 
.A1(n_6173),
.A2(n_5946),
.B1(n_5990),
.B2(n_5907),
.Y(n_6868)
);

OR2x2_ASAP7_75t_L g6869 ( 
.A(n_6252),
.B(n_5278),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_6412),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_6421),
.Y(n_6871)
);

INVx1_ASAP7_75t_L g6872 ( 
.A(n_6421),
.Y(n_6872)
);

BUFx3_ASAP7_75t_L g6873 ( 
.A(n_6221),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6425),
.Y(n_6874)
);

INVx1_ASAP7_75t_L g6875 ( 
.A(n_6425),
.Y(n_6875)
);

NAND2xp5_ASAP7_75t_L g6876 ( 
.A(n_6456),
.B(n_4638),
.Y(n_6876)
);

INVx1_ASAP7_75t_L g6877 ( 
.A(n_6431),
.Y(n_6877)
);

AOI22xp33_ASAP7_75t_L g6878 ( 
.A1(n_6341),
.A2(n_6120),
.B1(n_6253),
.B2(n_6200),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6431),
.Y(n_6879)
);

HB1xp67_ASAP7_75t_L g6880 ( 
.A(n_6483),
.Y(n_6880)
);

AND2x2_ASAP7_75t_L g6881 ( 
.A(n_6234),
.B(n_6059),
.Y(n_6881)
);

INVxp67_ASAP7_75t_L g6882 ( 
.A(n_6333),
.Y(n_6882)
);

AND2x2_ASAP7_75t_L g6883 ( 
.A(n_6284),
.B(n_6030),
.Y(n_6883)
);

NOR2xp33_ASAP7_75t_L g6884 ( 
.A(n_6221),
.B(n_5908),
.Y(n_6884)
);

BUFx3_ASAP7_75t_L g6885 ( 
.A(n_6311),
.Y(n_6885)
);

AND2x2_ASAP7_75t_L g6886 ( 
.A(n_6284),
.B(n_6033),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_6432),
.Y(n_6887)
);

OR2x2_ASAP7_75t_L g6888 ( 
.A(n_6280),
.B(n_5278),
.Y(n_6888)
);

AND2x4_ASAP7_75t_L g6889 ( 
.A(n_6387),
.B(n_5995),
.Y(n_6889)
);

INVxp67_ASAP7_75t_SL g6890 ( 
.A(n_6311),
.Y(n_6890)
);

INVx2_ASAP7_75t_L g6891 ( 
.A(n_6279),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_6432),
.Y(n_6892)
);

INVx2_ASAP7_75t_L g6893 ( 
.A(n_6396),
.Y(n_6893)
);

INVx1_ASAP7_75t_L g6894 ( 
.A(n_6434),
.Y(n_6894)
);

AND2x2_ASAP7_75t_L g6895 ( 
.A(n_6293),
.B(n_6041),
.Y(n_6895)
);

AND2x4_ASAP7_75t_L g6896 ( 
.A(n_6387),
.B(n_5995),
.Y(n_6896)
);

AOI22xp33_ASAP7_75t_L g6897 ( 
.A1(n_6341),
.A2(n_5538),
.B1(n_4801),
.B2(n_4701),
.Y(n_6897)
);

INVx2_ASAP7_75t_SL g6898 ( 
.A(n_6311),
.Y(n_6898)
);

INVx2_ASAP7_75t_L g6899 ( 
.A(n_6396),
.Y(n_6899)
);

BUFx2_ASAP7_75t_L g6900 ( 
.A(n_6784),
.Y(n_6900)
);

AND2x2_ASAP7_75t_L g6901 ( 
.A(n_6678),
.B(n_6498),
.Y(n_6901)
);

AND2x2_ASAP7_75t_L g6902 ( 
.A(n_6543),
.B(n_6498),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6551),
.Y(n_6903)
);

INVx3_ASAP7_75t_L g6904 ( 
.A(n_6851),
.Y(n_6904)
);

AND2x4_ASAP7_75t_SL g6905 ( 
.A(n_6528),
.B(n_6311),
.Y(n_6905)
);

NAND2xp5_ASAP7_75t_L g6906 ( 
.A(n_6722),
.B(n_6434),
.Y(n_6906)
);

INVx2_ASAP7_75t_L g6907 ( 
.A(n_6527),
.Y(n_6907)
);

AOI221xp5_ASAP7_75t_L g6908 ( 
.A1(n_6564),
.A2(n_6246),
.B1(n_6400),
.B2(n_6184),
.C(n_6178),
.Y(n_6908)
);

AND2x2_ASAP7_75t_L g6909 ( 
.A(n_6543),
.B(n_6275),
.Y(n_6909)
);

NOR2x1_ASAP7_75t_L g6910 ( 
.A(n_6730),
.B(n_6268),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_6551),
.Y(n_6911)
);

INVx1_ASAP7_75t_L g6912 ( 
.A(n_6556),
.Y(n_6912)
);

OR2x2_ASAP7_75t_L g6913 ( 
.A(n_6618),
.B(n_6283),
.Y(n_6913)
);

NAND2xp5_ASAP7_75t_L g6914 ( 
.A(n_6564),
.B(n_6436),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_6556),
.Y(n_6915)
);

HB1xp67_ASAP7_75t_L g6916 ( 
.A(n_6605),
.Y(n_6916)
);

INVx1_ASAP7_75t_L g6917 ( 
.A(n_6557),
.Y(n_6917)
);

NOR2x1_ASAP7_75t_L g6918 ( 
.A(n_6730),
.B(n_6854),
.Y(n_6918)
);

NAND2x1_ASAP7_75t_L g6919 ( 
.A(n_6629),
.B(n_6318),
.Y(n_6919)
);

AND2x2_ASAP7_75t_L g6920 ( 
.A(n_6538),
.B(n_6275),
.Y(n_6920)
);

INVx2_ASAP7_75t_L g6921 ( 
.A(n_6527),
.Y(n_6921)
);

AND2x2_ASAP7_75t_L g6922 ( 
.A(n_6538),
.B(n_6311),
.Y(n_6922)
);

HB1xp67_ASAP7_75t_L g6923 ( 
.A(n_6605),
.Y(n_6923)
);

AND2x4_ASAP7_75t_L g6924 ( 
.A(n_6639),
.B(n_6290),
.Y(n_6924)
);

AND2x2_ASAP7_75t_L g6925 ( 
.A(n_6549),
.B(n_6293),
.Y(n_6925)
);

INVx2_ASAP7_75t_L g6926 ( 
.A(n_6527),
.Y(n_6926)
);

INVx2_ASAP7_75t_L g6927 ( 
.A(n_6672),
.Y(n_6927)
);

INVx2_ASAP7_75t_SL g6928 ( 
.A(n_6628),
.Y(n_6928)
);

AND2x2_ASAP7_75t_L g6929 ( 
.A(n_6549),
.B(n_6295),
.Y(n_6929)
);

AND2x2_ASAP7_75t_L g6930 ( 
.A(n_6523),
.B(n_5797),
.Y(n_6930)
);

INVx1_ASAP7_75t_L g6931 ( 
.A(n_6557),
.Y(n_6931)
);

AND2x2_ASAP7_75t_L g6932 ( 
.A(n_6560),
.B(n_5809),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_6565),
.Y(n_6933)
);

AO21x2_ASAP7_75t_L g6934 ( 
.A1(n_6808),
.A2(n_6511),
.B(n_6464),
.Y(n_6934)
);

AND2x2_ASAP7_75t_L g6935 ( 
.A(n_6589),
.B(n_5809),
.Y(n_6935)
);

BUFx5_ASAP7_75t_L g6936 ( 
.A(n_6788),
.Y(n_6936)
);

NAND3xp33_ASAP7_75t_L g6937 ( 
.A(n_6540),
.B(n_6390),
.C(n_6511),
.Y(n_6937)
);

AND2x2_ASAP7_75t_L g6938 ( 
.A(n_6646),
.B(n_6360),
.Y(n_6938)
);

OR2x2_ASAP7_75t_L g6939 ( 
.A(n_6573),
.B(n_6283),
.Y(n_6939)
);

INVx2_ASAP7_75t_L g6940 ( 
.A(n_6672),
.Y(n_6940)
);

AND2x2_ASAP7_75t_L g6941 ( 
.A(n_6827),
.B(n_6360),
.Y(n_6941)
);

INVx2_ASAP7_75t_SL g6942 ( 
.A(n_6628),
.Y(n_6942)
);

INVx2_ASAP7_75t_L g6943 ( 
.A(n_6672),
.Y(n_6943)
);

AO21x2_ASAP7_75t_L g6944 ( 
.A1(n_6808),
.A2(n_6464),
.B(n_6462),
.Y(n_6944)
);

INVxp67_ASAP7_75t_SL g6945 ( 
.A(n_6516),
.Y(n_6945)
);

INVx2_ASAP7_75t_L g6946 ( 
.A(n_6746),
.Y(n_6946)
);

INVx2_ASAP7_75t_L g6947 ( 
.A(n_6746),
.Y(n_6947)
);

INVx2_ASAP7_75t_L g6948 ( 
.A(n_6746),
.Y(n_6948)
);

INVx1_ASAP7_75t_L g6949 ( 
.A(n_6565),
.Y(n_6949)
);

INVx3_ASAP7_75t_L g6950 ( 
.A(n_6608),
.Y(n_6950)
);

HB1xp67_ASAP7_75t_L g6951 ( 
.A(n_6608),
.Y(n_6951)
);

INVx2_ASAP7_75t_L g6952 ( 
.A(n_6533),
.Y(n_6952)
);

NOR2x1_ASAP7_75t_L g6953 ( 
.A(n_6730),
.B(n_6411),
.Y(n_6953)
);

INVx2_ASAP7_75t_SL g6954 ( 
.A(n_6711),
.Y(n_6954)
);

AND2x2_ASAP7_75t_L g6955 ( 
.A(n_6664),
.B(n_6860),
.Y(n_6955)
);

INVx5_ASAP7_75t_L g6956 ( 
.A(n_6568),
.Y(n_6956)
);

OR2x2_ASAP7_75t_L g6957 ( 
.A(n_6640),
.B(n_6280),
.Y(n_6957)
);

HB1xp67_ASAP7_75t_L g6958 ( 
.A(n_6620),
.Y(n_6958)
);

NAND2xp5_ASAP7_75t_L g6959 ( 
.A(n_6537),
.B(n_6436),
.Y(n_6959)
);

AND2x4_ASAP7_75t_L g6960 ( 
.A(n_6639),
.B(n_6290),
.Y(n_6960)
);

INVx2_ASAP7_75t_SL g6961 ( 
.A(n_6711),
.Y(n_6961)
);

NAND2xp5_ASAP7_75t_L g6962 ( 
.A(n_6546),
.B(n_6439),
.Y(n_6962)
);

NAND2xp5_ASAP7_75t_L g6963 ( 
.A(n_6569),
.B(n_6439),
.Y(n_6963)
);

BUFx3_ASAP7_75t_L g6964 ( 
.A(n_6689),
.Y(n_6964)
);

INVx1_ASAP7_75t_L g6965 ( 
.A(n_6620),
.Y(n_6965)
);

AND2x4_ASAP7_75t_L g6966 ( 
.A(n_6639),
.B(n_6387),
.Y(n_6966)
);

AND2x2_ASAP7_75t_L g6967 ( 
.A(n_6860),
.B(n_6295),
.Y(n_6967)
);

INVx3_ASAP7_75t_L g6968 ( 
.A(n_6788),
.Y(n_6968)
);

HB1xp67_ASAP7_75t_L g6969 ( 
.A(n_6643),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6643),
.Y(n_6970)
);

HB1xp67_ASAP7_75t_L g6971 ( 
.A(n_6734),
.Y(n_6971)
);

AND2x2_ASAP7_75t_L g6972 ( 
.A(n_6881),
.B(n_6381),
.Y(n_6972)
);

OAI321xp33_ASAP7_75t_L g6973 ( 
.A1(n_6574),
.A2(n_6146),
.A3(n_6232),
.B1(n_6314),
.B2(n_6336),
.C(n_6474),
.Y(n_6973)
);

NAND2x1_ASAP7_75t_L g6974 ( 
.A(n_6629),
.B(n_6411),
.Y(n_6974)
);

INVx1_ASAP7_75t_L g6975 ( 
.A(n_6734),
.Y(n_6975)
);

OR2x2_ASAP7_75t_L g6976 ( 
.A(n_6520),
.B(n_6443),
.Y(n_6976)
);

INVx1_ASAP7_75t_L g6977 ( 
.A(n_6747),
.Y(n_6977)
);

AND2x2_ASAP7_75t_L g6978 ( 
.A(n_6881),
.B(n_6381),
.Y(n_6978)
);

AOI21xp5_ASAP7_75t_L g6979 ( 
.A1(n_6574),
.A2(n_6079),
.B(n_6228),
.Y(n_6979)
);

INVx2_ASAP7_75t_L g6980 ( 
.A(n_6533),
.Y(n_6980)
);

INVx1_ASAP7_75t_L g6981 ( 
.A(n_6747),
.Y(n_6981)
);

BUFx3_ASAP7_75t_L g6982 ( 
.A(n_6689),
.Y(n_6982)
);

OR2x2_ASAP7_75t_L g6983 ( 
.A(n_6522),
.B(n_6443),
.Y(n_6983)
);

AND2x2_ASAP7_75t_L g6984 ( 
.A(n_6555),
.B(n_6366),
.Y(n_6984)
);

INVx1_ASAP7_75t_L g6985 ( 
.A(n_6796),
.Y(n_6985)
);

AND2x2_ASAP7_75t_L g6986 ( 
.A(n_6750),
.B(n_6366),
.Y(n_6986)
);

HB1xp67_ASAP7_75t_L g6987 ( 
.A(n_6796),
.Y(n_6987)
);

HB1xp67_ASAP7_75t_L g6988 ( 
.A(n_6850),
.Y(n_6988)
);

AND2x2_ASAP7_75t_L g6989 ( 
.A(n_6750),
.B(n_6757),
.Y(n_6989)
);

BUFx3_ASAP7_75t_L g6990 ( 
.A(n_6568),
.Y(n_6990)
);

INVx1_ASAP7_75t_L g6991 ( 
.A(n_6850),
.Y(n_6991)
);

AND2x4_ASAP7_75t_SL g6992 ( 
.A(n_6528),
.B(n_6381),
.Y(n_6992)
);

BUFx2_ASAP7_75t_L g6993 ( 
.A(n_6714),
.Y(n_6993)
);

AND2x2_ASAP7_75t_L g6994 ( 
.A(n_6765),
.B(n_6471),
.Y(n_6994)
);

INVx2_ASAP7_75t_L g6995 ( 
.A(n_6539),
.Y(n_6995)
);

OR2x2_ASAP7_75t_L g6996 ( 
.A(n_6535),
.B(n_6444),
.Y(n_6996)
);

OA21x2_ASAP7_75t_L g6997 ( 
.A1(n_6878),
.A2(n_6328),
.B(n_6323),
.Y(n_6997)
);

AO21x2_ASAP7_75t_L g6998 ( 
.A1(n_6880),
.A2(n_6470),
.B(n_6462),
.Y(n_6998)
);

INVx1_ASAP7_75t_L g6999 ( 
.A(n_6880),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6519),
.Y(n_7000)
);

INVx2_ASAP7_75t_L g7001 ( 
.A(n_6539),
.Y(n_7001)
);

HB1xp67_ASAP7_75t_L g7002 ( 
.A(n_6572),
.Y(n_7002)
);

INVx2_ASAP7_75t_L g7003 ( 
.A(n_6548),
.Y(n_7003)
);

INVx2_ASAP7_75t_L g7004 ( 
.A(n_6548),
.Y(n_7004)
);

INVx1_ASAP7_75t_L g7005 ( 
.A(n_6519),
.Y(n_7005)
);

AND2x2_ASAP7_75t_L g7006 ( 
.A(n_6600),
.B(n_6438),
.Y(n_7006)
);

INVx1_ASAP7_75t_SL g7007 ( 
.A(n_6716),
.Y(n_7007)
);

NAND3xp33_ASAP7_75t_L g7008 ( 
.A(n_6540),
.B(n_6120),
.C(n_6253),
.Y(n_7008)
);

BUFx6f_ASAP7_75t_L g7009 ( 
.A(n_6568),
.Y(n_7009)
);

HB1xp67_ASAP7_75t_L g7010 ( 
.A(n_6609),
.Y(n_7010)
);

INVx1_ASAP7_75t_L g7011 ( 
.A(n_6521),
.Y(n_7011)
);

AND2x2_ASAP7_75t_L g7012 ( 
.A(n_6612),
.B(n_6438),
.Y(n_7012)
);

INVx1_ASAP7_75t_L g7013 ( 
.A(n_6521),
.Y(n_7013)
);

AND2x2_ASAP7_75t_L g7014 ( 
.A(n_6619),
.B(n_6438),
.Y(n_7014)
);

BUFx2_ASAP7_75t_L g7015 ( 
.A(n_6714),
.Y(n_7015)
);

AND2x2_ASAP7_75t_L g7016 ( 
.A(n_6670),
.B(n_6471),
.Y(n_7016)
);

INVx2_ASAP7_75t_L g7017 ( 
.A(n_6526),
.Y(n_7017)
);

AND2x2_ASAP7_75t_L g7018 ( 
.A(n_6671),
.B(n_6224),
.Y(n_7018)
);

AOI22xp33_ASAP7_75t_L g7019 ( 
.A1(n_6878),
.A2(n_6680),
.B1(n_6804),
.B2(n_6659),
.Y(n_7019)
);

INVx1_ASAP7_75t_L g7020 ( 
.A(n_6526),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6740),
.Y(n_7021)
);

NAND2xp5_ASAP7_75t_SL g7022 ( 
.A(n_6733),
.B(n_5783),
.Y(n_7022)
);

NOR2x1_ASAP7_75t_L g7023 ( 
.A(n_6854),
.B(n_6010),
.Y(n_7023)
);

BUFx2_ASAP7_75t_L g7024 ( 
.A(n_6840),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6745),
.Y(n_7025)
);

INVx1_ASAP7_75t_L g7026 ( 
.A(n_6748),
.Y(n_7026)
);

AND2x4_ASAP7_75t_L g7027 ( 
.A(n_6616),
.B(n_6392),
.Y(n_7027)
);

AOI22xp33_ASAP7_75t_L g7028 ( 
.A1(n_6659),
.A2(n_6341),
.B1(n_6120),
.B2(n_6253),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6752),
.Y(n_7029)
);

INVx1_ASAP7_75t_L g7030 ( 
.A(n_6753),
.Y(n_7030)
);

INVx1_ASAP7_75t_L g7031 ( 
.A(n_6754),
.Y(n_7031)
);

AOI22xp33_ASAP7_75t_L g7032 ( 
.A1(n_6799),
.A2(n_6341),
.B1(n_6253),
.B2(n_6335),
.Y(n_7032)
);

AOI321xp33_ASAP7_75t_L g7033 ( 
.A1(n_6824),
.A2(n_6465),
.A3(n_6470),
.B1(n_6478),
.B2(n_6497),
.C(n_6485),
.Y(n_7033)
);

BUFx6f_ASAP7_75t_L g7034 ( 
.A(n_6568),
.Y(n_7034)
);

HB1xp67_ASAP7_75t_L g7035 ( 
.A(n_6611),
.Y(n_7035)
);

OR2x2_ASAP7_75t_L g7036 ( 
.A(n_6530),
.B(n_6444),
.Y(n_7036)
);

AND2x2_ASAP7_75t_L g7037 ( 
.A(n_6838),
.B(n_6224),
.Y(n_7037)
);

AND2x2_ASAP7_75t_L g7038 ( 
.A(n_6838),
.B(n_6225),
.Y(n_7038)
);

AND2x2_ASAP7_75t_L g7039 ( 
.A(n_6841),
.B(n_6225),
.Y(n_7039)
);

AND2x4_ASAP7_75t_L g7040 ( 
.A(n_6669),
.B(n_6392),
.Y(n_7040)
);

INVx2_ASAP7_75t_L g7041 ( 
.A(n_6829),
.Y(n_7041)
);

INVx1_ASAP7_75t_L g7042 ( 
.A(n_6755),
.Y(n_7042)
);

INVx1_ASAP7_75t_L g7043 ( 
.A(n_6759),
.Y(n_7043)
);

NOR2xp33_ASAP7_75t_SL g7044 ( 
.A(n_6516),
.B(n_6333),
.Y(n_7044)
);

INVx2_ASAP7_75t_L g7045 ( 
.A(n_6829),
.Y(n_7045)
);

AOI22xp33_ASAP7_75t_L g7046 ( 
.A1(n_6675),
.A2(n_6335),
.B1(n_6396),
.B2(n_6465),
.Y(n_7046)
);

AND2x2_ASAP7_75t_L g7047 ( 
.A(n_6841),
.B(n_5783),
.Y(n_7047)
);

AND2x2_ASAP7_75t_L g7048 ( 
.A(n_6847),
.B(n_6407),
.Y(n_7048)
);

OR2x2_ASAP7_75t_L g7049 ( 
.A(n_6532),
.B(n_6445),
.Y(n_7049)
);

INVx1_ASAP7_75t_SL g7050 ( 
.A(n_6592),
.Y(n_7050)
);

AND2x2_ASAP7_75t_L g7051 ( 
.A(n_6559),
.B(n_6547),
.Y(n_7051)
);

INVx5_ASAP7_75t_SL g7052 ( 
.A(n_6585),
.Y(n_7052)
);

INVx1_ASAP7_75t_SL g7053 ( 
.A(n_6592),
.Y(n_7053)
);

HB1xp67_ASAP7_75t_L g7054 ( 
.A(n_6668),
.Y(n_7054)
);

OR2x2_ASAP7_75t_L g7055 ( 
.A(n_6583),
.B(n_6445),
.Y(n_7055)
);

HB1xp67_ASAP7_75t_L g7056 ( 
.A(n_6558),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_6764),
.Y(n_7057)
);

AND2x4_ASAP7_75t_L g7058 ( 
.A(n_6629),
.B(n_6392),
.Y(n_7058)
);

INVx2_ASAP7_75t_L g7059 ( 
.A(n_6833),
.Y(n_7059)
);

AOI22xp33_ASAP7_75t_L g7060 ( 
.A1(n_6739),
.A2(n_6335),
.B1(n_6256),
.B2(n_6441),
.Y(n_7060)
);

AND2x2_ASAP7_75t_L g7061 ( 
.A(n_6559),
.B(n_6049),
.Y(n_7061)
);

BUFx2_ASAP7_75t_L g7062 ( 
.A(n_6840),
.Y(n_7062)
);

AND2x4_ASAP7_75t_L g7063 ( 
.A(n_6698),
.B(n_6427),
.Y(n_7063)
);

AND2x2_ASAP7_75t_L g7064 ( 
.A(n_6547),
.B(n_6424),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_6767),
.Y(n_7065)
);

INVx1_ASAP7_75t_L g7066 ( 
.A(n_6774),
.Y(n_7066)
);

AND2x2_ASAP7_75t_L g7067 ( 
.A(n_6743),
.B(n_6489),
.Y(n_7067)
);

INVxp67_ASAP7_75t_SL g7068 ( 
.A(n_6633),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_6777),
.Y(n_7069)
);

OR2x2_ASAP7_75t_L g7070 ( 
.A(n_6614),
.B(n_6460),
.Y(n_7070)
);

NAND2xp5_ASAP7_75t_L g7071 ( 
.A(n_6698),
.B(n_6460),
.Y(n_7071)
);

INVx2_ASAP7_75t_L g7072 ( 
.A(n_6833),
.Y(n_7072)
);

NAND2xp5_ASAP7_75t_L g7073 ( 
.A(n_6544),
.B(n_6441),
.Y(n_7073)
);

OR2x2_ASAP7_75t_L g7074 ( 
.A(n_6818),
.B(n_6484),
.Y(n_7074)
);

NAND2xp5_ASAP7_75t_L g7075 ( 
.A(n_6544),
.B(n_6463),
.Y(n_7075)
);

AND2x2_ASAP7_75t_L g7076 ( 
.A(n_6743),
.B(n_6489),
.Y(n_7076)
);

NOR2xp33_ASAP7_75t_L g7077 ( 
.A(n_6552),
.B(n_6370),
.Y(n_7077)
);

BUFx2_ASAP7_75t_L g7078 ( 
.A(n_6517),
.Y(n_7078)
);

AND2x2_ASAP7_75t_L g7079 ( 
.A(n_6517),
.B(n_6493),
.Y(n_7079)
);

BUFx3_ASAP7_75t_L g7080 ( 
.A(n_6585),
.Y(n_7080)
);

INVx5_ASAP7_75t_SL g7081 ( 
.A(n_6585),
.Y(n_7081)
);

INVx5_ASAP7_75t_L g7082 ( 
.A(n_6585),
.Y(n_7082)
);

AND2x4_ASAP7_75t_L g7083 ( 
.A(n_6528),
.B(n_6427),
.Y(n_7083)
);

AND2x2_ASAP7_75t_L g7084 ( 
.A(n_6517),
.B(n_6749),
.Y(n_7084)
);

AOI22xp33_ASAP7_75t_L g7085 ( 
.A1(n_6724),
.A2(n_6335),
.B1(n_6256),
.B2(n_6463),
.Y(n_7085)
);

INVx1_ASAP7_75t_L g7086 ( 
.A(n_6779),
.Y(n_7086)
);

INVxp67_ASAP7_75t_SL g7087 ( 
.A(n_6633),
.Y(n_7087)
);

INVx2_ASAP7_75t_L g7088 ( 
.A(n_6891),
.Y(n_7088)
);

INVx2_ASAP7_75t_L g7089 ( 
.A(n_6891),
.Y(n_7089)
);

NAND2xp5_ASAP7_75t_L g7090 ( 
.A(n_6783),
.B(n_6810),
.Y(n_7090)
);

INVx3_ASAP7_75t_L g7091 ( 
.A(n_6711),
.Y(n_7091)
);

AND2x2_ASAP7_75t_L g7092 ( 
.A(n_6749),
.B(n_6424),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6789),
.Y(n_7093)
);

AND2x2_ASAP7_75t_L g7094 ( 
.A(n_6751),
.B(n_6426),
.Y(n_7094)
);

INVxp67_ASAP7_75t_SL g7095 ( 
.A(n_6529),
.Y(n_7095)
);

INVx1_ASAP7_75t_L g7096 ( 
.A(n_6793),
.Y(n_7096)
);

HB1xp67_ASAP7_75t_L g7097 ( 
.A(n_6562),
.Y(n_7097)
);

HB1xp67_ASAP7_75t_L g7098 ( 
.A(n_6725),
.Y(n_7098)
);

NOR2xp33_ASAP7_75t_L g7099 ( 
.A(n_6552),
.B(n_6433),
.Y(n_7099)
);

INVx2_ASAP7_75t_L g7100 ( 
.A(n_6893),
.Y(n_7100)
);

NAND2xp5_ASAP7_75t_L g7101 ( 
.A(n_6822),
.B(n_6332),
.Y(n_7101)
);

AND2x2_ASAP7_75t_L g7102 ( 
.A(n_6741),
.B(n_6426),
.Y(n_7102)
);

OR2x2_ASAP7_75t_L g7103 ( 
.A(n_6666),
.B(n_6422),
.Y(n_7103)
);

AND2x2_ASAP7_75t_L g7104 ( 
.A(n_6741),
.B(n_6447),
.Y(n_7104)
);

INVx2_ASAP7_75t_L g7105 ( 
.A(n_6893),
.Y(n_7105)
);

INVx2_ASAP7_75t_L g7106 ( 
.A(n_6899),
.Y(n_7106)
);

BUFx3_ASAP7_75t_L g7107 ( 
.A(n_6770),
.Y(n_7107)
);

INVx3_ASAP7_75t_L g7108 ( 
.A(n_6711),
.Y(n_7108)
);

NAND2xp5_ASAP7_75t_L g7109 ( 
.A(n_6791),
.B(n_6514),
.Y(n_7109)
);

BUFx2_ASAP7_75t_L g7110 ( 
.A(n_6761),
.Y(n_7110)
);

AND2x2_ASAP7_75t_L g7111 ( 
.A(n_6795),
.B(n_6447),
.Y(n_7111)
);

AND2x4_ASAP7_75t_L g7112 ( 
.A(n_6761),
.B(n_6885),
.Y(n_7112)
);

HB1xp67_ASAP7_75t_L g7113 ( 
.A(n_6727),
.Y(n_7113)
);

INVx3_ASAP7_75t_L g7114 ( 
.A(n_6761),
.Y(n_7114)
);

INVx1_ASAP7_75t_L g7115 ( 
.A(n_6809),
.Y(n_7115)
);

INVx1_ASAP7_75t_L g7116 ( 
.A(n_6811),
.Y(n_7116)
);

INVx2_ASAP7_75t_L g7117 ( 
.A(n_6899),
.Y(n_7117)
);

INVx2_ASAP7_75t_L g7118 ( 
.A(n_6768),
.Y(n_7118)
);

INVx1_ASAP7_75t_L g7119 ( 
.A(n_6812),
.Y(n_7119)
);

AND2x2_ASAP7_75t_L g7120 ( 
.A(n_6883),
.B(n_6795),
.Y(n_7120)
);

INVxp67_ASAP7_75t_L g7121 ( 
.A(n_6601),
.Y(n_7121)
);

INVx1_ASAP7_75t_L g7122 ( 
.A(n_6813),
.Y(n_7122)
);

BUFx2_ASAP7_75t_L g7123 ( 
.A(n_6761),
.Y(n_7123)
);

INVx1_ASAP7_75t_L g7124 ( 
.A(n_6814),
.Y(n_7124)
);

INVx1_ASAP7_75t_L g7125 ( 
.A(n_6817),
.Y(n_7125)
);

HB1xp67_ASAP7_75t_L g7126 ( 
.A(n_6684),
.Y(n_7126)
);

INVx2_ASAP7_75t_L g7127 ( 
.A(n_6768),
.Y(n_7127)
);

AND2x2_ASAP7_75t_L g7128 ( 
.A(n_6883),
.B(n_6493),
.Y(n_7128)
);

NAND2xp5_ASAP7_75t_L g7129 ( 
.A(n_6760),
.B(n_6514),
.Y(n_7129)
);

AND2x2_ASAP7_75t_L g7130 ( 
.A(n_6798),
.B(n_6409),
.Y(n_7130)
);

INVx3_ASAP7_75t_L g7131 ( 
.A(n_6552),
.Y(n_7131)
);

INVx2_ASAP7_75t_SL g7132 ( 
.A(n_6648),
.Y(n_7132)
);

NOR2x1_ASAP7_75t_L g7133 ( 
.A(n_6854),
.B(n_6010),
.Y(n_7133)
);

NAND2xp5_ASAP7_75t_L g7134 ( 
.A(n_6769),
.B(n_6514),
.Y(n_7134)
);

AND2x2_ASAP7_75t_L g7135 ( 
.A(n_6798),
.B(n_6409),
.Y(n_7135)
);

BUFx2_ASAP7_75t_L g7136 ( 
.A(n_6889),
.Y(n_7136)
);

AND2x2_ASAP7_75t_L g7137 ( 
.A(n_6803),
.B(n_6016),
.Y(n_7137)
);

NAND2xp5_ASAP7_75t_L g7138 ( 
.A(n_6825),
.B(n_6455),
.Y(n_7138)
);

INVx4_ASAP7_75t_L g7139 ( 
.A(n_6885),
.Y(n_7139)
);

INVx4_ASAP7_75t_L g7140 ( 
.A(n_6873),
.Y(n_7140)
);

AND2x4_ASAP7_75t_L g7141 ( 
.A(n_6825),
.B(n_6427),
.Y(n_7141)
);

INVx1_ASAP7_75t_L g7142 ( 
.A(n_6820),
.Y(n_7142)
);

INVx2_ASAP7_75t_L g7143 ( 
.A(n_6772),
.Y(n_7143)
);

AND2x2_ASAP7_75t_L g7144 ( 
.A(n_6803),
.B(n_6806),
.Y(n_7144)
);

AND2x4_ASAP7_75t_L g7145 ( 
.A(n_6800),
.B(n_6124),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_6823),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_6835),
.Y(n_7147)
);

INVx2_ASAP7_75t_L g7148 ( 
.A(n_6772),
.Y(n_7148)
);

NOR2xp33_ASAP7_75t_L g7149 ( 
.A(n_6601),
.B(n_6433),
.Y(n_7149)
);

INVx1_ASAP7_75t_L g7150 ( 
.A(n_6842),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_6852),
.Y(n_7151)
);

OR2x2_ASAP7_75t_L g7152 ( 
.A(n_6697),
.B(n_6762),
.Y(n_7152)
);

AND2x2_ASAP7_75t_L g7153 ( 
.A(n_6806),
.B(n_6016),
.Y(n_7153)
);

AND2x2_ASAP7_75t_L g7154 ( 
.A(n_6623),
.B(n_5994),
.Y(n_7154)
);

INVx1_ASAP7_75t_L g7155 ( 
.A(n_6857),
.Y(n_7155)
);

AND2x2_ASAP7_75t_L g7156 ( 
.A(n_6623),
.B(n_5998),
.Y(n_7156)
);

NAND2x1p5_ASAP7_75t_L g7157 ( 
.A(n_6683),
.B(n_6756),
.Y(n_7157)
);

INVx1_ASAP7_75t_L g7158 ( 
.A(n_6861),
.Y(n_7158)
);

NAND2xp5_ASAP7_75t_L g7159 ( 
.A(n_6571),
.B(n_6455),
.Y(n_7159)
);

AND2x4_ASAP7_75t_L g7160 ( 
.A(n_6800),
.B(n_6124),
.Y(n_7160)
);

AND2x2_ASAP7_75t_L g7161 ( 
.A(n_6673),
.B(n_6011),
.Y(n_7161)
);

BUFx2_ASAP7_75t_L g7162 ( 
.A(n_6889),
.Y(n_7162)
);

AND2x4_ASAP7_75t_L g7163 ( 
.A(n_6800),
.B(n_6124),
.Y(n_7163)
);

BUFx2_ASAP7_75t_L g7164 ( 
.A(n_6889),
.Y(n_7164)
);

AND2x2_ASAP7_75t_L g7165 ( 
.A(n_6676),
.B(n_6017),
.Y(n_7165)
);

HB1xp67_ASAP7_75t_L g7166 ( 
.A(n_6737),
.Y(n_7166)
);

NAND4xp25_ASAP7_75t_L g7167 ( 
.A(n_6773),
.B(n_6500),
.C(n_5720),
.D(n_6294),
.Y(n_7167)
);

AOI22xp33_ASAP7_75t_L g7168 ( 
.A1(n_6662),
.A2(n_6256),
.B1(n_6259),
.B2(n_6258),
.Y(n_7168)
);

INVx2_ASAP7_75t_L g7169 ( 
.A(n_6780),
.Y(n_7169)
);

HB1xp67_ASAP7_75t_L g7170 ( 
.A(n_6625),
.Y(n_7170)
);

INVxp67_ASAP7_75t_SL g7171 ( 
.A(n_6713),
.Y(n_7171)
);

AND2x4_ASAP7_75t_L g7172 ( 
.A(n_6778),
.B(n_6124),
.Y(n_7172)
);

INVx1_ASAP7_75t_L g7173 ( 
.A(n_6863),
.Y(n_7173)
);

INVx5_ASAP7_75t_L g7174 ( 
.A(n_6844),
.Y(n_7174)
);

NAND2xp5_ASAP7_75t_L g7175 ( 
.A(n_6638),
.B(n_6455),
.Y(n_7175)
);

OAI33xp33_ASAP7_75t_L g7176 ( 
.A1(n_6792),
.A2(n_6422),
.A3(n_6428),
.B1(n_6358),
.B2(n_6485),
.B3(n_6478),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_6864),
.Y(n_7177)
);

BUFx3_ASAP7_75t_L g7178 ( 
.A(n_6770),
.Y(n_7178)
);

INVx1_ASAP7_75t_L g7179 ( 
.A(n_6866),
.Y(n_7179)
);

AND2x4_ASAP7_75t_L g7180 ( 
.A(n_6831),
.B(n_6160),
.Y(n_7180)
);

BUFx3_ASAP7_75t_L g7181 ( 
.A(n_6770),
.Y(n_7181)
);

NOR2x1_ASAP7_75t_SL g7182 ( 
.A(n_6683),
.B(n_6299),
.Y(n_7182)
);

AND2x2_ASAP7_75t_L g7183 ( 
.A(n_6658),
.B(n_6320),
.Y(n_7183)
);

INVxp67_ASAP7_75t_L g7184 ( 
.A(n_6677),
.Y(n_7184)
);

AND2x2_ASAP7_75t_L g7185 ( 
.A(n_6658),
.B(n_6320),
.Y(n_7185)
);

INVx2_ASAP7_75t_L g7186 ( 
.A(n_6780),
.Y(n_7186)
);

INVx1_ASAP7_75t_L g7187 ( 
.A(n_6870),
.Y(n_7187)
);

INVx2_ASAP7_75t_L g7188 ( 
.A(n_6807),
.Y(n_7188)
);

OR2x2_ASAP7_75t_L g7189 ( 
.A(n_6782),
.B(n_6428),
.Y(n_7189)
);

INVx1_ASAP7_75t_L g7190 ( 
.A(n_6871),
.Y(n_7190)
);

BUFx2_ASAP7_75t_L g7191 ( 
.A(n_6896),
.Y(n_7191)
);

NAND3xp33_ASAP7_75t_L g7192 ( 
.A(n_6786),
.B(n_6579),
.C(n_6830),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_6872),
.Y(n_7193)
);

BUFx2_ASAP7_75t_L g7194 ( 
.A(n_6896),
.Y(n_7194)
);

NAND2xp5_ASAP7_75t_L g7195 ( 
.A(n_6890),
.B(n_6458),
.Y(n_7195)
);

INVx2_ASAP7_75t_L g7196 ( 
.A(n_6807),
.Y(n_7196)
);

INVx5_ASAP7_75t_L g7197 ( 
.A(n_6844),
.Y(n_7197)
);

AND2x2_ASAP7_75t_L g7198 ( 
.A(n_6661),
.B(n_6349),
.Y(n_7198)
);

NAND4xp25_ASAP7_75t_L g7199 ( 
.A(n_6826),
.B(n_6626),
.C(n_6849),
.D(n_6781),
.Y(n_7199)
);

BUFx2_ASAP7_75t_L g7200 ( 
.A(n_6896),
.Y(n_7200)
);

INVx1_ASAP7_75t_L g7201 ( 
.A(n_6874),
.Y(n_7201)
);

INVx2_ASAP7_75t_L g7202 ( 
.A(n_6816),
.Y(n_7202)
);

OR2x2_ASAP7_75t_L g7203 ( 
.A(n_6797),
.B(n_5301),
.Y(n_7203)
);

AND2x2_ASAP7_75t_L g7204 ( 
.A(n_6661),
.B(n_6349),
.Y(n_7204)
);

HB1xp67_ASAP7_75t_L g7205 ( 
.A(n_6802),
.Y(n_7205)
);

AND2x2_ASAP7_75t_L g7206 ( 
.A(n_6663),
.B(n_6356),
.Y(n_7206)
);

INVx1_ASAP7_75t_L g7207 ( 
.A(n_6875),
.Y(n_7207)
);

HB1xp67_ASAP7_75t_L g7208 ( 
.A(n_6821),
.Y(n_7208)
);

AND2x2_ASAP7_75t_L g7209 ( 
.A(n_6663),
.B(n_6356),
.Y(n_7209)
);

INVx3_ASAP7_75t_L g7210 ( 
.A(n_6648),
.Y(n_7210)
);

INVx1_ASAP7_75t_L g7211 ( 
.A(n_6877),
.Y(n_7211)
);

INVx1_ASAP7_75t_L g7212 ( 
.A(n_6879),
.Y(n_7212)
);

INVx3_ASAP7_75t_L g7213 ( 
.A(n_6648),
.Y(n_7213)
);

OR2x2_ASAP7_75t_L g7214 ( 
.A(n_6703),
.B(n_5301),
.Y(n_7214)
);

INVx1_ASAP7_75t_L g7215 ( 
.A(n_6887),
.Y(n_7215)
);

INVx3_ASAP7_75t_L g7216 ( 
.A(n_6691),
.Y(n_7216)
);

BUFx2_ASAP7_75t_L g7217 ( 
.A(n_6518),
.Y(n_7217)
);

INVxp67_ASAP7_75t_SL g7218 ( 
.A(n_6677),
.Y(n_7218)
);

AND2x2_ASAP7_75t_L g7219 ( 
.A(n_6717),
.B(n_6373),
.Y(n_7219)
);

AND2x4_ASAP7_75t_L g7220 ( 
.A(n_6805),
.B(n_6160),
.Y(n_7220)
);

INVx2_ASAP7_75t_L g7221 ( 
.A(n_6816),
.Y(n_7221)
);

INVxp67_ASAP7_75t_SL g7222 ( 
.A(n_6700),
.Y(n_7222)
);

AND2x2_ASAP7_75t_L g7223 ( 
.A(n_6717),
.B(n_6373),
.Y(n_7223)
);

INVx1_ASAP7_75t_L g7224 ( 
.A(n_6892),
.Y(n_7224)
);

INVx5_ASAP7_75t_L g7225 ( 
.A(n_6873),
.Y(n_7225)
);

INVx2_ASAP7_75t_L g7226 ( 
.A(n_6819),
.Y(n_7226)
);

AND2x2_ASAP7_75t_L g7227 ( 
.A(n_6718),
.B(n_6382),
.Y(n_7227)
);

INVx2_ASAP7_75t_L g7228 ( 
.A(n_6819),
.Y(n_7228)
);

INVx2_ASAP7_75t_L g7229 ( 
.A(n_6964),
.Y(n_7229)
);

NAND2xp5_ASAP7_75t_L g7230 ( 
.A(n_7019),
.B(n_6894),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_6958),
.Y(n_7231)
);

NAND2xp5_ASAP7_75t_L g7232 ( 
.A(n_7019),
.B(n_6997),
.Y(n_7232)
);

NAND2xp5_ASAP7_75t_L g7233 ( 
.A(n_6997),
.B(n_6524),
.Y(n_7233)
);

INVx1_ASAP7_75t_L g7234 ( 
.A(n_6958),
.Y(n_7234)
);

AND2x2_ASAP7_75t_L g7235 ( 
.A(n_7007),
.B(n_6776),
.Y(n_7235)
);

INVxp67_ASAP7_75t_L g7236 ( 
.A(n_6900),
.Y(n_7236)
);

INVx2_ASAP7_75t_L g7237 ( 
.A(n_6964),
.Y(n_7237)
);

AND2x2_ASAP7_75t_L g7238 ( 
.A(n_6955),
.B(n_6593),
.Y(n_7238)
);

OR2x2_ASAP7_75t_L g7239 ( 
.A(n_7217),
.B(n_6655),
.Y(n_7239)
);

AOI22xp33_ASAP7_75t_L g7240 ( 
.A1(n_6908),
.A2(n_6830),
.B1(n_6626),
.B2(n_6865),
.Y(n_7240)
);

NAND2xp5_ASAP7_75t_L g7241 ( 
.A(n_6997),
.B(n_6525),
.Y(n_7241)
);

AND2x2_ASAP7_75t_L g7242 ( 
.A(n_6955),
.B(n_6596),
.Y(n_7242)
);

HB1xp67_ASAP7_75t_L g7243 ( 
.A(n_6969),
.Y(n_7243)
);

BUFx2_ASAP7_75t_SL g7244 ( 
.A(n_6982),
.Y(n_7244)
);

INVx1_ASAP7_75t_L g7245 ( 
.A(n_6969),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_6971),
.Y(n_7246)
);

NAND2x1p5_ASAP7_75t_L g7247 ( 
.A(n_6956),
.B(n_6837),
.Y(n_7247)
);

AND2x4_ASAP7_75t_L g7248 ( 
.A(n_6982),
.B(n_6832),
.Y(n_7248)
);

OR2x2_ASAP7_75t_L g7249 ( 
.A(n_6939),
.B(n_6709),
.Y(n_7249)
);

INVx1_ASAP7_75t_L g7250 ( 
.A(n_6971),
.Y(n_7250)
);

AND2x4_ASAP7_75t_L g7251 ( 
.A(n_6990),
.B(n_6834),
.Y(n_7251)
);

NAND2xp5_ASAP7_75t_L g7252 ( 
.A(n_7028),
.B(n_6536),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_6987),
.Y(n_7253)
);

INVx1_ASAP7_75t_L g7254 ( 
.A(n_6987),
.Y(n_7254)
);

AND2x2_ASAP7_75t_L g7255 ( 
.A(n_7120),
.B(n_6550),
.Y(n_7255)
);

INVxp67_ASAP7_75t_L g7256 ( 
.A(n_7002),
.Y(n_7256)
);

NAND3xp33_ASAP7_75t_L g7257 ( 
.A(n_7008),
.B(n_6786),
.C(n_6682),
.Y(n_7257)
);

INVx1_ASAP7_75t_L g7258 ( 
.A(n_7002),
.Y(n_7258)
);

NAND2xp5_ASAP7_75t_L g7259 ( 
.A(n_7028),
.B(n_6541),
.Y(n_7259)
);

AND2x2_ASAP7_75t_L g7260 ( 
.A(n_6989),
.B(n_6584),
.Y(n_7260)
);

INVx2_ASAP7_75t_L g7261 ( 
.A(n_7009),
.Y(n_7261)
);

INVx1_ASAP7_75t_L g7262 ( 
.A(n_7010),
.Y(n_7262)
);

AND2x2_ASAP7_75t_L g7263 ( 
.A(n_7051),
.B(n_6603),
.Y(n_7263)
);

INVx3_ASAP7_75t_L g7264 ( 
.A(n_7009),
.Y(n_7264)
);

AND2x2_ASAP7_75t_L g7265 ( 
.A(n_7144),
.B(n_6545),
.Y(n_7265)
);

OR2x2_ASAP7_75t_L g7266 ( 
.A(n_6913),
.B(n_6647),
.Y(n_7266)
);

INVx2_ASAP7_75t_L g7267 ( 
.A(n_7009),
.Y(n_7267)
);

INVx1_ASAP7_75t_L g7268 ( 
.A(n_7010),
.Y(n_7268)
);

INVx1_ASAP7_75t_L g7269 ( 
.A(n_7170),
.Y(n_7269)
);

AOI22xp33_ASAP7_75t_SL g7270 ( 
.A1(n_6937),
.A2(n_7192),
.B1(n_6914),
.B2(n_7097),
.Y(n_7270)
);

AND2x2_ASAP7_75t_L g7271 ( 
.A(n_7084),
.B(n_6545),
.Y(n_7271)
);

OR2x2_ASAP7_75t_L g7272 ( 
.A(n_7152),
.B(n_6869),
.Y(n_7272)
);

INVx2_ASAP7_75t_L g7273 ( 
.A(n_7009),
.Y(n_7273)
);

INVx2_ASAP7_75t_L g7274 ( 
.A(n_7034),
.Y(n_7274)
);

AND2x2_ASAP7_75t_L g7275 ( 
.A(n_6972),
.B(n_6718),
.Y(n_7275)
);

AND2x4_ASAP7_75t_L g7276 ( 
.A(n_6990),
.B(n_6859),
.Y(n_7276)
);

INVx1_ASAP7_75t_L g7277 ( 
.A(n_7170),
.Y(n_7277)
);

AND2x2_ASAP7_75t_L g7278 ( 
.A(n_6972),
.B(n_6886),
.Y(n_7278)
);

INVx3_ASAP7_75t_L g7279 ( 
.A(n_7034),
.Y(n_7279)
);

OR2x2_ASAP7_75t_L g7280 ( 
.A(n_6957),
.B(n_6888),
.Y(n_7280)
);

INVx1_ASAP7_75t_L g7281 ( 
.A(n_6916),
.Y(n_7281)
);

INVx1_ASAP7_75t_L g7282 ( 
.A(n_6916),
.Y(n_7282)
);

INVx1_ASAP7_75t_L g7283 ( 
.A(n_6923),
.Y(n_7283)
);

INVxp67_ASAP7_75t_L g7284 ( 
.A(n_7034),
.Y(n_7284)
);

NOR2xp33_ASAP7_75t_SL g7285 ( 
.A(n_7054),
.B(n_6770),
.Y(n_7285)
);

AND2x2_ASAP7_75t_L g7286 ( 
.A(n_6978),
.B(n_6886),
.Y(n_7286)
);

NAND2xp5_ASAP7_75t_L g7287 ( 
.A(n_7056),
.B(n_6542),
.Y(n_7287)
);

NAND2xp5_ASAP7_75t_L g7288 ( 
.A(n_7056),
.B(n_6553),
.Y(n_7288)
);

NAND2xp5_ASAP7_75t_L g7289 ( 
.A(n_7097),
.B(n_6554),
.Y(n_7289)
);

INVx1_ASAP7_75t_L g7290 ( 
.A(n_6923),
.Y(n_7290)
);

AND2x2_ASAP7_75t_L g7291 ( 
.A(n_6978),
.B(n_6895),
.Y(n_7291)
);

INVx1_ASAP7_75t_L g7292 ( 
.A(n_6951),
.Y(n_7292)
);

INVx2_ASAP7_75t_L g7293 ( 
.A(n_7034),
.Y(n_7293)
);

OR2x2_ASAP7_75t_L g7294 ( 
.A(n_7090),
.B(n_6801),
.Y(n_7294)
);

INVx1_ASAP7_75t_L g7295 ( 
.A(n_6951),
.Y(n_7295)
);

OR2x2_ASAP7_75t_L g7296 ( 
.A(n_6906),
.B(n_6815),
.Y(n_7296)
);

OAI221xp5_ASAP7_75t_SL g7297 ( 
.A1(n_7168),
.A2(n_6708),
.B1(n_6531),
.B2(n_6723),
.C(n_6865),
.Y(n_7297)
);

AND2x2_ASAP7_75t_L g7298 ( 
.A(n_6920),
.B(n_7079),
.Y(n_7298)
);

OR2x2_ASAP7_75t_L g7299 ( 
.A(n_7078),
.B(n_6561),
.Y(n_7299)
);

NAND2x1p5_ASAP7_75t_L g7300 ( 
.A(n_6956),
.B(n_6867),
.Y(n_7300)
);

INVx1_ASAP7_75t_L g7301 ( 
.A(n_7035),
.Y(n_7301)
);

INVxp67_ASAP7_75t_L g7302 ( 
.A(n_6993),
.Y(n_7302)
);

INVx1_ASAP7_75t_L g7303 ( 
.A(n_7035),
.Y(n_7303)
);

AND2x2_ASAP7_75t_L g7304 ( 
.A(n_6920),
.B(n_6895),
.Y(n_7304)
);

OR2x2_ASAP7_75t_L g7305 ( 
.A(n_7015),
.B(n_6597),
.Y(n_7305)
);

INVx1_ASAP7_75t_L g7306 ( 
.A(n_6903),
.Y(n_7306)
);

AND2x4_ASAP7_75t_L g7307 ( 
.A(n_7080),
.B(n_6695),
.Y(n_7307)
);

AOI211xp5_ASAP7_75t_L g7308 ( 
.A1(n_6973),
.A2(n_6979),
.B(n_7167),
.C(n_7149),
.Y(n_7308)
);

NAND2xp5_ASAP7_75t_L g7309 ( 
.A(n_7032),
.B(n_6563),
.Y(n_7309)
);

INVxp67_ASAP7_75t_L g7310 ( 
.A(n_7024),
.Y(n_7310)
);

AND2x4_ASAP7_75t_L g7311 ( 
.A(n_7080),
.B(n_6721),
.Y(n_7311)
);

NAND2x1p5_ASAP7_75t_L g7312 ( 
.A(n_6956),
.B(n_6898),
.Y(n_7312)
);

AND2x2_ASAP7_75t_L g7313 ( 
.A(n_6909),
.B(n_6721),
.Y(n_7313)
);

INVxp67_ASAP7_75t_SL g7314 ( 
.A(n_7054),
.Y(n_7314)
);

NOR2xp33_ASAP7_75t_L g7315 ( 
.A(n_6956),
.B(n_7082),
.Y(n_7315)
);

OR2x2_ASAP7_75t_L g7316 ( 
.A(n_7062),
.B(n_6634),
.Y(n_7316)
);

OAI21xp5_ASAP7_75t_L g7317 ( 
.A1(n_7168),
.A2(n_6682),
.B(n_6729),
.Y(n_7317)
);

AND2x2_ASAP7_75t_L g7318 ( 
.A(n_6909),
.B(n_6925),
.Y(n_7318)
);

HB1xp67_ASAP7_75t_L g7319 ( 
.A(n_6988),
.Y(n_7319)
);

INVx1_ASAP7_75t_L g7320 ( 
.A(n_6911),
.Y(n_7320)
);

OR2x2_ASAP7_75t_L g7321 ( 
.A(n_7203),
.B(n_6602),
.Y(n_7321)
);

HB1xp67_ASAP7_75t_L g7322 ( 
.A(n_6988),
.Y(n_7322)
);

NAND2xp5_ASAP7_75t_L g7323 ( 
.A(n_7032),
.B(n_6566),
.Y(n_7323)
);

BUFx3_ASAP7_75t_L g7324 ( 
.A(n_7082),
.Y(n_7324)
);

AND2x2_ASAP7_75t_L g7325 ( 
.A(n_6925),
.B(n_6787),
.Y(n_7325)
);

HB1xp67_ASAP7_75t_L g7326 ( 
.A(n_6912),
.Y(n_7326)
);

AND2x2_ASAP7_75t_L g7327 ( 
.A(n_6929),
.B(n_6787),
.Y(n_7327)
);

INVx1_ASAP7_75t_L g7328 ( 
.A(n_6915),
.Y(n_7328)
);

INVx1_ASAP7_75t_L g7329 ( 
.A(n_6917),
.Y(n_7329)
);

INVx2_ASAP7_75t_L g7330 ( 
.A(n_7082),
.Y(n_7330)
);

INVx2_ASAP7_75t_L g7331 ( 
.A(n_7082),
.Y(n_7331)
);

HB1xp67_ASAP7_75t_L g7332 ( 
.A(n_6931),
.Y(n_7332)
);

NAND2xp5_ASAP7_75t_L g7333 ( 
.A(n_7085),
.B(n_6567),
.Y(n_7333)
);

INVx1_ASAP7_75t_L g7334 ( 
.A(n_6933),
.Y(n_7334)
);

AND2x4_ASAP7_75t_L g7335 ( 
.A(n_7141),
.B(n_6882),
.Y(n_7335)
);

AND2x2_ASAP7_75t_L g7336 ( 
.A(n_6929),
.B(n_6790),
.Y(n_7336)
);

OR2x2_ASAP7_75t_L g7337 ( 
.A(n_7214),
.B(n_6610),
.Y(n_7337)
);

INVxp67_ASAP7_75t_L g7338 ( 
.A(n_6945),
.Y(n_7338)
);

NOR2x1_ASAP7_75t_L g7339 ( 
.A(n_7139),
.B(n_6826),
.Y(n_7339)
);

AND2x2_ASAP7_75t_L g7340 ( 
.A(n_7136),
.B(n_6790),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_6949),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_L g7342 ( 
.A(n_7085),
.B(n_6575),
.Y(n_7342)
);

AND2x2_ASAP7_75t_L g7343 ( 
.A(n_7162),
.B(n_6652),
.Y(n_7343)
);

INVx1_ASAP7_75t_L g7344 ( 
.A(n_6965),
.Y(n_7344)
);

INVx1_ASAP7_75t_L g7345 ( 
.A(n_6970),
.Y(n_7345)
);

HB1xp67_ASAP7_75t_L g7346 ( 
.A(n_6975),
.Y(n_7346)
);

AND2x2_ASAP7_75t_L g7347 ( 
.A(n_7164),
.B(n_6652),
.Y(n_7347)
);

INVx2_ASAP7_75t_L g7348 ( 
.A(n_7191),
.Y(n_7348)
);

NAND3xp33_ASAP7_75t_L g7349 ( 
.A(n_7033),
.B(n_6581),
.C(n_6577),
.Y(n_7349)
);

AND2x2_ASAP7_75t_L g7350 ( 
.A(n_7194),
.B(n_7200),
.Y(n_7350)
);

HB1xp67_ASAP7_75t_L g7351 ( 
.A(n_6977),
.Y(n_7351)
);

INVx2_ASAP7_75t_SL g7352 ( 
.A(n_6992),
.Y(n_7352)
);

NAND2xp5_ASAP7_75t_L g7353 ( 
.A(n_7205),
.B(n_6576),
.Y(n_7353)
);

AND2x4_ASAP7_75t_L g7354 ( 
.A(n_7141),
.B(n_6805),
.Y(n_7354)
);

NAND2xp5_ASAP7_75t_L g7355 ( 
.A(n_7205),
.B(n_6578),
.Y(n_7355)
);

NAND3xp33_ASAP7_75t_L g7356 ( 
.A(n_7060),
.B(n_7046),
.C(n_7099),
.Y(n_7356)
);

AND2x2_ASAP7_75t_L g7357 ( 
.A(n_7061),
.B(n_6922),
.Y(n_7357)
);

NAND2xp5_ASAP7_75t_L g7358 ( 
.A(n_7208),
.B(n_6582),
.Y(n_7358)
);

HB1xp67_ASAP7_75t_L g7359 ( 
.A(n_6981),
.Y(n_7359)
);

INVx1_ASAP7_75t_L g7360 ( 
.A(n_6985),
.Y(n_7360)
);

INVx2_ASAP7_75t_L g7361 ( 
.A(n_7210),
.Y(n_7361)
);

BUFx3_ASAP7_75t_L g7362 ( 
.A(n_6928),
.Y(n_7362)
);

BUFx2_ASAP7_75t_L g7363 ( 
.A(n_7083),
.Y(n_7363)
);

AND2x4_ASAP7_75t_L g7364 ( 
.A(n_7141),
.B(n_6805),
.Y(n_7364)
);

INVx1_ASAP7_75t_L g7365 ( 
.A(n_6907),
.Y(n_7365)
);

AND2x2_ASAP7_75t_L g7366 ( 
.A(n_6922),
.B(n_6653),
.Y(n_7366)
);

AND2x2_ASAP7_75t_L g7367 ( 
.A(n_6967),
.B(n_6653),
.Y(n_7367)
);

AND2x4_ASAP7_75t_SL g7368 ( 
.A(n_7063),
.B(n_6884),
.Y(n_7368)
);

AND2x2_ASAP7_75t_L g7369 ( 
.A(n_6967),
.B(n_6843),
.Y(n_7369)
);

AND2x2_ASAP7_75t_L g7370 ( 
.A(n_7128),
.B(n_6843),
.Y(n_7370)
);

OR2x2_ASAP7_75t_L g7371 ( 
.A(n_7049),
.B(n_6828),
.Y(n_7371)
);

INVx1_ASAP7_75t_L g7372 ( 
.A(n_6907),
.Y(n_7372)
);

AND2x4_ASAP7_75t_L g7373 ( 
.A(n_7063),
.B(n_6836),
.Y(n_7373)
);

AND2x2_ASAP7_75t_L g7374 ( 
.A(n_7083),
.B(n_6856),
.Y(n_7374)
);

AND2x2_ASAP7_75t_L g7375 ( 
.A(n_7083),
.B(n_6856),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_6921),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_6921),
.Y(n_7377)
);

AND2x2_ASAP7_75t_L g7378 ( 
.A(n_7016),
.B(n_6858),
.Y(n_7378)
);

NAND2xp5_ASAP7_75t_L g7379 ( 
.A(n_7208),
.B(n_6586),
.Y(n_7379)
);

INVxp67_ASAP7_75t_L g7380 ( 
.A(n_7068),
.Y(n_7380)
);

AND2x2_ASAP7_75t_L g7381 ( 
.A(n_7016),
.B(n_6858),
.Y(n_7381)
);

NAND2xp5_ASAP7_75t_L g7382 ( 
.A(n_7098),
.B(n_6587),
.Y(n_7382)
);

INVx1_ASAP7_75t_L g7383 ( 
.A(n_6926),
.Y(n_7383)
);

INVx1_ASAP7_75t_L g7384 ( 
.A(n_6926),
.Y(n_7384)
);

AND2x2_ASAP7_75t_L g7385 ( 
.A(n_7161),
.B(n_7165),
.Y(n_7385)
);

INVx1_ASAP7_75t_L g7386 ( 
.A(n_6950),
.Y(n_7386)
);

AND2x2_ASAP7_75t_L g7387 ( 
.A(n_7183),
.B(n_6645),
.Y(n_7387)
);

AND2x2_ASAP7_75t_L g7388 ( 
.A(n_7183),
.B(n_6645),
.Y(n_7388)
);

NAND2xp5_ASAP7_75t_L g7389 ( 
.A(n_7098),
.B(n_6588),
.Y(n_7389)
);

NAND2x1p5_ASAP7_75t_L g7390 ( 
.A(n_6968),
.B(n_6898),
.Y(n_7390)
);

INVx3_ASAP7_75t_L g7391 ( 
.A(n_6966),
.Y(n_7391)
);

INVx3_ASAP7_75t_L g7392 ( 
.A(n_6966),
.Y(n_7392)
);

AND2x4_ASAP7_75t_SL g7393 ( 
.A(n_6941),
.B(n_6935),
.Y(n_7393)
);

AND2x2_ASAP7_75t_L g7394 ( 
.A(n_7185),
.B(n_7198),
.Y(n_7394)
);

INVx2_ASAP7_75t_L g7395 ( 
.A(n_7210),
.Y(n_7395)
);

INVx2_ASAP7_75t_L g7396 ( 
.A(n_7210),
.Y(n_7396)
);

AND2x2_ASAP7_75t_L g7397 ( 
.A(n_7185),
.B(n_6650),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_6950),
.Y(n_7398)
);

AND2x2_ASAP7_75t_L g7399 ( 
.A(n_7198),
.B(n_6650),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_6950),
.Y(n_7400)
);

INVx1_ASAP7_75t_L g7401 ( 
.A(n_6927),
.Y(n_7401)
);

AND2x2_ASAP7_75t_L g7402 ( 
.A(n_7204),
.B(n_7206),
.Y(n_7402)
);

AND2x4_ASAP7_75t_L g7403 ( 
.A(n_7063),
.B(n_7058),
.Y(n_7403)
);

OR2x2_ASAP7_75t_L g7404 ( 
.A(n_7055),
.B(n_6570),
.Y(n_7404)
);

AND2x2_ASAP7_75t_L g7405 ( 
.A(n_7204),
.B(n_6884),
.Y(n_7405)
);

INVx1_ASAP7_75t_L g7406 ( 
.A(n_6927),
.Y(n_7406)
);

NAND2xp5_ASAP7_75t_L g7407 ( 
.A(n_7113),
.B(n_6595),
.Y(n_7407)
);

INVx1_ASAP7_75t_L g7408 ( 
.A(n_6940),
.Y(n_7408)
);

AND2x2_ASAP7_75t_L g7409 ( 
.A(n_7206),
.B(n_6794),
.Y(n_7409)
);

AND2x4_ASAP7_75t_L g7410 ( 
.A(n_7058),
.B(n_6836),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_6940),
.Y(n_7411)
);

INVx1_ASAP7_75t_L g7412 ( 
.A(n_6943),
.Y(n_7412)
);

AND2x4_ASAP7_75t_L g7413 ( 
.A(n_7058),
.B(n_6836),
.Y(n_7413)
);

INVx1_ASAP7_75t_L g7414 ( 
.A(n_6943),
.Y(n_7414)
);

AND2x2_ASAP7_75t_L g7415 ( 
.A(n_7209),
.B(n_6794),
.Y(n_7415)
);

NAND2x1p5_ASAP7_75t_L g7416 ( 
.A(n_6968),
.B(n_7139),
.Y(n_7416)
);

AND2x2_ASAP7_75t_L g7417 ( 
.A(n_7209),
.B(n_6631),
.Y(n_7417)
);

AND2x2_ASAP7_75t_L g7418 ( 
.A(n_7219),
.B(n_6631),
.Y(n_7418)
);

NAND2xp5_ASAP7_75t_L g7419 ( 
.A(n_7113),
.B(n_6598),
.Y(n_7419)
);

NAND2x1_ASAP7_75t_L g7420 ( 
.A(n_6953),
.B(n_6691),
.Y(n_7420)
);

INVx1_ASAP7_75t_L g7421 ( 
.A(n_6946),
.Y(n_7421)
);

NAND2x1_ASAP7_75t_SL g7422 ( 
.A(n_6966),
.B(n_6691),
.Y(n_7422)
);

INVx1_ASAP7_75t_L g7423 ( 
.A(n_6946),
.Y(n_7423)
);

NAND2xp5_ASAP7_75t_L g7424 ( 
.A(n_7126),
.B(n_6599),
.Y(n_7424)
);

AND2x2_ASAP7_75t_L g7425 ( 
.A(n_7219),
.B(n_6770),
.Y(n_7425)
);

AND2x2_ASAP7_75t_L g7426 ( 
.A(n_7223),
.B(n_6770),
.Y(n_7426)
);

AND2x2_ASAP7_75t_L g7427 ( 
.A(n_7223),
.B(n_6770),
.Y(n_7427)
);

INVx3_ASAP7_75t_L g7428 ( 
.A(n_6919),
.Y(n_7428)
);

INVx1_ASAP7_75t_L g7429 ( 
.A(n_6947),
.Y(n_7429)
);

BUFx6f_ASAP7_75t_L g7430 ( 
.A(n_7131),
.Y(n_7430)
);

AND2x2_ASAP7_75t_L g7431 ( 
.A(n_7227),
.B(n_6742),
.Y(n_7431)
);

INVx1_ASAP7_75t_L g7432 ( 
.A(n_6947),
.Y(n_7432)
);

NOR2xp67_ASAP7_75t_L g7433 ( 
.A(n_7213),
.B(n_6710),
.Y(n_7433)
);

NOR2xp33_ASAP7_75t_L g7434 ( 
.A(n_7139),
.B(n_6704),
.Y(n_7434)
);

INVx2_ASAP7_75t_L g7435 ( 
.A(n_7213),
.Y(n_7435)
);

AND2x2_ASAP7_75t_L g7436 ( 
.A(n_7227),
.B(n_6742),
.Y(n_7436)
);

INVx1_ASAP7_75t_L g7437 ( 
.A(n_6948),
.Y(n_7437)
);

AND2x2_ASAP7_75t_L g7438 ( 
.A(n_6986),
.B(n_6984),
.Y(n_7438)
);

NAND2xp5_ASAP7_75t_L g7439 ( 
.A(n_7126),
.B(n_6604),
.Y(n_7439)
);

NAND2xp5_ASAP7_75t_L g7440 ( 
.A(n_7006),
.B(n_6606),
.Y(n_7440)
);

AND2x4_ASAP7_75t_L g7441 ( 
.A(n_7213),
.B(n_6696),
.Y(n_7441)
);

NOR3xp33_ASAP7_75t_L g7442 ( 
.A(n_7171),
.B(n_6581),
.C(n_6577),
.Y(n_7442)
);

OR2x2_ASAP7_75t_L g7443 ( 
.A(n_7070),
.B(n_6839),
.Y(n_7443)
);

BUFx2_ASAP7_75t_L g7444 ( 
.A(n_7027),
.Y(n_7444)
);

AND2x2_ASAP7_75t_L g7445 ( 
.A(n_7154),
.B(n_6744),
.Y(n_7445)
);

NAND2xp5_ASAP7_75t_L g7446 ( 
.A(n_7006),
.B(n_6607),
.Y(n_7446)
);

AND2x2_ASAP7_75t_L g7447 ( 
.A(n_7156),
.B(n_6744),
.Y(n_7447)
);

AND2x4_ASAP7_75t_L g7448 ( 
.A(n_7216),
.B(n_7132),
.Y(n_7448)
);

INVx2_ASAP7_75t_L g7449 ( 
.A(n_7216),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_6948),
.Y(n_7450)
);

INVx2_ASAP7_75t_L g7451 ( 
.A(n_7216),
.Y(n_7451)
);

INVxp67_ASAP7_75t_SL g7452 ( 
.A(n_7149),
.Y(n_7452)
);

OR2x2_ASAP7_75t_L g7453 ( 
.A(n_7036),
.B(n_6862),
.Y(n_7453)
);

BUFx2_ASAP7_75t_L g7454 ( 
.A(n_7027),
.Y(n_7454)
);

AND2x2_ASAP7_75t_L g7455 ( 
.A(n_6994),
.B(n_6534),
.Y(n_7455)
);

NAND2xp5_ASAP7_75t_L g7456 ( 
.A(n_7012),
.B(n_6613),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_6944),
.Y(n_7457)
);

OR2x2_ASAP7_75t_L g7458 ( 
.A(n_6996),
.B(n_6848),
.Y(n_7458)
);

INVx1_ASAP7_75t_L g7459 ( 
.A(n_6944),
.Y(n_7459)
);

INVx2_ASAP7_75t_L g7460 ( 
.A(n_6992),
.Y(n_7460)
);

NOR2xp33_ASAP7_75t_L g7461 ( 
.A(n_7050),
.B(n_6687),
.Y(n_7461)
);

INVx2_ASAP7_75t_L g7462 ( 
.A(n_7052),
.Y(n_7462)
);

AND2x2_ASAP7_75t_L g7463 ( 
.A(n_7102),
.B(n_6696),
.Y(n_7463)
);

OR2x2_ASAP7_75t_L g7464 ( 
.A(n_7073),
.B(n_6702),
.Y(n_7464)
);

AND2x2_ASAP7_75t_L g7465 ( 
.A(n_7102),
.B(n_6696),
.Y(n_7465)
);

INVx2_ASAP7_75t_L g7466 ( 
.A(n_7052),
.Y(n_7466)
);

AND2x2_ASAP7_75t_L g7467 ( 
.A(n_7104),
.B(n_6756),
.Y(n_7467)
);

BUFx2_ASAP7_75t_L g7468 ( 
.A(n_7027),
.Y(n_7468)
);

NAND2xp5_ASAP7_75t_L g7469 ( 
.A(n_7012),
.B(n_6615),
.Y(n_7469)
);

AND2x2_ASAP7_75t_L g7470 ( 
.A(n_7104),
.B(n_6710),
.Y(n_7470)
);

INVx1_ASAP7_75t_L g7471 ( 
.A(n_6998),
.Y(n_7471)
);

AND2x2_ASAP7_75t_L g7472 ( 
.A(n_7111),
.B(n_6688),
.Y(n_7472)
);

INVx2_ASAP7_75t_L g7473 ( 
.A(n_7052),
.Y(n_7473)
);

OR2x2_ASAP7_75t_L g7474 ( 
.A(n_7075),
.B(n_6705),
.Y(n_7474)
);

AND2x2_ASAP7_75t_L g7475 ( 
.A(n_7111),
.B(n_6694),
.Y(n_7475)
);

AND2x2_ASAP7_75t_L g7476 ( 
.A(n_7064),
.B(n_6654),
.Y(n_7476)
);

NOR2x1_ASAP7_75t_L g7477 ( 
.A(n_7199),
.B(n_6758),
.Y(n_7477)
);

NOR2x1p5_ASAP7_75t_L g7478 ( 
.A(n_7087),
.B(n_6685),
.Y(n_7478)
);

INVxp67_ASAP7_75t_SL g7479 ( 
.A(n_7157),
.Y(n_7479)
);

INVxp67_ASAP7_75t_L g7480 ( 
.A(n_6928),
.Y(n_7480)
);

NOR2xp33_ASAP7_75t_L g7481 ( 
.A(n_7053),
.B(n_6785),
.Y(n_7481)
);

AND2x4_ASAP7_75t_SL g7482 ( 
.A(n_6924),
.B(n_6960),
.Y(n_7482)
);

INVx2_ASAP7_75t_L g7483 ( 
.A(n_7081),
.Y(n_7483)
);

OR2x2_ASAP7_75t_L g7484 ( 
.A(n_6959),
.B(n_6707),
.Y(n_7484)
);

INVx2_ASAP7_75t_L g7485 ( 
.A(n_7081),
.Y(n_7485)
);

NAND2xp5_ASAP7_75t_L g7486 ( 
.A(n_7014),
.B(n_6622),
.Y(n_7486)
);

INVx1_ASAP7_75t_L g7487 ( 
.A(n_6998),
.Y(n_7487)
);

AND2x2_ASAP7_75t_L g7488 ( 
.A(n_7064),
.B(n_6025),
.Y(n_7488)
);

AND2x2_ASAP7_75t_L g7489 ( 
.A(n_6902),
.B(n_6771),
.Y(n_7489)
);

INVx2_ASAP7_75t_L g7490 ( 
.A(n_7081),
.Y(n_7490)
);

INVx1_ASAP7_75t_L g7491 ( 
.A(n_6934),
.Y(n_7491)
);

NAND2xp5_ASAP7_75t_L g7492 ( 
.A(n_7014),
.B(n_6627),
.Y(n_7492)
);

NAND2xp5_ASAP7_75t_L g7493 ( 
.A(n_6942),
.B(n_6630),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_6934),
.Y(n_7494)
);

AND2x2_ASAP7_75t_L g7495 ( 
.A(n_6902),
.B(n_6715),
.Y(n_7495)
);

INVx1_ASAP7_75t_L g7496 ( 
.A(n_6962),
.Y(n_7496)
);

NAND2xp5_ASAP7_75t_L g7497 ( 
.A(n_6942),
.B(n_6635),
.Y(n_7497)
);

OR2x2_ASAP7_75t_L g7498 ( 
.A(n_6963),
.B(n_7103),
.Y(n_7498)
);

INVx1_ASAP7_75t_L g7499 ( 
.A(n_7166),
.Y(n_7499)
);

AND2x2_ASAP7_75t_L g7500 ( 
.A(n_7067),
.B(n_6726),
.Y(n_7500)
);

NOR2xp33_ASAP7_75t_L g7501 ( 
.A(n_7132),
.B(n_6728),
.Y(n_7501)
);

INVx1_ASAP7_75t_L g7502 ( 
.A(n_7166),
.Y(n_7502)
);

AND2x2_ASAP7_75t_L g7503 ( 
.A(n_7076),
.B(n_6732),
.Y(n_7503)
);

INVx2_ASAP7_75t_L g7504 ( 
.A(n_7091),
.Y(n_7504)
);

AND2x2_ASAP7_75t_L g7505 ( 
.A(n_7037),
.B(n_6735),
.Y(n_7505)
);

INVx1_ASAP7_75t_L g7506 ( 
.A(n_6991),
.Y(n_7506)
);

AND2x2_ASAP7_75t_L g7507 ( 
.A(n_7037),
.B(n_6110),
.Y(n_7507)
);

INVx1_ASAP7_75t_L g7508 ( 
.A(n_6999),
.Y(n_7508)
);

AND2x2_ASAP7_75t_L g7509 ( 
.A(n_7038),
.B(n_6112),
.Y(n_7509)
);

AND2x4_ASAP7_75t_L g7510 ( 
.A(n_6924),
.B(n_6960),
.Y(n_7510)
);

AND2x4_ASAP7_75t_L g7511 ( 
.A(n_6924),
.B(n_6960),
.Y(n_7511)
);

OR2x2_ASAP7_75t_L g7512 ( 
.A(n_7189),
.B(n_6636),
.Y(n_7512)
);

AND2x2_ASAP7_75t_L g7513 ( 
.A(n_7318),
.B(n_6905),
.Y(n_7513)
);

NOR2x1_ASAP7_75t_L g7514 ( 
.A(n_7324),
.B(n_7140),
.Y(n_7514)
);

OR2x2_ASAP7_75t_L g7515 ( 
.A(n_7272),
.B(n_7222),
.Y(n_7515)
);

NOR3xp33_ASAP7_75t_L g7516 ( 
.A(n_7232),
.B(n_7176),
.C(n_7099),
.Y(n_7516)
);

INVx1_ASAP7_75t_L g7517 ( 
.A(n_7243),
.Y(n_7517)
);

NOR3xp33_ASAP7_75t_SL g7518 ( 
.A(n_7479),
.B(n_7022),
.C(n_7218),
.Y(n_7518)
);

AND2x2_ASAP7_75t_L g7519 ( 
.A(n_7378),
.B(n_6905),
.Y(n_7519)
);

INVx1_ASAP7_75t_L g7520 ( 
.A(n_7243),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_7314),
.Y(n_7521)
);

BUFx3_ASAP7_75t_L g7522 ( 
.A(n_7362),
.Y(n_7522)
);

NAND2xp5_ASAP7_75t_L g7523 ( 
.A(n_7381),
.B(n_7110),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_7314),
.Y(n_7524)
);

AND2x2_ASAP7_75t_L g7525 ( 
.A(n_7369),
.B(n_7040),
.Y(n_7525)
);

NAND2xp5_ASAP7_75t_L g7526 ( 
.A(n_7367),
.B(n_7123),
.Y(n_7526)
);

AND2x2_ASAP7_75t_L g7527 ( 
.A(n_7304),
.B(n_7040),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_7319),
.Y(n_7528)
);

NAND2xp5_ASAP7_75t_L g7529 ( 
.A(n_7275),
.B(n_6938),
.Y(n_7529)
);

OR2x2_ASAP7_75t_L g7530 ( 
.A(n_7299),
.B(n_7101),
.Y(n_7530)
);

AND2x2_ASAP7_75t_L g7531 ( 
.A(n_7238),
.B(n_7242),
.Y(n_7531)
);

OR2x2_ASAP7_75t_L g7532 ( 
.A(n_7239),
.B(n_6976),
.Y(n_7532)
);

NAND2xp5_ASAP7_75t_L g7533 ( 
.A(n_7387),
.B(n_7095),
.Y(n_7533)
);

AND2x2_ASAP7_75t_L g7534 ( 
.A(n_7278),
.B(n_7040),
.Y(n_7534)
);

AND2x2_ASAP7_75t_L g7535 ( 
.A(n_7286),
.B(n_7092),
.Y(n_7535)
);

AND2x2_ASAP7_75t_L g7536 ( 
.A(n_7291),
.B(n_7325),
.Y(n_7536)
);

NOR2xp33_ASAP7_75t_L g7537 ( 
.A(n_7356),
.B(n_7131),
.Y(n_7537)
);

INVxp67_ASAP7_75t_L g7538 ( 
.A(n_7244),
.Y(n_7538)
);

INVx1_ASAP7_75t_L g7539 ( 
.A(n_7319),
.Y(n_7539)
);

AND2x4_ASAP7_75t_L g7540 ( 
.A(n_7403),
.B(n_7131),
.Y(n_7540)
);

NOR2xp33_ASAP7_75t_L g7541 ( 
.A(n_7356),
.B(n_7121),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7322),
.Y(n_7542)
);

OAI221xp5_ASAP7_75t_L g7543 ( 
.A1(n_7270),
.A2(n_7060),
.B1(n_7046),
.B2(n_6974),
.C(n_6845),
.Y(n_7543)
);

BUFx2_ASAP7_75t_L g7544 ( 
.A(n_7422),
.Y(n_7544)
);

INVx1_ASAP7_75t_L g7545 ( 
.A(n_7322),
.Y(n_7545)
);

AND2x2_ASAP7_75t_L g7546 ( 
.A(n_7327),
.B(n_7092),
.Y(n_7546)
);

AND2x2_ASAP7_75t_L g7547 ( 
.A(n_7336),
.B(n_7130),
.Y(n_7547)
);

INVx1_ASAP7_75t_L g7548 ( 
.A(n_7350),
.Y(n_7548)
);

OR2x6_ASAP7_75t_L g7549 ( 
.A(n_7284),
.B(n_6968),
.Y(n_7549)
);

OR2x2_ASAP7_75t_L g7550 ( 
.A(n_7249),
.B(n_6983),
.Y(n_7550)
);

INVx2_ASAP7_75t_SL g7551 ( 
.A(n_7482),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_7280),
.Y(n_7552)
);

AND2x2_ASAP7_75t_L g7553 ( 
.A(n_7394),
.B(n_7135),
.Y(n_7553)
);

AND2x2_ASAP7_75t_L g7554 ( 
.A(n_7402),
.B(n_7038),
.Y(n_7554)
);

NAND2xp5_ASAP7_75t_SL g7555 ( 
.A(n_7270),
.B(n_7232),
.Y(n_7555)
);

AND2x4_ASAP7_75t_L g7556 ( 
.A(n_7403),
.B(n_7112),
.Y(n_7556)
);

NAND2xp33_ASAP7_75t_SL g7557 ( 
.A(n_7420),
.B(n_7022),
.Y(n_7557)
);

AND2x2_ASAP7_75t_L g7558 ( 
.A(n_7438),
.B(n_7039),
.Y(n_7558)
);

INVx2_ASAP7_75t_L g7559 ( 
.A(n_7457),
.Y(n_7559)
);

INVx2_ASAP7_75t_L g7560 ( 
.A(n_7459),
.Y(n_7560)
);

AND2x2_ASAP7_75t_L g7561 ( 
.A(n_7340),
.B(n_7039),
.Y(n_7561)
);

OAI31xp33_ASAP7_75t_L g7562 ( 
.A1(n_7297),
.A2(n_6845),
.A3(n_7048),
.B(n_6580),
.Y(n_7562)
);

NAND2xp5_ASAP7_75t_L g7563 ( 
.A(n_7388),
.B(n_7397),
.Y(n_7563)
);

AND2x2_ASAP7_75t_L g7564 ( 
.A(n_7370),
.B(n_7094),
.Y(n_7564)
);

INVx1_ASAP7_75t_L g7565 ( 
.A(n_7363),
.Y(n_7565)
);

AND2x2_ASAP7_75t_L g7566 ( 
.A(n_7374),
.B(n_7094),
.Y(n_7566)
);

NAND2xp5_ASAP7_75t_L g7567 ( 
.A(n_7399),
.B(n_6954),
.Y(n_7567)
);

INVx1_ASAP7_75t_L g7568 ( 
.A(n_7326),
.Y(n_7568)
);

AND2x2_ASAP7_75t_L g7569 ( 
.A(n_7375),
.B(n_7343),
.Y(n_7569)
);

NAND2xp5_ASAP7_75t_L g7570 ( 
.A(n_7479),
.B(n_7347),
.Y(n_7570)
);

OR2x2_ASAP7_75t_L g7571 ( 
.A(n_7266),
.B(n_7071),
.Y(n_7571)
);

INVx2_ASAP7_75t_L g7572 ( 
.A(n_7471),
.Y(n_7572)
);

AND2x2_ASAP7_75t_L g7573 ( 
.A(n_7298),
.B(n_7409),
.Y(n_7573)
);

AND2x4_ASAP7_75t_L g7574 ( 
.A(n_7428),
.B(n_7112),
.Y(n_7574)
);

NOR2x1_ASAP7_75t_L g7575 ( 
.A(n_7324),
.B(n_7140),
.Y(n_7575)
);

AND2x2_ASAP7_75t_L g7576 ( 
.A(n_7415),
.B(n_7047),
.Y(n_7576)
);

INVx1_ASAP7_75t_L g7577 ( 
.A(n_7326),
.Y(n_7577)
);

BUFx2_ASAP7_75t_L g7578 ( 
.A(n_7354),
.Y(n_7578)
);

NAND2xp5_ASAP7_75t_L g7579 ( 
.A(n_7366),
.B(n_6954),
.Y(n_7579)
);

AND2x2_ASAP7_75t_L g7580 ( 
.A(n_7357),
.B(n_7018),
.Y(n_7580)
);

HB1xp67_ASAP7_75t_L g7581 ( 
.A(n_7487),
.Y(n_7581)
);

HB1xp67_ASAP7_75t_L g7582 ( 
.A(n_7491),
.Y(n_7582)
);

AND2x2_ASAP7_75t_L g7583 ( 
.A(n_7263),
.B(n_7018),
.Y(n_7583)
);

AND2x4_ASAP7_75t_L g7584 ( 
.A(n_7428),
.B(n_7112),
.Y(n_7584)
);

NAND2xp5_ASAP7_75t_L g7585 ( 
.A(n_7448),
.B(n_6961),
.Y(n_7585)
);

OR2x2_ASAP7_75t_L g7586 ( 
.A(n_7236),
.B(n_7159),
.Y(n_7586)
);

OR2x2_ASAP7_75t_L g7587 ( 
.A(n_7236),
.B(n_7074),
.Y(n_7587)
);

INVx2_ASAP7_75t_L g7588 ( 
.A(n_7494),
.Y(n_7588)
);

AND2x2_ASAP7_75t_L g7589 ( 
.A(n_7482),
.B(n_7137),
.Y(n_7589)
);

INVxp67_ASAP7_75t_L g7590 ( 
.A(n_7285),
.Y(n_7590)
);

OR2x2_ASAP7_75t_L g7591 ( 
.A(n_7294),
.B(n_7321),
.Y(n_7591)
);

INVxp67_ASAP7_75t_L g7592 ( 
.A(n_7285),
.Y(n_7592)
);

AND2x2_ASAP7_75t_L g7593 ( 
.A(n_7418),
.B(n_7153),
.Y(n_7593)
);

INVx3_ASAP7_75t_L g7594 ( 
.A(n_7354),
.Y(n_7594)
);

NAND2xp5_ASAP7_75t_L g7595 ( 
.A(n_7448),
.B(n_6961),
.Y(n_7595)
);

INVx1_ASAP7_75t_SL g7596 ( 
.A(n_7489),
.Y(n_7596)
);

OAI211xp5_ASAP7_75t_SL g7597 ( 
.A1(n_7308),
.A2(n_6910),
.B(n_7184),
.C(n_7077),
.Y(n_7597)
);

NOR2xp33_ASAP7_75t_L g7598 ( 
.A(n_7391),
.B(n_7140),
.Y(n_7598)
);

NOR2xp67_ASAP7_75t_L g7599 ( 
.A(n_7391),
.B(n_6904),
.Y(n_7599)
);

INVx1_ASAP7_75t_L g7600 ( 
.A(n_7332),
.Y(n_7600)
);

INVx1_ASAP7_75t_SL g7601 ( 
.A(n_7235),
.Y(n_7601)
);

AND2x2_ASAP7_75t_L g7602 ( 
.A(n_7385),
.B(n_6930),
.Y(n_7602)
);

AND2x2_ASAP7_75t_L g7603 ( 
.A(n_7417),
.B(n_6932),
.Y(n_7603)
);

AND2x2_ASAP7_75t_L g7604 ( 
.A(n_7463),
.B(n_6901),
.Y(n_7604)
);

INVx1_ASAP7_75t_L g7605 ( 
.A(n_7332),
.Y(n_7605)
);

AND2x2_ASAP7_75t_L g7606 ( 
.A(n_7465),
.B(n_6901),
.Y(n_7606)
);

INVx2_ASAP7_75t_L g7607 ( 
.A(n_7392),
.Y(n_7607)
);

AND2x2_ASAP7_75t_L g7608 ( 
.A(n_7431),
.B(n_7077),
.Y(n_7608)
);

AND2x2_ASAP7_75t_L g7609 ( 
.A(n_7436),
.B(n_7157),
.Y(n_7609)
);

OR2x2_ASAP7_75t_L g7610 ( 
.A(n_7337),
.B(n_7129),
.Y(n_7610)
);

HB1xp67_ASAP7_75t_L g7611 ( 
.A(n_7309),
.Y(n_7611)
);

INVx2_ASAP7_75t_L g7612 ( 
.A(n_7392),
.Y(n_7612)
);

AND2x2_ASAP7_75t_L g7613 ( 
.A(n_7265),
.B(n_7044),
.Y(n_7613)
);

INVx2_ASAP7_75t_L g7614 ( 
.A(n_7510),
.Y(n_7614)
);

NAND2xp5_ASAP7_75t_L g7615 ( 
.A(n_7362),
.B(n_7091),
.Y(n_7615)
);

INVx3_ASAP7_75t_L g7616 ( 
.A(n_7364),
.Y(n_7616)
);

AND2x2_ASAP7_75t_L g7617 ( 
.A(n_7271),
.B(n_7134),
.Y(n_7617)
);

NAND2xp5_ASAP7_75t_L g7618 ( 
.A(n_7495),
.B(n_7338),
.Y(n_7618)
);

INVx1_ASAP7_75t_L g7619 ( 
.A(n_7346),
.Y(n_7619)
);

NAND2xp5_ASAP7_75t_L g7620 ( 
.A(n_7338),
.B(n_7091),
.Y(n_7620)
);

INVx1_ASAP7_75t_L g7621 ( 
.A(n_7346),
.Y(n_7621)
);

NAND2xp5_ASAP7_75t_SL g7622 ( 
.A(n_7309),
.B(n_7197),
.Y(n_7622)
);

BUFx3_ASAP7_75t_L g7623 ( 
.A(n_7248),
.Y(n_7623)
);

AND2x2_ASAP7_75t_L g7624 ( 
.A(n_7313),
.B(n_7182),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_7351),
.Y(n_7625)
);

INVx3_ASAP7_75t_L g7626 ( 
.A(n_7364),
.Y(n_7626)
);

INVx1_ASAP7_75t_L g7627 ( 
.A(n_7351),
.Y(n_7627)
);

INVx1_ASAP7_75t_L g7628 ( 
.A(n_7359),
.Y(n_7628)
);

AND2x2_ASAP7_75t_L g7629 ( 
.A(n_7373),
.B(n_7510),
.Y(n_7629)
);

AND2x2_ASAP7_75t_L g7630 ( 
.A(n_7373),
.B(n_6936),
.Y(n_7630)
);

INVx1_ASAP7_75t_L g7631 ( 
.A(n_7359),
.Y(n_7631)
);

AND2x2_ASAP7_75t_L g7632 ( 
.A(n_7511),
.B(n_6936),
.Y(n_7632)
);

AND2x2_ASAP7_75t_L g7633 ( 
.A(n_7511),
.B(n_7488),
.Y(n_7633)
);

AND2x2_ASAP7_75t_L g7634 ( 
.A(n_7455),
.B(n_6936),
.Y(n_7634)
);

NAND2xp5_ASAP7_75t_L g7635 ( 
.A(n_7500),
.B(n_7108),
.Y(n_7635)
);

INVx1_ASAP7_75t_L g7636 ( 
.A(n_7258),
.Y(n_7636)
);

INVx2_ASAP7_75t_L g7637 ( 
.A(n_7444),
.Y(n_7637)
);

INVx1_ASAP7_75t_L g7638 ( 
.A(n_7262),
.Y(n_7638)
);

AND2x2_ASAP7_75t_L g7639 ( 
.A(n_7445),
.B(n_7447),
.Y(n_7639)
);

NAND2xp5_ASAP7_75t_SL g7640 ( 
.A(n_7323),
.B(n_7174),
.Y(n_7640)
);

OR2x2_ASAP7_75t_L g7641 ( 
.A(n_7453),
.B(n_7175),
.Y(n_7641)
);

NAND2xp5_ASAP7_75t_L g7642 ( 
.A(n_7503),
.B(n_7108),
.Y(n_7642)
);

AND2x2_ASAP7_75t_L g7643 ( 
.A(n_7260),
.B(n_6936),
.Y(n_7643)
);

HB1xp67_ASAP7_75t_L g7644 ( 
.A(n_7323),
.Y(n_7644)
);

INVx1_ASAP7_75t_L g7645 ( 
.A(n_7268),
.Y(n_7645)
);

INVx1_ASAP7_75t_L g7646 ( 
.A(n_7505),
.Y(n_7646)
);

NOR2xp33_ASAP7_75t_L g7647 ( 
.A(n_7454),
.B(n_7468),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_7348),
.Y(n_7648)
);

AND2x2_ASAP7_75t_L g7649 ( 
.A(n_7410),
.B(n_6936),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_7231),
.Y(n_7650)
);

AND2x4_ASAP7_75t_L g7651 ( 
.A(n_7410),
.B(n_7172),
.Y(n_7651)
);

INVx2_ASAP7_75t_L g7652 ( 
.A(n_7264),
.Y(n_7652)
);

INVx1_ASAP7_75t_L g7653 ( 
.A(n_7234),
.Y(n_7653)
);

NOR2xp33_ASAP7_75t_L g7654 ( 
.A(n_7452),
.B(n_6936),
.Y(n_7654)
);

AND2x2_ASAP7_75t_L g7655 ( 
.A(n_7413),
.B(n_6936),
.Y(n_7655)
);

AND2x2_ASAP7_75t_L g7656 ( 
.A(n_7413),
.B(n_7174),
.Y(n_7656)
);

OR2x2_ASAP7_75t_L g7657 ( 
.A(n_7296),
.B(n_7138),
.Y(n_7657)
);

AND2x2_ASAP7_75t_L g7658 ( 
.A(n_7393),
.B(n_7174),
.Y(n_7658)
);

INVx1_ASAP7_75t_L g7659 ( 
.A(n_7245),
.Y(n_7659)
);

INVx1_ASAP7_75t_L g7660 ( 
.A(n_7246),
.Y(n_7660)
);

AND2x2_ASAP7_75t_L g7661 ( 
.A(n_7467),
.B(n_7174),
.Y(n_7661)
);

INVx2_ASAP7_75t_L g7662 ( 
.A(n_7264),
.Y(n_7662)
);

AND2x2_ASAP7_75t_L g7663 ( 
.A(n_7507),
.B(n_7255),
.Y(n_7663)
);

OR2x2_ASAP7_75t_L g7664 ( 
.A(n_7371),
.B(n_7195),
.Y(n_7664)
);

INVx2_ASAP7_75t_L g7665 ( 
.A(n_7279),
.Y(n_7665)
);

AND2x2_ASAP7_75t_L g7666 ( 
.A(n_7470),
.B(n_7197),
.Y(n_7666)
);

AND2x2_ASAP7_75t_L g7667 ( 
.A(n_7509),
.B(n_7197),
.Y(n_7667)
);

INVx2_ASAP7_75t_L g7668 ( 
.A(n_7279),
.Y(n_7668)
);

INVx1_ASAP7_75t_L g7669 ( 
.A(n_7250),
.Y(n_7669)
);

AOI221xp5_ASAP7_75t_L g7670 ( 
.A1(n_7297),
.A2(n_7257),
.B1(n_7452),
.B2(n_7252),
.C(n_7259),
.Y(n_7670)
);

OR2x2_ASAP7_75t_L g7671 ( 
.A(n_7458),
.B(n_7109),
.Y(n_7671)
);

NAND2xp5_ASAP7_75t_L g7672 ( 
.A(n_7480),
.B(n_7108),
.Y(n_7672)
);

NAND2xp5_ASAP7_75t_L g7673 ( 
.A(n_7480),
.B(n_7114),
.Y(n_7673)
);

INVx1_ASAP7_75t_L g7674 ( 
.A(n_7253),
.Y(n_7674)
);

AND2x2_ASAP7_75t_L g7675 ( 
.A(n_7405),
.B(n_7197),
.Y(n_7675)
);

INVx1_ASAP7_75t_L g7676 ( 
.A(n_7254),
.Y(n_7676)
);

INVx1_ASAP7_75t_L g7677 ( 
.A(n_7281),
.Y(n_7677)
);

INVx1_ASAP7_75t_L g7678 ( 
.A(n_7282),
.Y(n_7678)
);

INVx1_ASAP7_75t_L g7679 ( 
.A(n_7283),
.Y(n_7679)
);

INVxp67_ASAP7_75t_L g7680 ( 
.A(n_7481),
.Y(n_7680)
);

INVx1_ASAP7_75t_SL g7681 ( 
.A(n_7368),
.Y(n_7681)
);

INVx2_ASAP7_75t_L g7682 ( 
.A(n_7307),
.Y(n_7682)
);

AND2x2_ASAP7_75t_L g7683 ( 
.A(n_7368),
.B(n_7225),
.Y(n_7683)
);

INVx1_ASAP7_75t_L g7684 ( 
.A(n_7290),
.Y(n_7684)
);

INVx1_ASAP7_75t_L g7685 ( 
.A(n_7292),
.Y(n_7685)
);

AND2x2_ASAP7_75t_L g7686 ( 
.A(n_7248),
.B(n_7225),
.Y(n_7686)
);

INVx1_ASAP7_75t_L g7687 ( 
.A(n_7295),
.Y(n_7687)
);

INVx1_ASAP7_75t_L g7688 ( 
.A(n_7440),
.Y(n_7688)
);

O2A1O1Ixp33_ASAP7_75t_L g7689 ( 
.A1(n_7252),
.A2(n_7025),
.B(n_7026),
.C(n_7021),
.Y(n_7689)
);

AND2x2_ASAP7_75t_L g7690 ( 
.A(n_7307),
.B(n_7225),
.Y(n_7690)
);

AND2x2_ASAP7_75t_L g7691 ( 
.A(n_7352),
.B(n_7225),
.Y(n_7691)
);

NAND2xp5_ASAP7_75t_L g7692 ( 
.A(n_7302),
.B(n_7114),
.Y(n_7692)
);

NAND2xp5_ASAP7_75t_L g7693 ( 
.A(n_7302),
.B(n_7114),
.Y(n_7693)
);

AND2x2_ASAP7_75t_L g7694 ( 
.A(n_7311),
.B(n_6904),
.Y(n_7694)
);

INVx2_ASAP7_75t_L g7695 ( 
.A(n_7441),
.Y(n_7695)
);

AND2x2_ASAP7_75t_L g7696 ( 
.A(n_7311),
.B(n_6904),
.Y(n_7696)
);

INVx3_ASAP7_75t_L g7697 ( 
.A(n_7441),
.Y(n_7697)
);

INVxp67_ASAP7_75t_SL g7698 ( 
.A(n_7259),
.Y(n_7698)
);

AND2x2_ASAP7_75t_L g7699 ( 
.A(n_7335),
.B(n_7172),
.Y(n_7699)
);

AND2x2_ASAP7_75t_L g7700 ( 
.A(n_7335),
.B(n_7172),
.Y(n_7700)
);

BUFx2_ASAP7_75t_L g7701 ( 
.A(n_7339),
.Y(n_7701)
);

OR2x2_ASAP7_75t_L g7702 ( 
.A(n_7498),
.B(n_7029),
.Y(n_7702)
);

INVx2_ASAP7_75t_L g7703 ( 
.A(n_7233),
.Y(n_7703)
);

INVx1_ASAP7_75t_L g7704 ( 
.A(n_7440),
.Y(n_7704)
);

INVx2_ASAP7_75t_L g7705 ( 
.A(n_7233),
.Y(n_7705)
);

AND2x2_ASAP7_75t_L g7706 ( 
.A(n_7251),
.B(n_7180),
.Y(n_7706)
);

NAND2xp5_ASAP7_75t_SL g7707 ( 
.A(n_7333),
.B(n_7180),
.Y(n_7707)
);

AND2x2_ASAP7_75t_L g7708 ( 
.A(n_7251),
.B(n_7180),
.Y(n_7708)
);

OR2x2_ASAP7_75t_L g7709 ( 
.A(n_7380),
.B(n_7030),
.Y(n_7709)
);

NAND2xp5_ASAP7_75t_L g7710 ( 
.A(n_7310),
.B(n_7145),
.Y(n_7710)
);

AND2x2_ASAP7_75t_L g7711 ( 
.A(n_7460),
.B(n_6918),
.Y(n_7711)
);

OR2x6_ASAP7_75t_L g7712 ( 
.A(n_7284),
.B(n_7145),
.Y(n_7712)
);

INVx1_ASAP7_75t_L g7713 ( 
.A(n_7446),
.Y(n_7713)
);

AND2x2_ASAP7_75t_L g7714 ( 
.A(n_7229),
.B(n_7023),
.Y(n_7714)
);

INVx2_ASAP7_75t_L g7715 ( 
.A(n_7241),
.Y(n_7715)
);

OR2x2_ASAP7_75t_L g7716 ( 
.A(n_7380),
.B(n_7031),
.Y(n_7716)
);

AND2x2_ASAP7_75t_L g7717 ( 
.A(n_7425),
.B(n_7133),
.Y(n_7717)
);

INVx1_ASAP7_75t_L g7718 ( 
.A(n_7446),
.Y(n_7718)
);

INVx1_ASAP7_75t_L g7719 ( 
.A(n_7456),
.Y(n_7719)
);

NOR2xp67_ASAP7_75t_L g7720 ( 
.A(n_7310),
.B(n_6699),
.Y(n_7720)
);

INVx1_ASAP7_75t_SL g7721 ( 
.A(n_7316),
.Y(n_7721)
);

AND2x2_ASAP7_75t_L g7722 ( 
.A(n_7426),
.B(n_7107),
.Y(n_7722)
);

AND2x2_ASAP7_75t_L g7723 ( 
.A(n_7427),
.B(n_7107),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_7456),
.Y(n_7724)
);

AND2x4_ASAP7_75t_SL g7725 ( 
.A(n_7237),
.B(n_7145),
.Y(n_7725)
);

INVx2_ASAP7_75t_L g7726 ( 
.A(n_7241),
.Y(n_7726)
);

AND2x2_ASAP7_75t_L g7727 ( 
.A(n_7472),
.B(n_7178),
.Y(n_7727)
);

NAND2xp5_ASAP7_75t_L g7728 ( 
.A(n_7276),
.B(n_7160),
.Y(n_7728)
);

AND2x2_ASAP7_75t_L g7729 ( 
.A(n_7475),
.B(n_7476),
.Y(n_7729)
);

BUFx2_ASAP7_75t_L g7730 ( 
.A(n_7276),
.Y(n_7730)
);

INVx2_ASAP7_75t_L g7731 ( 
.A(n_7247),
.Y(n_7731)
);

AOI22xp33_ASAP7_75t_L g7732 ( 
.A1(n_7257),
.A2(n_6591),
.B1(n_6624),
.B2(n_6617),
.Y(n_7732)
);

INVx1_ASAP7_75t_L g7733 ( 
.A(n_7469),
.Y(n_7733)
);

AND2x2_ASAP7_75t_L g7734 ( 
.A(n_7477),
.B(n_7178),
.Y(n_7734)
);

AND2x4_ASAP7_75t_L g7735 ( 
.A(n_7433),
.B(n_7160),
.Y(n_7735)
);

AND2x2_ASAP7_75t_L g7736 ( 
.A(n_7481),
.B(n_7181),
.Y(n_7736)
);

INVx1_ASAP7_75t_L g7737 ( 
.A(n_7469),
.Y(n_7737)
);

AND2x2_ASAP7_75t_L g7738 ( 
.A(n_7434),
.B(n_7181),
.Y(n_7738)
);

NAND2xp5_ASAP7_75t_L g7739 ( 
.A(n_7261),
.B(n_7160),
.Y(n_7739)
);

INVx2_ASAP7_75t_L g7740 ( 
.A(n_7247),
.Y(n_7740)
);

INVx2_ASAP7_75t_L g7741 ( 
.A(n_7300),
.Y(n_7741)
);

NAND2xp5_ASAP7_75t_SL g7742 ( 
.A(n_7333),
.B(n_7163),
.Y(n_7742)
);

INVx1_ASAP7_75t_L g7743 ( 
.A(n_7486),
.Y(n_7743)
);

NAND2xp5_ASAP7_75t_L g7744 ( 
.A(n_7267),
.B(n_7163),
.Y(n_7744)
);

INVx1_ASAP7_75t_SL g7745 ( 
.A(n_7305),
.Y(n_7745)
);

INVx1_ASAP7_75t_SL g7746 ( 
.A(n_7443),
.Y(n_7746)
);

AND2x2_ASAP7_75t_L g7747 ( 
.A(n_7434),
.B(n_7163),
.Y(n_7747)
);

INVx2_ASAP7_75t_L g7748 ( 
.A(n_7300),
.Y(n_7748)
);

AND2x2_ASAP7_75t_L g7749 ( 
.A(n_7462),
.B(n_7220),
.Y(n_7749)
);

NAND2xp5_ASAP7_75t_L g7750 ( 
.A(n_7273),
.B(n_7220),
.Y(n_7750)
);

NAND2xp5_ASAP7_75t_L g7751 ( 
.A(n_7274),
.B(n_7220),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_7486),
.Y(n_7752)
);

AND2x2_ASAP7_75t_L g7753 ( 
.A(n_7361),
.B(n_7042),
.Y(n_7753)
);

NOR5xp2_ASAP7_75t_SL g7754 ( 
.A(n_7478),
.B(n_6868),
.C(n_7057),
.D(n_7065),
.E(n_7043),
.Y(n_7754)
);

AND2x2_ASAP7_75t_L g7755 ( 
.A(n_7395),
.B(n_7066),
.Y(n_7755)
);

AND2x2_ASAP7_75t_L g7756 ( 
.A(n_7396),
.B(n_7069),
.Y(n_7756)
);

AND3x2_ASAP7_75t_L g7757 ( 
.A(n_7315),
.B(n_7045),
.C(n_7041),
.Y(n_7757)
);

NAND2xp5_ASAP7_75t_L g7758 ( 
.A(n_7293),
.B(n_7086),
.Y(n_7758)
);

AND2x2_ASAP7_75t_L g7759 ( 
.A(n_7435),
.B(n_7093),
.Y(n_7759)
);

INVx1_ASAP7_75t_L g7760 ( 
.A(n_7492),
.Y(n_7760)
);

NAND2xp5_ASAP7_75t_L g7761 ( 
.A(n_7269),
.B(n_7277),
.Y(n_7761)
);

INVx2_ASAP7_75t_L g7762 ( 
.A(n_7312),
.Y(n_7762)
);

INVx1_ASAP7_75t_L g7763 ( 
.A(n_7492),
.Y(n_7763)
);

INVx1_ASAP7_75t_L g7764 ( 
.A(n_7449),
.Y(n_7764)
);

AND2x2_ASAP7_75t_L g7765 ( 
.A(n_7466),
.B(n_7096),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_7451),
.Y(n_7766)
);

INVx2_ASAP7_75t_L g7767 ( 
.A(n_7312),
.Y(n_7767)
);

INVx2_ASAP7_75t_L g7768 ( 
.A(n_7430),
.Y(n_7768)
);

AND2x2_ASAP7_75t_L g7769 ( 
.A(n_7473),
.B(n_7115),
.Y(n_7769)
);

NOR2x1_ASAP7_75t_L g7770 ( 
.A(n_7315),
.B(n_7116),
.Y(n_7770)
);

AND2x2_ASAP7_75t_L g7771 ( 
.A(n_7580),
.B(n_7483),
.Y(n_7771)
);

XNOR2xp5_ASAP7_75t_L g7772 ( 
.A(n_7561),
.B(n_7240),
.Y(n_7772)
);

AND2x4_ASAP7_75t_L g7773 ( 
.A(n_7623),
.B(n_7485),
.Y(n_7773)
);

XNOR2xp5_ASAP7_75t_L g7774 ( 
.A(n_7569),
.B(n_7240),
.Y(n_7774)
);

AND2x2_ASAP7_75t_L g7775 ( 
.A(n_7580),
.B(n_7490),
.Y(n_7775)
);

NAND2xp5_ASAP7_75t_L g7776 ( 
.A(n_7583),
.B(n_7301),
.Y(n_7776)
);

NAND3xp33_ASAP7_75t_SL g7777 ( 
.A(n_7670),
.B(n_7555),
.C(n_7516),
.Y(n_7777)
);

AND2x2_ASAP7_75t_L g7778 ( 
.A(n_7569),
.B(n_7390),
.Y(n_7778)
);

NAND4xp75_ASAP7_75t_L g7779 ( 
.A(n_7555),
.B(n_7317),
.C(n_7230),
.D(n_7342),
.Y(n_7779)
);

AND2x2_ASAP7_75t_L g7780 ( 
.A(n_7573),
.B(n_7390),
.Y(n_7780)
);

XNOR2x2_ASAP7_75t_L g7781 ( 
.A(n_7541),
.B(n_7317),
.Y(n_7781)
);

INVx2_ASAP7_75t_L g7782 ( 
.A(n_7623),
.Y(n_7782)
);

INVx1_ASAP7_75t_L g7783 ( 
.A(n_7757),
.Y(n_7783)
);

NOR2xp33_ASAP7_75t_L g7784 ( 
.A(n_7538),
.B(n_7416),
.Y(n_7784)
);

BUFx2_ASAP7_75t_L g7785 ( 
.A(n_7712),
.Y(n_7785)
);

NAND2xp5_ASAP7_75t_L g7786 ( 
.A(n_7583),
.B(n_7303),
.Y(n_7786)
);

BUFx2_ASAP7_75t_L g7787 ( 
.A(n_7712),
.Y(n_7787)
);

INVx1_ASAP7_75t_L g7788 ( 
.A(n_7757),
.Y(n_7788)
);

AND2x2_ASAP7_75t_L g7789 ( 
.A(n_7573),
.B(n_7461),
.Y(n_7789)
);

NAND4xp75_ASAP7_75t_SL g7790 ( 
.A(n_7609),
.B(n_7461),
.C(n_7501),
.D(n_6369),
.Y(n_7790)
);

INVx4_ASAP7_75t_L g7791 ( 
.A(n_7549),
.Y(n_7791)
);

XNOR2xp5_ASAP7_75t_L g7792 ( 
.A(n_7746),
.B(n_7404),
.Y(n_7792)
);

NAND4xp75_ASAP7_75t_SL g7793 ( 
.A(n_7531),
.B(n_7501),
.C(n_6369),
.D(n_6491),
.Y(n_7793)
);

INVx1_ASAP7_75t_L g7794 ( 
.A(n_7591),
.Y(n_7794)
);

NAND2xp5_ASAP7_75t_L g7795 ( 
.A(n_7729),
.B(n_7256),
.Y(n_7795)
);

AOI22xp5_ASAP7_75t_L g7796 ( 
.A1(n_7698),
.A2(n_7342),
.B1(n_7230),
.B2(n_7349),
.Y(n_7796)
);

XOR2x2_ASAP7_75t_L g7797 ( 
.A(n_7541),
.B(n_7349),
.Y(n_7797)
);

NAND4xp75_ASAP7_75t_L g7798 ( 
.A(n_7518),
.B(n_7499),
.C(n_7502),
.D(n_7496),
.Y(n_7798)
);

NAND4xp75_ASAP7_75t_L g7799 ( 
.A(n_7518),
.B(n_7562),
.C(n_7647),
.D(n_7599),
.Y(n_7799)
);

INVx1_ASAP7_75t_L g7800 ( 
.A(n_7550),
.Y(n_7800)
);

AND2x2_ASAP7_75t_L g7801 ( 
.A(n_7593),
.B(n_7416),
.Y(n_7801)
);

INVx1_ASAP7_75t_L g7802 ( 
.A(n_7515),
.Y(n_7802)
);

NAND4xp75_ASAP7_75t_L g7803 ( 
.A(n_7647),
.B(n_7398),
.C(n_7400),
.D(n_7386),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_7554),
.Y(n_7804)
);

OR2x2_ASAP7_75t_L g7805 ( 
.A(n_7532),
.B(n_7512),
.Y(n_7805)
);

INVx2_ASAP7_75t_L g7806 ( 
.A(n_7556),
.Y(n_7806)
);

INVx2_ASAP7_75t_SL g7807 ( 
.A(n_7725),
.Y(n_7807)
);

BUFx2_ASAP7_75t_L g7808 ( 
.A(n_7712),
.Y(n_7808)
);

INVx1_ASAP7_75t_L g7809 ( 
.A(n_7611),
.Y(n_7809)
);

NAND3xp33_ASAP7_75t_L g7810 ( 
.A(n_7516),
.B(n_7442),
.C(n_7256),
.Y(n_7810)
);

NAND4xp75_ASAP7_75t_L g7811 ( 
.A(n_7661),
.B(n_7742),
.C(n_7570),
.D(n_7707),
.Y(n_7811)
);

INVx1_ASAP7_75t_L g7812 ( 
.A(n_7611),
.Y(n_7812)
);

AND2x2_ASAP7_75t_L g7813 ( 
.A(n_7593),
.B(n_7330),
.Y(n_7813)
);

AND2x2_ASAP7_75t_L g7814 ( 
.A(n_7639),
.B(n_7331),
.Y(n_7814)
);

XOR2xp5_ASAP7_75t_L g7815 ( 
.A(n_7610),
.B(n_7484),
.Y(n_7815)
);

AND2x2_ASAP7_75t_L g7816 ( 
.A(n_7535),
.B(n_7504),
.Y(n_7816)
);

INVx3_ASAP7_75t_L g7817 ( 
.A(n_7574),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_7644),
.Y(n_7818)
);

NAND4xp75_ASAP7_75t_L g7819 ( 
.A(n_7742),
.B(n_7372),
.C(n_7376),
.D(n_7365),
.Y(n_7819)
);

NOR3xp33_ASAP7_75t_L g7820 ( 
.A(n_7680),
.B(n_7442),
.C(n_7288),
.Y(n_7820)
);

OAI21xp5_ASAP7_75t_L g7821 ( 
.A1(n_7698),
.A2(n_7439),
.B(n_7424),
.Y(n_7821)
);

INVx1_ASAP7_75t_L g7822 ( 
.A(n_7644),
.Y(n_7822)
);

INVx1_ASAP7_75t_L g7823 ( 
.A(n_7581),
.Y(n_7823)
);

NAND4xp75_ASAP7_75t_L g7824 ( 
.A(n_7707),
.B(n_7383),
.C(n_7384),
.D(n_7377),
.Y(n_7824)
);

NAND2xp5_ASAP7_75t_L g7825 ( 
.A(n_7546),
.B(n_7430),
.Y(n_7825)
);

OAI22xp33_ASAP7_75t_L g7826 ( 
.A1(n_7543),
.A2(n_6227),
.B1(n_6351),
.B2(n_7287),
.Y(n_7826)
);

NAND4xp75_ASAP7_75t_SL g7827 ( 
.A(n_7604),
.B(n_6369),
.C(n_6491),
.D(n_6389),
.Y(n_7827)
);

INVx2_ASAP7_75t_SL g7828 ( 
.A(n_7725),
.Y(n_7828)
);

INVx2_ASAP7_75t_L g7829 ( 
.A(n_7556),
.Y(n_7829)
);

BUFx2_ASAP7_75t_L g7830 ( 
.A(n_7522),
.Y(n_7830)
);

AND2x4_ASAP7_75t_L g7831 ( 
.A(n_7556),
.B(n_7430),
.Y(n_7831)
);

AND2x2_ASAP7_75t_L g7832 ( 
.A(n_7558),
.B(n_7306),
.Y(n_7832)
);

INVx2_ASAP7_75t_L g7833 ( 
.A(n_7574),
.Y(n_7833)
);

NAND4xp75_ASAP7_75t_L g7834 ( 
.A(n_7747),
.B(n_7406),
.C(n_7408),
.D(n_7401),
.Y(n_7834)
);

OR2x2_ASAP7_75t_L g7835 ( 
.A(n_7601),
.B(n_7464),
.Y(n_7835)
);

INVx3_ASAP7_75t_L g7836 ( 
.A(n_7574),
.Y(n_7836)
);

AOI22xp5_ASAP7_75t_L g7837 ( 
.A1(n_7703),
.A2(n_6591),
.B1(n_6624),
.B2(n_6617),
.Y(n_7837)
);

INVx2_ASAP7_75t_L g7838 ( 
.A(n_7584),
.Y(n_7838)
);

NAND4xp75_ASAP7_75t_L g7839 ( 
.A(n_7699),
.B(n_7412),
.C(n_7414),
.D(n_7411),
.Y(n_7839)
);

NAND2xp5_ASAP7_75t_L g7840 ( 
.A(n_7536),
.B(n_7424),
.Y(n_7840)
);

XNOR2xp5_ASAP7_75t_L g7841 ( 
.A(n_7566),
.B(n_7474),
.Y(n_7841)
);

INVx3_ASAP7_75t_L g7842 ( 
.A(n_7584),
.Y(n_7842)
);

OR2x2_ASAP7_75t_L g7843 ( 
.A(n_7637),
.B(n_7439),
.Y(n_7843)
);

INVx1_ASAP7_75t_L g7844 ( 
.A(n_7637),
.Y(n_7844)
);

AND2x2_ASAP7_75t_L g7845 ( 
.A(n_7663),
.B(n_7320),
.Y(n_7845)
);

AND2x2_ASAP7_75t_L g7846 ( 
.A(n_7606),
.B(n_7328),
.Y(n_7846)
);

INVx1_ASAP7_75t_L g7847 ( 
.A(n_7522),
.Y(n_7847)
);

HB1xp67_ASAP7_75t_L g7848 ( 
.A(n_7578),
.Y(n_7848)
);

AND2x2_ASAP7_75t_L g7849 ( 
.A(n_7553),
.B(n_7329),
.Y(n_7849)
);

OR2x2_ASAP7_75t_L g7850 ( 
.A(n_7721),
.B(n_7493),
.Y(n_7850)
);

XNOR2xp5_ASAP7_75t_L g7851 ( 
.A(n_7564),
.B(n_7493),
.Y(n_7851)
);

AND2x4_ASAP7_75t_L g7852 ( 
.A(n_7651),
.B(n_7594),
.Y(n_7852)
);

INVx5_ASAP7_75t_L g7853 ( 
.A(n_7549),
.Y(n_7853)
);

NAND2xp5_ASAP7_75t_L g7854 ( 
.A(n_7594),
.B(n_7334),
.Y(n_7854)
);

INVx1_ASAP7_75t_L g7855 ( 
.A(n_7607),
.Y(n_7855)
);

INVx2_ASAP7_75t_SL g7856 ( 
.A(n_7651),
.Y(n_7856)
);

NAND4xp75_ASAP7_75t_L g7857 ( 
.A(n_7700),
.B(n_7423),
.C(n_7429),
.D(n_7421),
.Y(n_7857)
);

NAND4xp75_ASAP7_75t_L g7858 ( 
.A(n_7706),
.B(n_7437),
.C(n_7450),
.D(n_7432),
.Y(n_7858)
);

AND2x4_ASAP7_75t_L g7859 ( 
.A(n_7651),
.B(n_7497),
.Y(n_7859)
);

AND2x2_ASAP7_75t_L g7860 ( 
.A(n_7547),
.B(n_7344),
.Y(n_7860)
);

INVx2_ASAP7_75t_SL g7861 ( 
.A(n_7589),
.Y(n_7861)
);

NAND4xp75_ASAP7_75t_L g7862 ( 
.A(n_7708),
.B(n_7345),
.C(n_7360),
.D(n_7341),
.Y(n_7862)
);

NOR4xp25_ASAP7_75t_L g7863 ( 
.A(n_7597),
.B(n_7288),
.C(n_7289),
.D(n_7287),
.Y(n_7863)
);

NAND2xp5_ASAP7_75t_L g7864 ( 
.A(n_7594),
.B(n_7497),
.Y(n_7864)
);

AOI22xp5_ASAP7_75t_L g7865 ( 
.A1(n_7703),
.A2(n_6632),
.B1(n_6580),
.B2(n_6258),
.Y(n_7865)
);

AND2x2_ASAP7_75t_L g7866 ( 
.A(n_7589),
.B(n_7382),
.Y(n_7866)
);

OAI31xp33_ASAP7_75t_L g7867 ( 
.A1(n_7537),
.A2(n_6637),
.A3(n_7289),
.B(n_6621),
.Y(n_7867)
);

XOR2x2_ASAP7_75t_L g7868 ( 
.A(n_7641),
.B(n_7382),
.Y(n_7868)
);

NOR2x1_ASAP7_75t_SL g7869 ( 
.A(n_7549),
.B(n_6299),
.Y(n_7869)
);

INVx2_ASAP7_75t_L g7870 ( 
.A(n_7584),
.Y(n_7870)
);

AND2x2_ASAP7_75t_L g7871 ( 
.A(n_7525),
.B(n_7527),
.Y(n_7871)
);

INVx2_ASAP7_75t_L g7872 ( 
.A(n_7616),
.Y(n_7872)
);

NAND3xp33_ASAP7_75t_L g7873 ( 
.A(n_7537),
.B(n_7355),
.C(n_7353),
.Y(n_7873)
);

INVx1_ASAP7_75t_L g7874 ( 
.A(n_7581),
.Y(n_7874)
);

INVx1_ASAP7_75t_L g7875 ( 
.A(n_7582),
.Y(n_7875)
);

NAND4xp75_ASAP7_75t_SL g7876 ( 
.A(n_7608),
.B(n_7613),
.C(n_7602),
.D(n_7603),
.Y(n_7876)
);

NAND4xp75_ASAP7_75t_SL g7877 ( 
.A(n_7519),
.B(n_7513),
.C(n_7576),
.D(n_7534),
.Y(n_7877)
);

XOR2x2_ASAP7_75t_L g7878 ( 
.A(n_7530),
.B(n_7389),
.Y(n_7878)
);

AND2x2_ASAP7_75t_L g7879 ( 
.A(n_7513),
.B(n_7519),
.Y(n_7879)
);

NAND2xp5_ASAP7_75t_L g7880 ( 
.A(n_7616),
.B(n_7389),
.Y(n_7880)
);

BUFx2_ASAP7_75t_L g7881 ( 
.A(n_7544),
.Y(n_7881)
);

INVxp67_ASAP7_75t_L g7882 ( 
.A(n_7730),
.Y(n_7882)
);

BUFx2_ASAP7_75t_L g7883 ( 
.A(n_7735),
.Y(n_7883)
);

HB1xp67_ASAP7_75t_L g7884 ( 
.A(n_7616),
.Y(n_7884)
);

OA22x2_ASAP7_75t_L g7885 ( 
.A1(n_7551),
.A2(n_7508),
.B1(n_7506),
.B2(n_7122),
.Y(n_7885)
);

INVx1_ASAP7_75t_L g7886 ( 
.A(n_7582),
.Y(n_7886)
);

OR2x2_ASAP7_75t_L g7887 ( 
.A(n_7745),
.B(n_7407),
.Y(n_7887)
);

AND2x2_ASAP7_75t_L g7888 ( 
.A(n_7633),
.B(n_7407),
.Y(n_7888)
);

INVx1_ASAP7_75t_SL g7889 ( 
.A(n_7675),
.Y(n_7889)
);

XNOR2x2_ASAP7_75t_L g7890 ( 
.A(n_7622),
.B(n_7353),
.Y(n_7890)
);

NAND4xp75_ASAP7_75t_L g7891 ( 
.A(n_7643),
.B(n_7358),
.C(n_7379),
.D(n_7355),
.Y(n_7891)
);

INVx1_ASAP7_75t_L g7892 ( 
.A(n_7705),
.Y(n_7892)
);

AOI22xp5_ASAP7_75t_L g7893 ( 
.A1(n_7705),
.A2(n_6632),
.B1(n_6258),
.B2(n_6637),
.Y(n_7893)
);

AND4x1_ASAP7_75t_L g7894 ( 
.A(n_7548),
.B(n_7379),
.C(n_7358),
.D(n_7419),
.Y(n_7894)
);

INVx1_ASAP7_75t_L g7895 ( 
.A(n_7715),
.Y(n_7895)
);

XNOR2xp5_ASAP7_75t_L g7896 ( 
.A(n_7596),
.B(n_7419),
.Y(n_7896)
);

NAND4xp75_ASAP7_75t_SL g7897 ( 
.A(n_7576),
.B(n_6369),
.C(n_6389),
.D(n_6382),
.Y(n_7897)
);

XOR2xp5_ASAP7_75t_L g7898 ( 
.A(n_7552),
.B(n_6590),
.Y(n_7898)
);

OAI22x1_ASAP7_75t_L g7899 ( 
.A1(n_7551),
.A2(n_7124),
.B1(n_7125),
.B2(n_7119),
.Y(n_7899)
);

NAND3xp33_ASAP7_75t_L g7900 ( 
.A(n_7597),
.B(n_7146),
.C(n_7142),
.Y(n_7900)
);

AND2x2_ASAP7_75t_SL g7901 ( 
.A(n_7624),
.B(n_7147),
.Y(n_7901)
);

INVx2_ASAP7_75t_SL g7902 ( 
.A(n_7735),
.Y(n_7902)
);

XNOR2xp5_ASAP7_75t_L g7903 ( 
.A(n_7629),
.B(n_7150),
.Y(n_7903)
);

NAND2xp5_ASAP7_75t_SL g7904 ( 
.A(n_7735),
.B(n_5951),
.Y(n_7904)
);

NOR2xp33_ASAP7_75t_L g7905 ( 
.A(n_7538),
.B(n_7151),
.Y(n_7905)
);

INVx1_ASAP7_75t_L g7906 ( 
.A(n_7715),
.Y(n_7906)
);

INVx2_ASAP7_75t_SL g7907 ( 
.A(n_7694),
.Y(n_7907)
);

INVx1_ASAP7_75t_L g7908 ( 
.A(n_7726),
.Y(n_7908)
);

AND2x4_ASAP7_75t_L g7909 ( 
.A(n_7626),
.B(n_7155),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_7726),
.Y(n_7910)
);

XNOR2x2_ASAP7_75t_L g7911 ( 
.A(n_7622),
.B(n_7158),
.Y(n_7911)
);

XOR2x2_ASAP7_75t_L g7912 ( 
.A(n_7533),
.B(n_7640),
.Y(n_7912)
);

INVx5_ASAP7_75t_L g7913 ( 
.A(n_7697),
.Y(n_7913)
);

NAND4xp75_ASAP7_75t_SL g7914 ( 
.A(n_7667),
.B(n_6405),
.C(n_6510),
.D(n_6413),
.Y(n_7914)
);

AND2x2_ASAP7_75t_L g7915 ( 
.A(n_7658),
.B(n_7173),
.Y(n_7915)
);

OR2x2_ASAP7_75t_L g7916 ( 
.A(n_7571),
.B(n_7563),
.Y(n_7916)
);

OR3x1_ASAP7_75t_L g7917 ( 
.A(n_7565),
.B(n_6656),
.C(n_6642),
.Y(n_7917)
);

INVx1_ASAP7_75t_SL g7918 ( 
.A(n_7696),
.Y(n_7918)
);

XNOR2xp5_ASAP7_75t_L g7919 ( 
.A(n_7617),
.B(n_7177),
.Y(n_7919)
);

AND2x2_ASAP7_75t_L g7920 ( 
.A(n_7681),
.B(n_7179),
.Y(n_7920)
);

INVx2_ASAP7_75t_L g7921 ( 
.A(n_7626),
.Y(n_7921)
);

INVx1_ASAP7_75t_L g7922 ( 
.A(n_7521),
.Y(n_7922)
);

NAND4xp75_ASAP7_75t_SL g7923 ( 
.A(n_7749),
.B(n_6405),
.C(n_6510),
.D(n_6413),
.Y(n_7923)
);

INVx4_ASAP7_75t_L g7924 ( 
.A(n_7697),
.Y(n_7924)
);

NAND2xp5_ASAP7_75t_L g7925 ( 
.A(n_7626),
.B(n_7187),
.Y(n_7925)
);

XNOR2xp5_ASAP7_75t_L g7926 ( 
.A(n_7529),
.B(n_7190),
.Y(n_7926)
);

INVx1_ASAP7_75t_L g7927 ( 
.A(n_7524),
.Y(n_7927)
);

BUFx2_ASAP7_75t_L g7928 ( 
.A(n_7697),
.Y(n_7928)
);

NAND2xp5_ASAP7_75t_L g7929 ( 
.A(n_7682),
.B(n_7193),
.Y(n_7929)
);

NAND4xp75_ASAP7_75t_L g7930 ( 
.A(n_7736),
.B(n_7710),
.C(n_7634),
.D(n_7728),
.Y(n_7930)
);

XNOR2x2_ASAP7_75t_L g7931 ( 
.A(n_7640),
.B(n_7201),
.Y(n_7931)
);

INVx1_ASAP7_75t_L g7932 ( 
.A(n_7607),
.Y(n_7932)
);

INVx2_ASAP7_75t_L g7933 ( 
.A(n_7540),
.Y(n_7933)
);

AND2x2_ASAP7_75t_L g7934 ( 
.A(n_7666),
.B(n_7207),
.Y(n_7934)
);

INVx2_ASAP7_75t_L g7935 ( 
.A(n_7540),
.Y(n_7935)
);

NAND4xp75_ASAP7_75t_SL g7936 ( 
.A(n_7656),
.B(n_6413),
.C(n_6398),
.D(n_6354),
.Y(n_7936)
);

AOI22xp33_ASAP7_75t_L g7937 ( 
.A1(n_7732),
.A2(n_6897),
.B1(n_6621),
.B2(n_6501),
.Y(n_7937)
);

NAND2xp5_ASAP7_75t_L g7938 ( 
.A(n_7682),
.B(n_7211),
.Y(n_7938)
);

INVx3_ASAP7_75t_L g7939 ( 
.A(n_7540),
.Y(n_7939)
);

AO22x2_ASAP7_75t_L g7940 ( 
.A1(n_7568),
.A2(n_6980),
.B1(n_6995),
.B2(n_6952),
.Y(n_7940)
);

NOR4xp25_ASAP7_75t_L g7941 ( 
.A(n_7689),
.B(n_7215),
.C(n_7224),
.D(n_7212),
.Y(n_7941)
);

NAND4xp75_ASAP7_75t_L g7942 ( 
.A(n_7770),
.B(n_7005),
.C(n_7011),
.D(n_7000),
.Y(n_7942)
);

AND2x2_ASAP7_75t_L g7943 ( 
.A(n_7614),
.B(n_6657),
.Y(n_7943)
);

AND2x2_ASAP7_75t_L g7944 ( 
.A(n_7614),
.B(n_6665),
.Y(n_7944)
);

AND2x2_ASAP7_75t_L g7945 ( 
.A(n_7727),
.B(n_6679),
.Y(n_7945)
);

OR2x2_ASAP7_75t_L g7946 ( 
.A(n_7618),
.B(n_6681),
.Y(n_7946)
);

INVx1_ASAP7_75t_L g7947 ( 
.A(n_7612),
.Y(n_7947)
);

XNOR2xp5_ASAP7_75t_L g7948 ( 
.A(n_7646),
.B(n_6686),
.Y(n_7948)
);

NAND3xp33_ASAP7_75t_L g7949 ( 
.A(n_7557),
.B(n_6692),
.C(n_6690),
.Y(n_7949)
);

AND2x2_ASAP7_75t_L g7950 ( 
.A(n_7727),
.B(n_6701),
.Y(n_7950)
);

XNOR2x2_ASAP7_75t_L g7951 ( 
.A(n_7734),
.B(n_7013),
.Y(n_7951)
);

NAND2xp5_ASAP7_75t_L g7952 ( 
.A(n_7695),
.B(n_6458),
.Y(n_7952)
);

NAND4xp75_ASAP7_75t_L g7953 ( 
.A(n_7739),
.B(n_7020),
.C(n_7045),
.D(n_7041),
.Y(n_7953)
);

INVx3_ASAP7_75t_L g7954 ( 
.A(n_7612),
.Y(n_7954)
);

BUFx2_ASAP7_75t_L g7955 ( 
.A(n_7557),
.Y(n_7955)
);

NAND4xp75_ASAP7_75t_L g7956 ( 
.A(n_7744),
.B(n_7072),
.C(n_7088),
.D(n_7059),
.Y(n_7956)
);

INVx2_ASAP7_75t_SL g7957 ( 
.A(n_7686),
.Y(n_7957)
);

HB1xp67_ASAP7_75t_L g7958 ( 
.A(n_7701),
.Y(n_7958)
);

AND2x2_ASAP7_75t_L g7959 ( 
.A(n_7695),
.B(n_6068),
.Y(n_7959)
);

XNOR2xp5_ASAP7_75t_L g7960 ( 
.A(n_7526),
.B(n_7579),
.Y(n_7960)
);

INVx2_ASAP7_75t_L g7961 ( 
.A(n_7683),
.Y(n_7961)
);

INVx1_ASAP7_75t_L g7962 ( 
.A(n_7702),
.Y(n_7962)
);

NOR3xp33_ASAP7_75t_L g7963 ( 
.A(n_7680),
.B(n_7127),
.C(n_7118),
.Y(n_7963)
);

INVx1_ASAP7_75t_L g7964 ( 
.A(n_7577),
.Y(n_7964)
);

AND2x2_ASAP7_75t_L g7965 ( 
.A(n_7690),
.B(n_6077),
.Y(n_7965)
);

AND4x1_ASAP7_75t_L g7966 ( 
.A(n_7598),
.B(n_6476),
.C(n_5377),
.D(n_5310),
.Y(n_7966)
);

XNOR2xp5_ASAP7_75t_L g7967 ( 
.A(n_7567),
.B(n_6235),
.Y(n_7967)
);

AND2x2_ASAP7_75t_L g7968 ( 
.A(n_7691),
.B(n_6086),
.Y(n_7968)
);

NOR3xp33_ASAP7_75t_L g7969 ( 
.A(n_7750),
.B(n_7127),
.C(n_7118),
.Y(n_7969)
);

BUFx3_ASAP7_75t_L g7970 ( 
.A(n_7523),
.Y(n_7970)
);

INVx1_ASAP7_75t_L g7971 ( 
.A(n_7559),
.Y(n_7971)
);

AND2x2_ASAP7_75t_L g7972 ( 
.A(n_7648),
.B(n_6097),
.Y(n_7972)
);

INVx1_ASAP7_75t_L g7973 ( 
.A(n_7559),
.Y(n_7973)
);

NAND2xp5_ASAP7_75t_L g7974 ( 
.A(n_7753),
.B(n_7755),
.Y(n_7974)
);

INVx1_ASAP7_75t_L g7975 ( 
.A(n_7560),
.Y(n_7975)
);

NAND2xp5_ASAP7_75t_L g7976 ( 
.A(n_7753),
.B(n_6458),
.Y(n_7976)
);

NAND4xp75_ASAP7_75t_L g7977 ( 
.A(n_7751),
.B(n_7072),
.C(n_7088),
.D(n_7059),
.Y(n_7977)
);

AND2x2_ASAP7_75t_L g7978 ( 
.A(n_7714),
.B(n_6594),
.Y(n_7978)
);

NAND4xp75_ASAP7_75t_L g7979 ( 
.A(n_7720),
.B(n_7100),
.C(n_7105),
.D(n_7089),
.Y(n_7979)
);

INVx1_ASAP7_75t_L g7980 ( 
.A(n_7560),
.Y(n_7980)
);

NAND4xp75_ASAP7_75t_L g7981 ( 
.A(n_7738),
.B(n_7100),
.C(n_7105),
.D(n_7089),
.Y(n_7981)
);

NAND3xp33_ASAP7_75t_SL g7982 ( 
.A(n_7689),
.B(n_6855),
.C(n_6649),
.Y(n_7982)
);

OR2x2_ASAP7_75t_L g7983 ( 
.A(n_7587),
.B(n_6876),
.Y(n_7983)
);

INVx2_ASAP7_75t_SL g7984 ( 
.A(n_7717),
.Y(n_7984)
);

XNOR2xp5_ASAP7_75t_L g7985 ( 
.A(n_7657),
.B(n_6235),
.Y(n_7985)
);

INVx3_ASAP7_75t_L g7986 ( 
.A(n_7762),
.Y(n_7986)
);

INVx2_ASAP7_75t_L g7987 ( 
.A(n_7717),
.Y(n_7987)
);

AND2x4_ASAP7_75t_L g7988 ( 
.A(n_7649),
.B(n_6506),
.Y(n_7988)
);

AND2x2_ASAP7_75t_L g7989 ( 
.A(n_7789),
.B(n_7711),
.Y(n_7989)
);

INVxp67_ASAP7_75t_L g7990 ( 
.A(n_7883),
.Y(n_7990)
);

INVx1_ASAP7_75t_L g7991 ( 
.A(n_7928),
.Y(n_7991)
);

INVx1_ASAP7_75t_L g7992 ( 
.A(n_7884),
.Y(n_7992)
);

AND2x2_ASAP7_75t_L g7993 ( 
.A(n_7871),
.B(n_7655),
.Y(n_7993)
);

NOR2x1_ASAP7_75t_SL g7994 ( 
.A(n_7853),
.B(n_7762),
.Y(n_7994)
);

AND2x2_ASAP7_75t_L g7995 ( 
.A(n_7879),
.B(n_7630),
.Y(n_7995)
);

AND2x2_ASAP7_75t_L g7996 ( 
.A(n_7780),
.B(n_7632),
.Y(n_7996)
);

OR2x2_ASAP7_75t_L g7997 ( 
.A(n_7974),
.B(n_7664),
.Y(n_7997)
);

NAND2xp5_ASAP7_75t_L g7998 ( 
.A(n_7796),
.B(n_7600),
.Y(n_7998)
);

AND2x2_ASAP7_75t_L g7999 ( 
.A(n_7778),
.B(n_7722),
.Y(n_7999)
);

INVx1_ASAP7_75t_L g8000 ( 
.A(n_7940),
.Y(n_8000)
);

NAND2xp5_ASAP7_75t_L g8001 ( 
.A(n_7779),
.B(n_7605),
.Y(n_8001)
);

OR2x2_ASAP7_75t_L g8002 ( 
.A(n_7805),
.B(n_7586),
.Y(n_8002)
);

NOR2xp33_ASAP7_75t_L g8003 ( 
.A(n_7791),
.B(n_7615),
.Y(n_8003)
);

AND2x2_ASAP7_75t_L g8004 ( 
.A(n_7801),
.B(n_7722),
.Y(n_8004)
);

AND2x2_ASAP7_75t_L g8005 ( 
.A(n_7813),
.B(n_7723),
.Y(n_8005)
);

NAND2xp5_ASAP7_75t_L g8006 ( 
.A(n_7863),
.B(n_7619),
.Y(n_8006)
);

INVx2_ASAP7_75t_L g8007 ( 
.A(n_7913),
.Y(n_8007)
);

INVx2_ASAP7_75t_L g8008 ( 
.A(n_7913),
.Y(n_8008)
);

NAND2xp5_ASAP7_75t_L g8009 ( 
.A(n_7797),
.B(n_7621),
.Y(n_8009)
);

O2A1O1Ixp33_ASAP7_75t_L g8010 ( 
.A1(n_7777),
.A2(n_7592),
.B(n_7590),
.C(n_7625),
.Y(n_8010)
);

NAND2xp5_ASAP7_75t_L g8011 ( 
.A(n_7940),
.B(n_7954),
.Y(n_8011)
);

INVx1_ASAP7_75t_SL g8012 ( 
.A(n_7781),
.Y(n_8012)
);

AND2x2_ASAP7_75t_L g8013 ( 
.A(n_7816),
.B(n_7723),
.Y(n_8013)
);

AND2x2_ASAP7_75t_L g8014 ( 
.A(n_7888),
.B(n_7765),
.Y(n_8014)
);

OR2x2_ASAP7_75t_L g8015 ( 
.A(n_7848),
.B(n_7671),
.Y(n_8015)
);

AND2x2_ASAP7_75t_L g8016 ( 
.A(n_7866),
.B(n_7755),
.Y(n_8016)
);

NAND2xp5_ASAP7_75t_L g8017 ( 
.A(n_7954),
.B(n_7627),
.Y(n_8017)
);

INVx1_ASAP7_75t_L g8018 ( 
.A(n_7792),
.Y(n_8018)
);

AOI22xp33_ASAP7_75t_L g8019 ( 
.A1(n_7810),
.A2(n_6897),
.B1(n_7732),
.B2(n_7588),
.Y(n_8019)
);

INVx2_ASAP7_75t_L g8020 ( 
.A(n_7913),
.Y(n_8020)
);

INVx1_ASAP7_75t_L g8021 ( 
.A(n_7830),
.Y(n_8021)
);

INVx1_ASAP7_75t_L g8022 ( 
.A(n_7815),
.Y(n_8022)
);

AND2x2_ASAP7_75t_L g8023 ( 
.A(n_7807),
.B(n_7828),
.Y(n_8023)
);

INVx1_ASAP7_75t_L g8024 ( 
.A(n_7924),
.Y(n_8024)
);

AND2x2_ASAP7_75t_L g8025 ( 
.A(n_7861),
.B(n_7756),
.Y(n_8025)
);

INVx1_ASAP7_75t_L g8026 ( 
.A(n_7924),
.Y(n_8026)
);

AND2x2_ASAP7_75t_L g8027 ( 
.A(n_7814),
.B(n_7756),
.Y(n_8027)
);

AND2x2_ASAP7_75t_L g8028 ( 
.A(n_7771),
.B(n_7759),
.Y(n_8028)
);

CKINVDCx16_ASAP7_75t_R g8029 ( 
.A(n_7970),
.Y(n_8029)
);

NAND2xp5_ASAP7_75t_L g8030 ( 
.A(n_7809),
.B(n_7628),
.Y(n_8030)
);

INVx2_ASAP7_75t_L g8031 ( 
.A(n_7817),
.Y(n_8031)
);

NAND2xp5_ASAP7_75t_L g8032 ( 
.A(n_7809),
.B(n_7631),
.Y(n_8032)
);

OR2x2_ASAP7_75t_L g8033 ( 
.A(n_7887),
.B(n_7688),
.Y(n_8033)
);

NAND2xp33_ASAP7_75t_L g8034 ( 
.A(n_7811),
.B(n_7635),
.Y(n_8034)
);

INVx1_ASAP7_75t_L g8035 ( 
.A(n_7817),
.Y(n_8035)
);

AND2x2_ASAP7_75t_L g8036 ( 
.A(n_7775),
.B(n_7759),
.Y(n_8036)
);

OR2x2_ASAP7_75t_L g8037 ( 
.A(n_7916),
.B(n_7704),
.Y(n_8037)
);

NAND2xp5_ASAP7_75t_L g8038 ( 
.A(n_7812),
.B(n_7517),
.Y(n_8038)
);

INVx1_ASAP7_75t_L g8039 ( 
.A(n_7836),
.Y(n_8039)
);

INVx2_ASAP7_75t_L g8040 ( 
.A(n_7836),
.Y(n_8040)
);

AND2x2_ASAP7_75t_L g8041 ( 
.A(n_7845),
.B(n_7769),
.Y(n_8041)
);

AND2x2_ASAP7_75t_L g8042 ( 
.A(n_7846),
.B(n_7769),
.Y(n_8042)
);

OR2x2_ASAP7_75t_L g8043 ( 
.A(n_7850),
.B(n_7713),
.Y(n_8043)
);

INVx2_ASAP7_75t_L g8044 ( 
.A(n_7842),
.Y(n_8044)
);

INVx1_ASAP7_75t_L g8045 ( 
.A(n_7842),
.Y(n_8045)
);

NAND2x1p5_ASAP7_75t_L g8046 ( 
.A(n_7853),
.B(n_7514),
.Y(n_8046)
);

NAND2xp5_ASAP7_75t_L g8047 ( 
.A(n_7812),
.B(n_7520),
.Y(n_8047)
);

INVx1_ASAP7_75t_L g8048 ( 
.A(n_7785),
.Y(n_8048)
);

OR2x2_ASAP7_75t_L g8049 ( 
.A(n_7794),
.B(n_7718),
.Y(n_8049)
);

INVx2_ASAP7_75t_L g8050 ( 
.A(n_7852),
.Y(n_8050)
);

INVxp67_ASAP7_75t_L g8051 ( 
.A(n_7955),
.Y(n_8051)
);

AND2x2_ASAP7_75t_L g8052 ( 
.A(n_7856),
.B(n_7642),
.Y(n_8052)
);

NAND2x1_ASAP7_75t_SL g8053 ( 
.A(n_7852),
.B(n_7575),
.Y(n_8053)
);

INVx2_ASAP7_75t_L g8054 ( 
.A(n_7853),
.Y(n_8054)
);

INVx1_ASAP7_75t_L g8055 ( 
.A(n_7787),
.Y(n_8055)
);

INVx1_ASAP7_75t_L g8056 ( 
.A(n_7808),
.Y(n_8056)
);

NAND2xp33_ASAP7_75t_R g8057 ( 
.A(n_7881),
.B(n_7754),
.Y(n_8057)
);

INVx1_ASAP7_75t_L g8058 ( 
.A(n_7818),
.Y(n_8058)
);

INVx1_ASAP7_75t_L g8059 ( 
.A(n_7818),
.Y(n_8059)
);

AND2x2_ASAP7_75t_L g8060 ( 
.A(n_7832),
.B(n_7719),
.Y(n_8060)
);

OR2x2_ASAP7_75t_L g8061 ( 
.A(n_7795),
.B(n_7724),
.Y(n_8061)
);

NAND2xp5_ASAP7_75t_L g8062 ( 
.A(n_7939),
.B(n_7598),
.Y(n_8062)
);

OR2x2_ASAP7_75t_L g8063 ( 
.A(n_7840),
.B(n_7733),
.Y(n_8063)
);

AND2x2_ASAP7_75t_L g8064 ( 
.A(n_7849),
.B(n_7737),
.Y(n_8064)
);

NAND3xp33_ASAP7_75t_SL g8065 ( 
.A(n_7820),
.B(n_7595),
.C(n_7585),
.Y(n_8065)
);

AND2x2_ASAP7_75t_L g8066 ( 
.A(n_7860),
.B(n_7743),
.Y(n_8066)
);

AND2x2_ASAP7_75t_L g8067 ( 
.A(n_7918),
.B(n_7752),
.Y(n_8067)
);

AND2x2_ASAP7_75t_L g8068 ( 
.A(n_7959),
.B(n_7760),
.Y(n_8068)
);

OR2x2_ASAP7_75t_L g8069 ( 
.A(n_7835),
.B(n_7763),
.Y(n_8069)
);

AND2x4_ASAP7_75t_L g8070 ( 
.A(n_7831),
.B(n_7764),
.Y(n_8070)
);

INVx1_ASAP7_75t_L g8071 ( 
.A(n_7822),
.Y(n_8071)
);

NAND2xp5_ASAP7_75t_L g8072 ( 
.A(n_7822),
.B(n_7528),
.Y(n_8072)
);

NOR2xp33_ASAP7_75t_L g8073 ( 
.A(n_7791),
.B(n_7831),
.Y(n_8073)
);

HB1xp67_ASAP7_75t_L g8074 ( 
.A(n_7890),
.Y(n_8074)
);

NAND2xp5_ASAP7_75t_L g8075 ( 
.A(n_7774),
.B(n_7539),
.Y(n_8075)
);

INVx2_ASAP7_75t_SL g8076 ( 
.A(n_7859),
.Y(n_8076)
);

INVx1_ASAP7_75t_L g8077 ( 
.A(n_7843),
.Y(n_8077)
);

INVx1_ASAP7_75t_L g8078 ( 
.A(n_7919),
.Y(n_8078)
);

NAND2xp5_ASAP7_75t_L g8079 ( 
.A(n_7939),
.B(n_7768),
.Y(n_8079)
);

INVxp67_ASAP7_75t_L g8080 ( 
.A(n_7859),
.Y(n_8080)
);

INVx1_ASAP7_75t_L g8081 ( 
.A(n_7958),
.Y(n_8081)
);

INVx1_ASAP7_75t_L g8082 ( 
.A(n_7880),
.Y(n_8082)
);

INVx1_ASAP7_75t_L g8083 ( 
.A(n_7864),
.Y(n_8083)
);

AND2x2_ASAP7_75t_L g8084 ( 
.A(n_7907),
.B(n_7766),
.Y(n_8084)
);

HB1xp67_ASAP7_75t_L g8085 ( 
.A(n_7841),
.Y(n_8085)
);

OR2x2_ASAP7_75t_SL g8086 ( 
.A(n_7982),
.B(n_7767),
.Y(n_8086)
);

INVx1_ASAP7_75t_SL g8087 ( 
.A(n_7911),
.Y(n_8087)
);

AND2x2_ASAP7_75t_L g8088 ( 
.A(n_7782),
.B(n_7767),
.Y(n_8088)
);

INVx3_ASAP7_75t_L g8089 ( 
.A(n_7773),
.Y(n_8089)
);

INVx2_ASAP7_75t_L g8090 ( 
.A(n_7902),
.Y(n_8090)
);

NAND2xp5_ASAP7_75t_L g8091 ( 
.A(n_7892),
.B(n_7542),
.Y(n_8091)
);

INVx1_ASAP7_75t_L g8092 ( 
.A(n_7872),
.Y(n_8092)
);

AND2x4_ASAP7_75t_L g8093 ( 
.A(n_7833),
.B(n_7768),
.Y(n_8093)
);

AND2x2_ASAP7_75t_L g8094 ( 
.A(n_7972),
.B(n_7731),
.Y(n_8094)
);

INVx1_ASAP7_75t_L g8095 ( 
.A(n_7921),
.Y(n_8095)
);

NOR2xp33_ASAP7_75t_L g8096 ( 
.A(n_7889),
.B(n_7672),
.Y(n_8096)
);

NAND2xp5_ASAP7_75t_SL g8097 ( 
.A(n_7901),
.B(n_7731),
.Y(n_8097)
);

INVx1_ASAP7_75t_L g8098 ( 
.A(n_7776),
.Y(n_8098)
);

NAND2xp5_ASAP7_75t_L g8099 ( 
.A(n_7892),
.B(n_7545),
.Y(n_8099)
);

OR2x2_ASAP7_75t_L g8100 ( 
.A(n_7786),
.B(n_7692),
.Y(n_8100)
);

INVx1_ASAP7_75t_SL g8101 ( 
.A(n_7931),
.Y(n_8101)
);

AND3x2_ASAP7_75t_L g8102 ( 
.A(n_7882),
.B(n_7592),
.C(n_7590),
.Y(n_8102)
);

OR2x2_ASAP7_75t_L g8103 ( 
.A(n_7804),
.B(n_7693),
.Y(n_8103)
);

AND2x2_ASAP7_75t_L g8104 ( 
.A(n_7968),
.B(n_7740),
.Y(n_8104)
);

NAND2xp5_ASAP7_75t_L g8105 ( 
.A(n_7895),
.B(n_7652),
.Y(n_8105)
);

AND2x2_ASAP7_75t_L g8106 ( 
.A(n_7978),
.B(n_7740),
.Y(n_8106)
);

AND2x2_ASAP7_75t_L g8107 ( 
.A(n_7800),
.B(n_7741),
.Y(n_8107)
);

INVx2_ASAP7_75t_L g8108 ( 
.A(n_7838),
.Y(n_8108)
);

AND2x2_ASAP7_75t_L g8109 ( 
.A(n_7806),
.B(n_7741),
.Y(n_8109)
);

NAND2xp5_ASAP7_75t_L g8110 ( 
.A(n_7895),
.B(n_7652),
.Y(n_8110)
);

INVx2_ASAP7_75t_L g8111 ( 
.A(n_7870),
.Y(n_8111)
);

INVx4_ASAP7_75t_L g8112 ( 
.A(n_7773),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_7896),
.Y(n_8113)
);

OR2x2_ASAP7_75t_L g8114 ( 
.A(n_7829),
.B(n_7620),
.Y(n_8114)
);

NAND2xp5_ASAP7_75t_L g8115 ( 
.A(n_7906),
.B(n_7908),
.Y(n_8115)
);

INVx2_ASAP7_75t_L g8116 ( 
.A(n_7986),
.Y(n_8116)
);

INVx1_ASAP7_75t_L g8117 ( 
.A(n_7986),
.Y(n_8117)
);

OR2x2_ASAP7_75t_L g8118 ( 
.A(n_7844),
.B(n_7761),
.Y(n_8118)
);

AOI22xp5_ASAP7_75t_L g8119 ( 
.A1(n_7799),
.A2(n_7588),
.B1(n_7572),
.B2(n_7654),
.Y(n_8119)
);

A2O1A1Ixp33_ASAP7_75t_L g8120 ( 
.A1(n_7867),
.A2(n_7572),
.B(n_7654),
.C(n_6130),
.Y(n_8120)
);

INVx2_ASAP7_75t_L g8121 ( 
.A(n_7984),
.Y(n_8121)
);

AND2x2_ASAP7_75t_L g8122 ( 
.A(n_7965),
.B(n_7748),
.Y(n_8122)
);

OR2x2_ASAP7_75t_L g8123 ( 
.A(n_7962),
.B(n_7673),
.Y(n_8123)
);

INVx1_ASAP7_75t_SL g8124 ( 
.A(n_7877),
.Y(n_8124)
);

AND2x2_ASAP7_75t_L g8125 ( 
.A(n_7920),
.B(n_7748),
.Y(n_8125)
);

AND2x2_ASAP7_75t_L g8126 ( 
.A(n_7987),
.B(n_7662),
.Y(n_8126)
);

NAND2xp5_ASAP7_75t_L g8127 ( 
.A(n_7851),
.B(n_7662),
.Y(n_8127)
);

AND2x2_ASAP7_75t_L g8128 ( 
.A(n_7988),
.B(n_7665),
.Y(n_8128)
);

INVx2_ASAP7_75t_L g8129 ( 
.A(n_7933),
.Y(n_8129)
);

AND2x2_ASAP7_75t_L g8130 ( 
.A(n_7988),
.B(n_7665),
.Y(n_8130)
);

NAND2x1p5_ASAP7_75t_L g8131 ( 
.A(n_7847),
.B(n_7668),
.Y(n_8131)
);

AND2x2_ASAP7_75t_L g8132 ( 
.A(n_7802),
.B(n_7668),
.Y(n_8132)
);

INVx1_ASAP7_75t_L g8133 ( 
.A(n_7932),
.Y(n_8133)
);

NAND2xp5_ASAP7_75t_L g8134 ( 
.A(n_7945),
.B(n_7677),
.Y(n_8134)
);

INVx2_ASAP7_75t_SL g8135 ( 
.A(n_7935),
.Y(n_8135)
);

AND2x2_ASAP7_75t_L g8136 ( 
.A(n_7957),
.B(n_7636),
.Y(n_8136)
);

OR2x2_ASAP7_75t_L g8137 ( 
.A(n_7854),
.B(n_7709),
.Y(n_8137)
);

INVxp67_ASAP7_75t_L g8138 ( 
.A(n_7824),
.Y(n_8138)
);

AND2x4_ASAP7_75t_L g8139 ( 
.A(n_7909),
.B(n_7638),
.Y(n_8139)
);

AND2x2_ASAP7_75t_L g8140 ( 
.A(n_7868),
.B(n_7645),
.Y(n_8140)
);

NAND2xp5_ASAP7_75t_L g8141 ( 
.A(n_7906),
.B(n_7678),
.Y(n_8141)
);

INVx1_ASAP7_75t_L g8142 ( 
.A(n_7932),
.Y(n_8142)
);

NAND2xp5_ASAP7_75t_L g8143 ( 
.A(n_7908),
.B(n_7679),
.Y(n_8143)
);

NAND2x1p5_ASAP7_75t_L g8144 ( 
.A(n_7961),
.B(n_7716),
.Y(n_8144)
);

INVx1_ASAP7_75t_L g8145 ( 
.A(n_7947),
.Y(n_8145)
);

NAND2xp5_ASAP7_75t_L g8146 ( 
.A(n_7910),
.B(n_7684),
.Y(n_8146)
);

INVx1_ASAP7_75t_L g8147 ( 
.A(n_7947),
.Y(n_8147)
);

INVx2_ASAP7_75t_L g8148 ( 
.A(n_7909),
.Y(n_8148)
);

AND2x2_ASAP7_75t_L g8149 ( 
.A(n_7878),
.B(n_7685),
.Y(n_8149)
);

OR2x2_ASAP7_75t_L g8150 ( 
.A(n_7873),
.B(n_7929),
.Y(n_8150)
);

INVx1_ASAP7_75t_L g8151 ( 
.A(n_7910),
.Y(n_8151)
);

NAND2xp5_ASAP7_75t_L g8152 ( 
.A(n_7772),
.B(n_7941),
.Y(n_8152)
);

OR2x2_ASAP7_75t_L g8153 ( 
.A(n_7938),
.B(n_7758),
.Y(n_8153)
);

AND2x2_ASAP7_75t_L g8154 ( 
.A(n_7934),
.B(n_7687),
.Y(n_8154)
);

INVx1_ASAP7_75t_L g8155 ( 
.A(n_7885),
.Y(n_8155)
);

INVx1_ASAP7_75t_L g8156 ( 
.A(n_7950),
.Y(n_8156)
);

OAI22xp5_ASAP7_75t_L g8157 ( 
.A1(n_7798),
.A2(n_7653),
.B1(n_7659),
.B2(n_7650),
.Y(n_8157)
);

AND2x2_ASAP7_75t_L g8158 ( 
.A(n_7915),
.B(n_7660),
.Y(n_8158)
);

INVx1_ASAP7_75t_L g8159 ( 
.A(n_7979),
.Y(n_8159)
);

NAND2xp5_ASAP7_75t_L g8160 ( 
.A(n_7783),
.B(n_7669),
.Y(n_8160)
);

INVxp67_ASAP7_75t_L g8161 ( 
.A(n_7819),
.Y(n_8161)
);

INVx2_ASAP7_75t_L g8162 ( 
.A(n_7839),
.Y(n_8162)
);

OR2x2_ASAP7_75t_L g8163 ( 
.A(n_7855),
.B(n_7674),
.Y(n_8163)
);

OR2x2_ASAP7_75t_L g8164 ( 
.A(n_7925),
.B(n_7946),
.Y(n_8164)
);

INVx1_ASAP7_75t_L g8165 ( 
.A(n_7917),
.Y(n_8165)
);

INVx1_ASAP7_75t_L g8166 ( 
.A(n_7943),
.Y(n_8166)
);

OR2x2_ASAP7_75t_L g8167 ( 
.A(n_7825),
.B(n_7676),
.Y(n_8167)
);

INVx1_ASAP7_75t_L g8168 ( 
.A(n_7944),
.Y(n_8168)
);

INVx1_ASAP7_75t_L g8169 ( 
.A(n_7956),
.Y(n_8169)
);

NAND2xp5_ASAP7_75t_L g8170 ( 
.A(n_7783),
.B(n_7106),
.Y(n_8170)
);

NAND2xp5_ASAP7_75t_L g8171 ( 
.A(n_7788),
.B(n_7106),
.Y(n_8171)
);

INVxp67_ASAP7_75t_L g8172 ( 
.A(n_7857),
.Y(n_8172)
);

AND2x2_ASAP7_75t_L g8173 ( 
.A(n_7960),
.B(n_6594),
.Y(n_8173)
);

HB1xp67_ASAP7_75t_L g8174 ( 
.A(n_7876),
.Y(n_8174)
);

AND2x2_ASAP7_75t_L g8175 ( 
.A(n_7912),
.B(n_6649),
.Y(n_8175)
);

OR2x2_ASAP7_75t_L g8176 ( 
.A(n_7821),
.B(n_6855),
.Y(n_8176)
);

OR2x2_ASAP7_75t_L g8177 ( 
.A(n_7900),
.B(n_6506),
.Y(n_8177)
);

INVx1_ASAP7_75t_L g8178 ( 
.A(n_7977),
.Y(n_8178)
);

INVx2_ASAP7_75t_L g8179 ( 
.A(n_7858),
.Y(n_8179)
);

NOR2x1_ASAP7_75t_L g8180 ( 
.A(n_7930),
.B(n_7117),
.Y(n_8180)
);

INVx1_ASAP7_75t_L g8181 ( 
.A(n_7926),
.Y(n_8181)
);

INVx1_ASAP7_75t_L g8182 ( 
.A(n_7981),
.Y(n_8182)
);

NOR2xp33_ASAP7_75t_L g8183 ( 
.A(n_7904),
.B(n_6075),
.Y(n_8183)
);

AND2x2_ASAP7_75t_L g8184 ( 
.A(n_7903),
.B(n_6502),
.Y(n_8184)
);

NAND2xp5_ASAP7_75t_L g8185 ( 
.A(n_7788),
.B(n_7117),
.Y(n_8185)
);

AND2x2_ASAP7_75t_L g8186 ( 
.A(n_7784),
.B(n_7894),
.Y(n_8186)
);

OR2x2_ASAP7_75t_L g8187 ( 
.A(n_7983),
.B(n_6506),
.Y(n_8187)
);

NAND2xp5_ASAP7_75t_L g8188 ( 
.A(n_7969),
.B(n_6475),
.Y(n_8188)
);

AND2x2_ASAP7_75t_L g8189 ( 
.A(n_7834),
.B(n_6502),
.Y(n_8189)
);

NAND2xp5_ASAP7_75t_L g8190 ( 
.A(n_8029),
.B(n_7891),
.Y(n_8190)
);

INVx1_ASAP7_75t_L g8191 ( 
.A(n_8089),
.Y(n_8191)
);

NAND2xp5_ASAP7_75t_L g8192 ( 
.A(n_8089),
.B(n_7985),
.Y(n_8192)
);

NOR2xp33_ASAP7_75t_L g8193 ( 
.A(n_8112),
.B(n_7967),
.Y(n_8193)
);

INVx2_ASAP7_75t_SL g8194 ( 
.A(n_8053),
.Y(n_8194)
);

INVx1_ASAP7_75t_SL g8195 ( 
.A(n_8012),
.Y(n_8195)
);

NAND2xp5_ASAP7_75t_L g8196 ( 
.A(n_8112),
.B(n_7948),
.Y(n_8196)
);

NAND2xp33_ASAP7_75t_L g8197 ( 
.A(n_8085),
.B(n_7862),
.Y(n_8197)
);

INVx1_ASAP7_75t_L g8198 ( 
.A(n_8016),
.Y(n_8198)
);

NAND2xp5_ASAP7_75t_L g8199 ( 
.A(n_8028),
.B(n_7803),
.Y(n_8199)
);

INVx1_ASAP7_75t_L g8200 ( 
.A(n_8036),
.Y(n_8200)
);

AND2x2_ASAP7_75t_L g8201 ( 
.A(n_8027),
.B(n_7905),
.Y(n_8201)
);

INVx1_ASAP7_75t_L g8202 ( 
.A(n_8042),
.Y(n_8202)
);

OR2x2_ASAP7_75t_L g8203 ( 
.A(n_8002),
.B(n_8015),
.Y(n_8203)
);

NAND2x1_ASAP7_75t_L g8204 ( 
.A(n_8041),
.B(n_7976),
.Y(n_8204)
);

OAI22xp5_ASAP7_75t_L g8205 ( 
.A1(n_8074),
.A2(n_7952),
.B1(n_7898),
.B2(n_7949),
.Y(n_8205)
);

INVx1_ASAP7_75t_L g8206 ( 
.A(n_8025),
.Y(n_8206)
);

OR2x2_ASAP7_75t_L g8207 ( 
.A(n_8087),
.B(n_7964),
.Y(n_8207)
);

INVx1_ASAP7_75t_L g8208 ( 
.A(n_8011),
.Y(n_8208)
);

INVx1_ASAP7_75t_L g8209 ( 
.A(n_8011),
.Y(n_8209)
);

OAI21xp33_ASAP7_75t_L g8210 ( 
.A1(n_8152),
.A2(n_8101),
.B(n_8087),
.Y(n_8210)
);

AND2x2_ASAP7_75t_L g8211 ( 
.A(n_8005),
.B(n_7899),
.Y(n_8211)
);

NOR2xp33_ASAP7_75t_L g8212 ( 
.A(n_8012),
.B(n_7953),
.Y(n_8212)
);

NAND4xp25_ASAP7_75t_L g8213 ( 
.A(n_8057),
.B(n_7823),
.C(n_7875),
.D(n_7874),
.Y(n_8213)
);

OAI32xp33_ASAP7_75t_L g8214 ( 
.A1(n_8101),
.A2(n_7874),
.A3(n_7886),
.B1(n_7875),
.B2(n_7823),
.Y(n_8214)
);

AND2x2_ASAP7_75t_L g8215 ( 
.A(n_8013),
.B(n_7869),
.Y(n_8215)
);

NAND2xp5_ASAP7_75t_L g8216 ( 
.A(n_8014),
.B(n_7963),
.Y(n_8216)
);

INVx1_ASAP7_75t_L g8217 ( 
.A(n_8144),
.Y(n_8217)
);

AND2x2_ASAP7_75t_L g8218 ( 
.A(n_7989),
.B(n_7922),
.Y(n_8218)
);

INVx1_ASAP7_75t_L g8219 ( 
.A(n_7997),
.Y(n_8219)
);

NAND2xp5_ASAP7_75t_L g8220 ( 
.A(n_8102),
.B(n_7942),
.Y(n_8220)
);

INVxp67_ASAP7_75t_SL g8221 ( 
.A(n_8180),
.Y(n_8221)
);

AND2x2_ASAP7_75t_L g8222 ( 
.A(n_7999),
.B(n_7922),
.Y(n_8222)
);

HB1xp67_ASAP7_75t_L g8223 ( 
.A(n_8004),
.Y(n_8223)
);

NOR2xp67_ASAP7_75t_SL g8224 ( 
.A(n_8022),
.B(n_7927),
.Y(n_8224)
);

INVx2_ASAP7_75t_L g8225 ( 
.A(n_8046),
.Y(n_8225)
);

INVx2_ASAP7_75t_L g8226 ( 
.A(n_7994),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_8115),
.Y(n_8227)
);

OAI22xp5_ASAP7_75t_L g8228 ( 
.A1(n_8138),
.A2(n_7927),
.B1(n_7886),
.B2(n_7826),
.Y(n_8228)
);

INVx2_ASAP7_75t_L g8229 ( 
.A(n_7995),
.Y(n_8229)
);

NAND2xp5_ASAP7_75t_L g8230 ( 
.A(n_8076),
.B(n_7971),
.Y(n_8230)
);

AND2x2_ASAP7_75t_L g8231 ( 
.A(n_7993),
.B(n_7966),
.Y(n_8231)
);

INVx1_ASAP7_75t_L g8232 ( 
.A(n_8115),
.Y(n_8232)
);

HB1xp67_ASAP7_75t_L g8233 ( 
.A(n_8125),
.Y(n_8233)
);

INVx1_ASAP7_75t_L g8234 ( 
.A(n_8158),
.Y(n_8234)
);

AND2x2_ASAP7_75t_L g8235 ( 
.A(n_8104),
.B(n_6255),
.Y(n_8235)
);

INVx1_ASAP7_75t_L g8236 ( 
.A(n_8105),
.Y(n_8236)
);

NAND2xp5_ASAP7_75t_SL g8237 ( 
.A(n_8139),
.B(n_7971),
.Y(n_8237)
);

AND2x2_ASAP7_75t_L g8238 ( 
.A(n_8122),
.B(n_6255),
.Y(n_8238)
);

AOI22xp5_ASAP7_75t_L g8239 ( 
.A1(n_8152),
.A2(n_7975),
.B1(n_7980),
.B2(n_7973),
.Y(n_8239)
);

HB1xp67_ASAP7_75t_L g8240 ( 
.A(n_8070),
.Y(n_8240)
);

INVx2_ASAP7_75t_L g8241 ( 
.A(n_8131),
.Y(n_8241)
);

AND2x2_ASAP7_75t_L g8242 ( 
.A(n_8094),
.B(n_6255),
.Y(n_8242)
);

HB1xp67_ASAP7_75t_L g8243 ( 
.A(n_8070),
.Y(n_8243)
);

HB1xp67_ASAP7_75t_L g8244 ( 
.A(n_7990),
.Y(n_8244)
);

INVx1_ASAP7_75t_SL g8245 ( 
.A(n_8037),
.Y(n_8245)
);

NAND2xp5_ASAP7_75t_L g8246 ( 
.A(n_8060),
.B(n_7973),
.Y(n_8246)
);

AND2x2_ASAP7_75t_L g8247 ( 
.A(n_8064),
.B(n_6294),
.Y(n_8247)
);

INVx1_ASAP7_75t_L g8248 ( 
.A(n_8105),
.Y(n_8248)
);

OR2x2_ASAP7_75t_L g8249 ( 
.A(n_8050),
.B(n_7951),
.Y(n_8249)
);

AND2x2_ASAP7_75t_L g8250 ( 
.A(n_8066),
.B(n_6294),
.Y(n_8250)
);

NAND2xp5_ASAP7_75t_L g8251 ( 
.A(n_8139),
.B(n_7975),
.Y(n_8251)
);

INVx1_ASAP7_75t_L g8252 ( 
.A(n_8110),
.Y(n_8252)
);

NAND2xp5_ASAP7_75t_L g8253 ( 
.A(n_8093),
.B(n_7980),
.Y(n_8253)
);

AND2x2_ASAP7_75t_L g8254 ( 
.A(n_8106),
.B(n_6506),
.Y(n_8254)
);

NOR2xp67_ASAP7_75t_L g8255 ( 
.A(n_8080),
.B(n_7865),
.Y(n_8255)
);

INVx2_ASAP7_75t_L g8256 ( 
.A(n_8164),
.Y(n_8256)
);

OR2x2_ASAP7_75t_L g8257 ( 
.A(n_8135),
.B(n_8033),
.Y(n_8257)
);

INVx1_ASAP7_75t_L g8258 ( 
.A(n_8110),
.Y(n_8258)
);

INVx1_ASAP7_75t_L g8259 ( 
.A(n_8154),
.Y(n_8259)
);

INVx1_ASAP7_75t_L g8260 ( 
.A(n_8126),
.Y(n_8260)
);

INVxp67_ASAP7_75t_SL g8261 ( 
.A(n_8034),
.Y(n_8261)
);

OAI211xp5_ASAP7_75t_SL g8262 ( 
.A1(n_8161),
.A2(n_7893),
.B(n_7754),
.C(n_7937),
.Y(n_8262)
);

NAND2x1_ASAP7_75t_L g8263 ( 
.A(n_8093),
.B(n_5931),
.Y(n_8263)
);

INVxp67_ASAP7_75t_L g8264 ( 
.A(n_8073),
.Y(n_8264)
);

INVx1_ASAP7_75t_L g8265 ( 
.A(n_8068),
.Y(n_8265)
);

OAI21xp33_ASAP7_75t_L g8266 ( 
.A1(n_8006),
.A2(n_7790),
.B(n_7837),
.Y(n_8266)
);

AND2x2_ASAP7_75t_L g8267 ( 
.A(n_8052),
.B(n_6106),
.Y(n_8267)
);

INVxp67_ASAP7_75t_L g8268 ( 
.A(n_8128),
.Y(n_8268)
);

NAND3xp33_ASAP7_75t_L g8269 ( 
.A(n_8006),
.B(n_7148),
.C(n_7143),
.Y(n_8269)
);

INVx2_ASAP7_75t_SL g8270 ( 
.A(n_8130),
.Y(n_8270)
);

INVx1_ASAP7_75t_L g8271 ( 
.A(n_8109),
.Y(n_8271)
);

NAND2xp5_ASAP7_75t_L g8272 ( 
.A(n_8116),
.B(n_7143),
.Y(n_8272)
);

INVx1_ASAP7_75t_L g8273 ( 
.A(n_8107),
.Y(n_8273)
);

INVx1_ASAP7_75t_L g8274 ( 
.A(n_8043),
.Y(n_8274)
);

NAND2xp5_ASAP7_75t_L g8275 ( 
.A(n_8077),
.B(n_7148),
.Y(n_8275)
);

INVx1_ASAP7_75t_L g8276 ( 
.A(n_8132),
.Y(n_8276)
);

INVx3_ASAP7_75t_L g8277 ( 
.A(n_8148),
.Y(n_8277)
);

INVxp67_ASAP7_75t_L g8278 ( 
.A(n_7996),
.Y(n_8278)
);

AND2x2_ASAP7_75t_L g8279 ( 
.A(n_8023),
.B(n_6106),
.Y(n_8279)
);

INVx1_ASAP7_75t_L g8280 ( 
.A(n_8017),
.Y(n_8280)
);

OR2x6_ASAP7_75t_L g8281 ( 
.A(n_8054),
.B(n_7169),
.Y(n_8281)
);

INVx2_ASAP7_75t_L g8282 ( 
.A(n_8153),
.Y(n_8282)
);

NAND2xp5_ASAP7_75t_L g8283 ( 
.A(n_8031),
.B(n_7169),
.Y(n_8283)
);

INVx2_ASAP7_75t_L g8284 ( 
.A(n_8069),
.Y(n_8284)
);

INVxp67_ASAP7_75t_SL g8285 ( 
.A(n_8075),
.Y(n_8285)
);

INVx1_ASAP7_75t_L g8286 ( 
.A(n_8017),
.Y(n_8286)
);

INVxp67_ASAP7_75t_SL g8287 ( 
.A(n_8075),
.Y(n_8287)
);

INVx1_ASAP7_75t_L g8288 ( 
.A(n_8067),
.Y(n_8288)
);

OR2x2_ASAP7_75t_L g8289 ( 
.A(n_8040),
.B(n_8044),
.Y(n_8289)
);

INVx1_ASAP7_75t_L g8290 ( 
.A(n_8084),
.Y(n_8290)
);

INVx1_ASAP7_75t_L g8291 ( 
.A(n_8079),
.Y(n_8291)
);

NAND2xp5_ASAP7_75t_L g8292 ( 
.A(n_8166),
.B(n_7186),
.Y(n_8292)
);

INVx1_ASAP7_75t_L g8293 ( 
.A(n_8000),
.Y(n_8293)
);

INVx1_ASAP7_75t_L g8294 ( 
.A(n_8127),
.Y(n_8294)
);

NAND2xp5_ASAP7_75t_SL g8295 ( 
.A(n_8124),
.B(n_5911),
.Y(n_8295)
);

NAND2xp5_ASAP7_75t_L g8296 ( 
.A(n_8168),
.B(n_7186),
.Y(n_8296)
);

NAND2xp33_ASAP7_75t_L g8297 ( 
.A(n_8124),
.B(n_5867),
.Y(n_8297)
);

INVx1_ASAP7_75t_L g8298 ( 
.A(n_8088),
.Y(n_8298)
);

INVx1_ASAP7_75t_L g8299 ( 
.A(n_8117),
.Y(n_8299)
);

AND2x2_ASAP7_75t_L g8300 ( 
.A(n_8175),
.B(n_6414),
.Y(n_8300)
);

AND2x2_ASAP7_75t_L g8301 ( 
.A(n_8173),
.B(n_6414),
.Y(n_8301)
);

AND2x2_ASAP7_75t_L g8302 ( 
.A(n_8186),
.B(n_5753),
.Y(n_8302)
);

INVx2_ASAP7_75t_L g8303 ( 
.A(n_8137),
.Y(n_8303)
);

OAI21xp5_ASAP7_75t_SL g8304 ( 
.A1(n_8001),
.A2(n_7793),
.B(n_7923),
.Y(n_8304)
);

NAND2xp5_ASAP7_75t_L g8305 ( 
.A(n_8156),
.B(n_7188),
.Y(n_8305)
);

AOI22xp5_ASAP7_75t_L g8306 ( 
.A1(n_8001),
.A2(n_7196),
.B1(n_7202),
.B2(n_7188),
.Y(n_8306)
);

OR2x2_ASAP7_75t_L g8307 ( 
.A(n_8018),
.B(n_6323),
.Y(n_8307)
);

NAND2xp5_ASAP7_75t_L g8308 ( 
.A(n_8090),
.B(n_7196),
.Y(n_8308)
);

NAND3xp33_ASAP7_75t_L g8309 ( 
.A(n_8119),
.B(n_7221),
.C(n_7202),
.Y(n_8309)
);

INVx1_ASAP7_75t_SL g8310 ( 
.A(n_8118),
.Y(n_8310)
);

A2O1A1Ixp33_ASAP7_75t_L g8311 ( 
.A1(n_8120),
.A2(n_8019),
.B(n_8178),
.C(n_8169),
.Y(n_8311)
);

AND2x2_ASAP7_75t_L g8312 ( 
.A(n_8184),
.B(n_8140),
.Y(n_8312)
);

INVx3_ASAP7_75t_L g8313 ( 
.A(n_8007),
.Y(n_8313)
);

INVx1_ASAP7_75t_L g8314 ( 
.A(n_8114),
.Y(n_8314)
);

AND2x2_ASAP7_75t_L g8315 ( 
.A(n_8149),
.B(n_5775),
.Y(n_8315)
);

INVx2_ASAP7_75t_L g8316 ( 
.A(n_8100),
.Y(n_8316)
);

INVx1_ASAP7_75t_L g8317 ( 
.A(n_8129),
.Y(n_8317)
);

NOR2xp33_ASAP7_75t_L g8318 ( 
.A(n_8051),
.B(n_5911),
.Y(n_8318)
);

OAI31xp33_ASAP7_75t_L g8319 ( 
.A1(n_8182),
.A2(n_7936),
.A3(n_6980),
.B(n_6995),
.Y(n_8319)
);

AND2x4_ASAP7_75t_L g8320 ( 
.A(n_7991),
.B(n_6160),
.Y(n_8320)
);

INVx2_ASAP7_75t_L g8321 ( 
.A(n_8061),
.Y(n_8321)
);

INVx2_ASAP7_75t_L g8322 ( 
.A(n_8049),
.Y(n_8322)
);

A2O1A1Ixp33_ASAP7_75t_R g8323 ( 
.A1(n_8189),
.A2(n_7914),
.B(n_7827),
.C(n_7897),
.Y(n_8323)
);

OR2x2_ASAP7_75t_L g8324 ( 
.A(n_8150),
.B(n_6334),
.Y(n_8324)
);

INVx2_ASAP7_75t_SL g8325 ( 
.A(n_8136),
.Y(n_8325)
);

AND2x2_ASAP7_75t_L g8326 ( 
.A(n_8174),
.B(n_6113),
.Y(n_8326)
);

INVxp67_ASAP7_75t_L g8327 ( 
.A(n_8096),
.Y(n_8327)
);

INVx1_ASAP7_75t_L g8328 ( 
.A(n_8108),
.Y(n_8328)
);

AND2x2_ASAP7_75t_L g8329 ( 
.A(n_8121),
.B(n_6090),
.Y(n_8329)
);

INVx2_ASAP7_75t_L g8330 ( 
.A(n_8111),
.Y(n_8330)
);

INVx1_ASAP7_75t_L g8331 ( 
.A(n_8091),
.Y(n_8331)
);

NAND2xp5_ASAP7_75t_L g8332 ( 
.A(n_8035),
.B(n_7221),
.Y(n_8332)
);

INVx1_ASAP7_75t_SL g8333 ( 
.A(n_8063),
.Y(n_8333)
);

AOI22xp5_ASAP7_75t_L g8334 ( 
.A1(n_8159),
.A2(n_7228),
.B1(n_7226),
.B2(n_7001),
.Y(n_8334)
);

OAI22xp5_ASAP7_75t_L g8335 ( 
.A1(n_8172),
.A2(n_6160),
.B1(n_6181),
.B2(n_6846),
.Y(n_8335)
);

NAND2xp5_ASAP7_75t_L g8336 ( 
.A(n_8039),
.B(n_7226),
.Y(n_8336)
);

INVx1_ASAP7_75t_L g8337 ( 
.A(n_8091),
.Y(n_8337)
);

NAND2xp5_ASAP7_75t_L g8338 ( 
.A(n_8045),
.B(n_7228),
.Y(n_8338)
);

NOR2x1_ASAP7_75t_L g8339 ( 
.A(n_8065),
.B(n_6952),
.Y(n_8339)
);

OAI22xp5_ASAP7_75t_L g8340 ( 
.A1(n_8086),
.A2(n_6181),
.B1(n_6846),
.B2(n_6075),
.Y(n_8340)
);

AND2x2_ASAP7_75t_L g8341 ( 
.A(n_8021),
.B(n_6181),
.Y(n_8341)
);

NAND2xp5_ASAP7_75t_L g8342 ( 
.A(n_7992),
.B(n_7001),
.Y(n_8342)
);

OAI22xp5_ASAP7_75t_L g8343 ( 
.A1(n_8162),
.A2(n_6181),
.B1(n_6075),
.B2(n_6009),
.Y(n_8343)
);

INVx2_ASAP7_75t_L g8344 ( 
.A(n_8163),
.Y(n_8344)
);

NAND2xp5_ASAP7_75t_L g8345 ( 
.A(n_8098),
.B(n_7003),
.Y(n_8345)
);

BUFx2_ASAP7_75t_L g8346 ( 
.A(n_8092),
.Y(n_8346)
);

NAND2x1p5_ASAP7_75t_L g8347 ( 
.A(n_8081),
.B(n_6075),
.Y(n_8347)
);

NAND2xp5_ASAP7_75t_L g8348 ( 
.A(n_8095),
.B(n_7003),
.Y(n_8348)
);

INVx1_ASAP7_75t_L g8349 ( 
.A(n_8099),
.Y(n_8349)
);

AOI211xp5_ASAP7_75t_L g8350 ( 
.A1(n_8157),
.A2(n_7004),
.B(n_7017),
.C(n_5669),
.Y(n_8350)
);

OR2x2_ASAP7_75t_L g8351 ( 
.A(n_8134),
.B(n_6334),
.Y(n_8351)
);

INVx1_ASAP7_75t_L g8352 ( 
.A(n_8099),
.Y(n_8352)
);

NOR2xp33_ASAP7_75t_L g8353 ( 
.A(n_8062),
.B(n_5911),
.Y(n_8353)
);

INVx2_ASAP7_75t_L g8354 ( 
.A(n_8008),
.Y(n_8354)
);

OR2x2_ASAP7_75t_L g8355 ( 
.A(n_8203),
.B(n_7998),
.Y(n_8355)
);

INVx1_ASAP7_75t_L g8356 ( 
.A(n_8223),
.Y(n_8356)
);

NAND2x1p5_ASAP7_75t_L g8357 ( 
.A(n_8257),
.B(n_8048),
.Y(n_8357)
);

NAND2x1p5_ASAP7_75t_L g8358 ( 
.A(n_8217),
.B(n_8055),
.Y(n_8358)
);

OR2x2_ASAP7_75t_L g8359 ( 
.A(n_8195),
.B(n_7998),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_8240),
.Y(n_8360)
);

INVx1_ASAP7_75t_L g8361 ( 
.A(n_8243),
.Y(n_8361)
);

AOI22xp5_ASAP7_75t_L g8362 ( 
.A1(n_8210),
.A2(n_8179),
.B1(n_8119),
.B2(n_8009),
.Y(n_8362)
);

OR2x2_ASAP7_75t_L g8363 ( 
.A(n_8195),
.B(n_8233),
.Y(n_8363)
);

AND2x2_ASAP7_75t_L g8364 ( 
.A(n_8218),
.B(n_8056),
.Y(n_8364)
);

BUFx2_ASAP7_75t_L g8365 ( 
.A(n_8222),
.Y(n_8365)
);

NAND2xp5_ASAP7_75t_L g8366 ( 
.A(n_8333),
.B(n_8003),
.Y(n_8366)
);

INVx1_ASAP7_75t_L g8367 ( 
.A(n_8253),
.Y(n_8367)
);

INVx2_ASAP7_75t_L g8368 ( 
.A(n_8316),
.Y(n_8368)
);

INVxp67_ASAP7_75t_L g8369 ( 
.A(n_8237),
.Y(n_8369)
);

NAND2xp5_ASAP7_75t_L g8370 ( 
.A(n_8333),
.B(n_8097),
.Y(n_8370)
);

NOR2xp33_ASAP7_75t_L g8371 ( 
.A(n_8245),
.B(n_8113),
.Y(n_8371)
);

INVx1_ASAP7_75t_L g8372 ( 
.A(n_8251),
.Y(n_8372)
);

NAND2xp33_ASAP7_75t_L g8373 ( 
.A(n_8194),
.B(n_8009),
.Y(n_8373)
);

NOR2xp33_ASAP7_75t_L g8374 ( 
.A(n_8310),
.B(n_8268),
.Y(n_8374)
);

NAND2xp5_ASAP7_75t_SL g8375 ( 
.A(n_8210),
.B(n_8157),
.Y(n_8375)
);

NOR2xp33_ASAP7_75t_L g8376 ( 
.A(n_8310),
.B(n_8123),
.Y(n_8376)
);

INVx1_ASAP7_75t_L g8377 ( 
.A(n_8246),
.Y(n_8377)
);

INVx1_ASAP7_75t_L g8378 ( 
.A(n_8346),
.Y(n_8378)
);

INVx2_ASAP7_75t_L g8379 ( 
.A(n_8321),
.Y(n_8379)
);

NOR2xp33_ASAP7_75t_L g8380 ( 
.A(n_8270),
.B(n_8285),
.Y(n_8380)
);

INVx1_ASAP7_75t_SL g8381 ( 
.A(n_8249),
.Y(n_8381)
);

NAND2xp5_ASAP7_75t_L g8382 ( 
.A(n_8277),
.B(n_8082),
.Y(n_8382)
);

AND2x2_ASAP7_75t_L g8383 ( 
.A(n_8201),
.B(n_8181),
.Y(n_8383)
);

INVx2_ASAP7_75t_L g8384 ( 
.A(n_8277),
.Y(n_8384)
);

AND2x2_ASAP7_75t_L g8385 ( 
.A(n_8235),
.B(n_8078),
.Y(n_8385)
);

INVx1_ASAP7_75t_L g8386 ( 
.A(n_8339),
.Y(n_8386)
);

INVx1_ASAP7_75t_L g8387 ( 
.A(n_8221),
.Y(n_8387)
);

NOR2xp33_ASAP7_75t_L g8388 ( 
.A(n_8287),
.B(n_8177),
.Y(n_8388)
);

INVx2_ASAP7_75t_SL g8389 ( 
.A(n_8238),
.Y(n_8389)
);

AND2x2_ASAP7_75t_L g8390 ( 
.A(n_8211),
.B(n_8155),
.Y(n_8390)
);

INVx1_ASAP7_75t_L g8391 ( 
.A(n_8271),
.Y(n_8391)
);

INVx1_ASAP7_75t_L g8392 ( 
.A(n_8273),
.Y(n_8392)
);

AND2x2_ASAP7_75t_L g8393 ( 
.A(n_8242),
.B(n_8183),
.Y(n_8393)
);

INVx1_ASAP7_75t_L g8394 ( 
.A(n_8207),
.Y(n_8394)
);

NAND2xp5_ASAP7_75t_L g8395 ( 
.A(n_8261),
.B(n_8083),
.Y(n_8395)
);

INVx2_ASAP7_75t_L g8396 ( 
.A(n_8282),
.Y(n_8396)
);

OR2x6_ASAP7_75t_L g8397 ( 
.A(n_8226),
.B(n_8020),
.Y(n_8397)
);

OAI32xp33_ASAP7_75t_L g8398 ( 
.A1(n_8212),
.A2(n_8176),
.A3(n_8165),
.B1(n_8188),
.B2(n_8143),
.Y(n_8398)
);

INVx2_ASAP7_75t_L g8399 ( 
.A(n_8256),
.Y(n_8399)
);

NOR2xp33_ASAP7_75t_SL g8400 ( 
.A(n_8284),
.B(n_8010),
.Y(n_8400)
);

INVx2_ASAP7_75t_L g8401 ( 
.A(n_8303),
.Y(n_8401)
);

INVx2_ASAP7_75t_L g8402 ( 
.A(n_8281),
.Y(n_8402)
);

INVx1_ASAP7_75t_SL g8403 ( 
.A(n_8267),
.Y(n_8403)
);

NAND2xp5_ASAP7_75t_L g8404 ( 
.A(n_8219),
.B(n_8133),
.Y(n_8404)
);

AND2x2_ASAP7_75t_L g8405 ( 
.A(n_8279),
.B(n_8103),
.Y(n_8405)
);

NAND2xp5_ASAP7_75t_L g8406 ( 
.A(n_8314),
.B(n_8142),
.Y(n_8406)
);

NOR2x1_ASAP7_75t_L g8407 ( 
.A(n_8213),
.B(n_8151),
.Y(n_8407)
);

AND2x2_ASAP7_75t_L g8408 ( 
.A(n_8215),
.B(n_8167),
.Y(n_8408)
);

INVx1_ASAP7_75t_SL g8409 ( 
.A(n_8289),
.Y(n_8409)
);

INVx1_ASAP7_75t_SL g8410 ( 
.A(n_8312),
.Y(n_8410)
);

NAND2xp5_ASAP7_75t_L g8411 ( 
.A(n_8298),
.B(n_8145),
.Y(n_8411)
);

NOR2xp33_ASAP7_75t_L g8412 ( 
.A(n_8241),
.B(n_8288),
.Y(n_8412)
);

INVx1_ASAP7_75t_L g8413 ( 
.A(n_8281),
.Y(n_8413)
);

AOI221xp5_ASAP7_75t_L g8414 ( 
.A1(n_8266),
.A2(n_8146),
.B1(n_8143),
.B2(n_8141),
.C(n_8147),
.Y(n_8414)
);

INVx1_ASAP7_75t_L g8415 ( 
.A(n_8281),
.Y(n_8415)
);

AND2x2_ASAP7_75t_L g8416 ( 
.A(n_8247),
.B(n_8024),
.Y(n_8416)
);

INVx1_ASAP7_75t_L g8417 ( 
.A(n_8276),
.Y(n_8417)
);

OR2x2_ASAP7_75t_L g8418 ( 
.A(n_8229),
.B(n_8141),
.Y(n_8418)
);

NAND2xp5_ASAP7_75t_L g8419 ( 
.A(n_8278),
.B(n_8325),
.Y(n_8419)
);

NAND2xp5_ASAP7_75t_L g8420 ( 
.A(n_8198),
.B(n_8026),
.Y(n_8420)
);

NAND2xp33_ASAP7_75t_SL g8421 ( 
.A(n_8204),
.B(n_8146),
.Y(n_8421)
);

OR2x2_ASAP7_75t_L g8422 ( 
.A(n_8322),
.B(n_8038),
.Y(n_8422)
);

OR2x2_ASAP7_75t_L g8423 ( 
.A(n_8260),
.B(n_8038),
.Y(n_8423)
);

NAND2xp5_ASAP7_75t_L g8424 ( 
.A(n_8200),
.B(n_8058),
.Y(n_8424)
);

NAND2xp5_ASAP7_75t_L g8425 ( 
.A(n_8330),
.B(n_8059),
.Y(n_8425)
);

NOR4xp25_ASAP7_75t_L g8426 ( 
.A(n_8262),
.B(n_8171),
.C(n_8185),
.D(n_8170),
.Y(n_8426)
);

AND2x4_ASAP7_75t_L g8427 ( 
.A(n_8320),
.B(n_8071),
.Y(n_8427)
);

OR2x2_ASAP7_75t_L g8428 ( 
.A(n_8230),
.B(n_8047),
.Y(n_8428)
);

AOI21xp5_ASAP7_75t_SL g8429 ( 
.A1(n_8216),
.A2(n_8072),
.B(n_8047),
.Y(n_8429)
);

OR2x2_ASAP7_75t_L g8430 ( 
.A(n_8202),
.B(n_8072),
.Y(n_8430)
);

NAND2xp5_ASAP7_75t_L g8431 ( 
.A(n_8274),
.B(n_8030),
.Y(n_8431)
);

INVx1_ASAP7_75t_SL g8432 ( 
.A(n_8190),
.Y(n_8432)
);

HB1xp67_ASAP7_75t_L g8433 ( 
.A(n_8254),
.Y(n_8433)
);

NOR2xp33_ASAP7_75t_SL g8434 ( 
.A(n_8213),
.B(n_8030),
.Y(n_8434)
);

NAND3xp33_ASAP7_75t_L g8435 ( 
.A(n_8239),
.B(n_8032),
.C(n_8170),
.Y(n_8435)
);

INVx1_ASAP7_75t_L g8436 ( 
.A(n_8244),
.Y(n_8436)
);

OR2x2_ASAP7_75t_L g8437 ( 
.A(n_8344),
.B(n_8032),
.Y(n_8437)
);

NAND2xp5_ASAP7_75t_L g8438 ( 
.A(n_8265),
.B(n_8160),
.Y(n_8438)
);

INVx1_ASAP7_75t_L g8439 ( 
.A(n_8239),
.Y(n_8439)
);

BUFx2_ASAP7_75t_L g8440 ( 
.A(n_8347),
.Y(n_8440)
);

AND2x2_ASAP7_75t_SL g8441 ( 
.A(n_8197),
.B(n_8160),
.Y(n_8441)
);

NAND2xp5_ASAP7_75t_L g8442 ( 
.A(n_8313),
.B(n_8187),
.Y(n_8442)
);

HB1xp67_ASAP7_75t_L g8443 ( 
.A(n_8250),
.Y(n_8443)
);

AND2x4_ASAP7_75t_L g8444 ( 
.A(n_8320),
.B(n_8171),
.Y(n_8444)
);

OR2x2_ASAP7_75t_L g8445 ( 
.A(n_8234),
.B(n_8185),
.Y(n_8445)
);

AND2x2_ASAP7_75t_L g8446 ( 
.A(n_8315),
.B(n_6235),
.Y(n_8446)
);

INVxp67_ASAP7_75t_L g8447 ( 
.A(n_8224),
.Y(n_8447)
);

NAND2xp5_ASAP7_75t_L g8448 ( 
.A(n_8313),
.B(n_7004),
.Y(n_8448)
);

INVx1_ASAP7_75t_L g8449 ( 
.A(n_8317),
.Y(n_8449)
);

INVx1_ASAP7_75t_L g8450 ( 
.A(n_8328),
.Y(n_8450)
);

INVx1_ASAP7_75t_L g8451 ( 
.A(n_8236),
.Y(n_8451)
);

INVx1_ASAP7_75t_L g8452 ( 
.A(n_8248),
.Y(n_8452)
);

NAND2xp5_ASAP7_75t_L g8453 ( 
.A(n_8252),
.B(n_7017),
.Y(n_8453)
);

NAND2xp5_ASAP7_75t_L g8454 ( 
.A(n_8258),
.B(n_6641),
.Y(n_8454)
);

AND2x4_ASAP7_75t_L g8455 ( 
.A(n_8191),
.B(n_5975),
.Y(n_8455)
);

NAND2xp5_ASAP7_75t_L g8456 ( 
.A(n_8259),
.B(n_6641),
.Y(n_8456)
);

NAND2xp5_ASAP7_75t_L g8457 ( 
.A(n_8331),
.B(n_8337),
.Y(n_8457)
);

INVx1_ASAP7_75t_L g8458 ( 
.A(n_8309),
.Y(n_8458)
);

INVx2_ASAP7_75t_L g8459 ( 
.A(n_8263),
.Y(n_8459)
);

NAND2xp5_ASAP7_75t_L g8460 ( 
.A(n_8349),
.B(n_6644),
.Y(n_8460)
);

AOI31xp33_ASAP7_75t_L g8461 ( 
.A1(n_8327),
.A2(n_6047),
.A3(n_6651),
.B(n_6644),
.Y(n_8461)
);

INVx1_ASAP7_75t_L g8462 ( 
.A(n_8309),
.Y(n_8462)
);

INVx2_ASAP7_75t_L g8463 ( 
.A(n_8227),
.Y(n_8463)
);

INVxp67_ASAP7_75t_SL g8464 ( 
.A(n_8220),
.Y(n_8464)
);

OR2x2_ASAP7_75t_L g8465 ( 
.A(n_8290),
.B(n_6383),
.Y(n_8465)
);

AOI22xp5_ASAP7_75t_L g8466 ( 
.A1(n_8266),
.A2(n_6651),
.B1(n_6667),
.B2(n_6660),
.Y(n_8466)
);

NAND2xp5_ASAP7_75t_L g8467 ( 
.A(n_8352),
.B(n_8232),
.Y(n_8467)
);

NAND2xp5_ASAP7_75t_L g8468 ( 
.A(n_8206),
.B(n_6660),
.Y(n_8468)
);

INVx1_ASAP7_75t_L g8469 ( 
.A(n_8308),
.Y(n_8469)
);

AOI22xp5_ASAP7_75t_L g8470 ( 
.A1(n_8304),
.A2(n_6667),
.B1(n_6693),
.B2(n_6674),
.Y(n_8470)
);

INVx1_ASAP7_75t_L g8471 ( 
.A(n_8283),
.Y(n_8471)
);

OR2x2_ASAP7_75t_L g8472 ( 
.A(n_8196),
.B(n_6383),
.Y(n_8472)
);

AND2x2_ASAP7_75t_L g8473 ( 
.A(n_8302),
.B(n_8231),
.Y(n_8473)
);

NAND2xp5_ASAP7_75t_L g8474 ( 
.A(n_8341),
.B(n_6674),
.Y(n_8474)
);

AND2x2_ASAP7_75t_L g8475 ( 
.A(n_8326),
.B(n_6235),
.Y(n_8475)
);

OAI211xp5_ASAP7_75t_L g8476 ( 
.A1(n_8214),
.A2(n_5951),
.B(n_5867),
.C(n_5993),
.Y(n_8476)
);

NOR2xp33_ASAP7_75t_L g8477 ( 
.A(n_8264),
.B(n_6763),
.Y(n_8477)
);

NAND2xp5_ASAP7_75t_L g8478 ( 
.A(n_8291),
.B(n_6693),
.Y(n_8478)
);

AND2x2_ASAP7_75t_L g8479 ( 
.A(n_8329),
.B(n_6386),
.Y(n_8479)
);

NAND2xp5_ASAP7_75t_L g8480 ( 
.A(n_8280),
.B(n_6706),
.Y(n_8480)
);

AND2x2_ASAP7_75t_L g8481 ( 
.A(n_8294),
.B(n_6386),
.Y(n_8481)
);

AND2x2_ASAP7_75t_L g8482 ( 
.A(n_8300),
.B(n_6386),
.Y(n_8482)
);

INVx1_ASAP7_75t_L g8483 ( 
.A(n_8275),
.Y(n_8483)
);

AND2x2_ASAP7_75t_L g8484 ( 
.A(n_8225),
.B(n_6386),
.Y(n_8484)
);

NAND2xp5_ASAP7_75t_L g8485 ( 
.A(n_8286),
.B(n_6706),
.Y(n_8485)
);

INVx1_ASAP7_75t_L g8486 ( 
.A(n_8348),
.Y(n_8486)
);

INVxp67_ASAP7_75t_L g8487 ( 
.A(n_8193),
.Y(n_8487)
);

AND2x2_ASAP7_75t_L g8488 ( 
.A(n_8301),
.B(n_6477),
.Y(n_8488)
);

AND2x4_ASAP7_75t_SL g8489 ( 
.A(n_8354),
.B(n_5929),
.Y(n_8489)
);

AND2x2_ASAP7_75t_L g8490 ( 
.A(n_8353),
.B(n_6477),
.Y(n_8490)
);

INVx2_ASAP7_75t_SL g8491 ( 
.A(n_8295),
.Y(n_8491)
);

INVxp67_ASAP7_75t_L g8492 ( 
.A(n_8199),
.Y(n_8492)
);

AND2x2_ASAP7_75t_SL g8493 ( 
.A(n_8297),
.B(n_6712),
.Y(n_8493)
);

NAND2xp5_ASAP7_75t_L g8494 ( 
.A(n_8228),
.B(n_6712),
.Y(n_8494)
);

NAND2xp5_ASAP7_75t_L g8495 ( 
.A(n_8350),
.B(n_6719),
.Y(n_8495)
);

AND2x2_ASAP7_75t_L g8496 ( 
.A(n_8318),
.B(n_6477),
.Y(n_8496)
);

OR2x2_ASAP7_75t_L g8497 ( 
.A(n_8305),
.B(n_6398),
.Y(n_8497)
);

INVx2_ASAP7_75t_L g8498 ( 
.A(n_8351),
.Y(n_8498)
);

INVx2_ASAP7_75t_SL g8499 ( 
.A(n_8272),
.Y(n_8499)
);

INVx1_ASAP7_75t_SL g8500 ( 
.A(n_8192),
.Y(n_8500)
);

AOI22xp33_ASAP7_75t_L g8501 ( 
.A1(n_8269),
.A2(n_6448),
.B1(n_6501),
.B2(n_6497),
.Y(n_8501)
);

NOR2xp33_ASAP7_75t_L g8502 ( 
.A(n_8307),
.B(n_6719),
.Y(n_8502)
);

NAND2xp5_ASAP7_75t_L g8503 ( 
.A(n_8350),
.B(n_6720),
.Y(n_8503)
);

AND2x2_ASAP7_75t_L g8504 ( 
.A(n_8205),
.B(n_6477),
.Y(n_8504)
);

OAI221xp5_ASAP7_75t_L g8505 ( 
.A1(n_8434),
.A2(n_8319),
.B1(n_8304),
.B2(n_8311),
.C(n_8209),
.Y(n_8505)
);

INVx1_ASAP7_75t_L g8506 ( 
.A(n_8365),
.Y(n_8506)
);

NAND2xp5_ASAP7_75t_L g8507 ( 
.A(n_8409),
.B(n_8319),
.Y(n_8507)
);

AOI22xp5_ASAP7_75t_L g8508 ( 
.A1(n_8432),
.A2(n_8208),
.B1(n_8293),
.B2(n_8255),
.Y(n_8508)
);

NAND2xp5_ASAP7_75t_L g8509 ( 
.A(n_8409),
.B(n_8306),
.Y(n_8509)
);

NAND2xp5_ASAP7_75t_SL g8510 ( 
.A(n_8355),
.B(n_8340),
.Y(n_8510)
);

INVx1_ASAP7_75t_L g8511 ( 
.A(n_8359),
.Y(n_8511)
);

INVx1_ASAP7_75t_L g8512 ( 
.A(n_8363),
.Y(n_8512)
);

INVx2_ASAP7_75t_L g8513 ( 
.A(n_8357),
.Y(n_8513)
);

INVx1_ASAP7_75t_L g8514 ( 
.A(n_8364),
.Y(n_8514)
);

INVxp33_ASAP7_75t_L g8515 ( 
.A(n_8376),
.Y(n_8515)
);

NAND2xp5_ASAP7_75t_L g8516 ( 
.A(n_8410),
.B(n_8306),
.Y(n_8516)
);

INVx1_ASAP7_75t_L g8517 ( 
.A(n_8422),
.Y(n_8517)
);

OAI21xp33_ASAP7_75t_L g8518 ( 
.A1(n_8400),
.A2(n_8343),
.B(n_8296),
.Y(n_8518)
);

INVx2_ASAP7_75t_L g8519 ( 
.A(n_8437),
.Y(n_8519)
);

OR2x2_ASAP7_75t_L g8520 ( 
.A(n_8381),
.B(n_8292),
.Y(n_8520)
);

OAI22xp5_ASAP7_75t_L g8521 ( 
.A1(n_8362),
.A2(n_8299),
.B1(n_8342),
.B2(n_8324),
.Y(n_8521)
);

NAND2xp5_ASAP7_75t_SL g8522 ( 
.A(n_8441),
.B(n_8345),
.Y(n_8522)
);

OAI21xp33_ASAP7_75t_L g8523 ( 
.A1(n_8400),
.A2(n_8336),
.B(n_8332),
.Y(n_8523)
);

OAI21xp5_ASAP7_75t_L g8524 ( 
.A1(n_8369),
.A2(n_8269),
.B(n_8338),
.Y(n_8524)
);

NAND2xp5_ASAP7_75t_L g8525 ( 
.A(n_8444),
.B(n_8255),
.Y(n_8525)
);

INVx1_ASAP7_75t_L g8526 ( 
.A(n_8433),
.Y(n_8526)
);

OAI22xp33_ASAP7_75t_L g8527 ( 
.A1(n_8434),
.A2(n_8334),
.B1(n_8335),
.B2(n_8323),
.Y(n_8527)
);

INVx3_ASAP7_75t_L g8528 ( 
.A(n_8427),
.Y(n_8528)
);

NAND2xp5_ASAP7_75t_L g8529 ( 
.A(n_8444),
.B(n_8334),
.Y(n_8529)
);

AOI21xp5_ASAP7_75t_L g8530 ( 
.A1(n_8375),
.A2(n_6731),
.B(n_6720),
.Y(n_8530)
);

NAND2xp5_ASAP7_75t_L g8531 ( 
.A(n_8405),
.B(n_6731),
.Y(n_8531)
);

NAND2xp5_ASAP7_75t_L g8532 ( 
.A(n_8408),
.B(n_8384),
.Y(n_8532)
);

INVxp67_ASAP7_75t_SL g8533 ( 
.A(n_8366),
.Y(n_8533)
);

NAND2xp5_ASAP7_75t_L g8534 ( 
.A(n_8439),
.B(n_6736),
.Y(n_8534)
);

INVx1_ASAP7_75t_L g8535 ( 
.A(n_8443),
.Y(n_8535)
);

NAND2xp5_ASAP7_75t_L g8536 ( 
.A(n_8427),
.B(n_6736),
.Y(n_8536)
);

NAND4xp25_ASAP7_75t_SL g8537 ( 
.A(n_8362),
.B(n_6763),
.C(n_6766),
.D(n_6738),
.Y(n_8537)
);

NAND3xp33_ASAP7_75t_L g8538 ( 
.A(n_8373),
.B(n_6766),
.C(n_6738),
.Y(n_8538)
);

INVx1_ASAP7_75t_L g8539 ( 
.A(n_8418),
.Y(n_8539)
);

AOI21xp5_ASAP7_75t_L g8540 ( 
.A1(n_8421),
.A2(n_8435),
.B(n_8429),
.Y(n_8540)
);

INVx1_ASAP7_75t_L g8541 ( 
.A(n_8435),
.Y(n_8541)
);

INVx1_ASAP7_75t_L g8542 ( 
.A(n_8448),
.Y(n_8542)
);

XNOR2xp5_ASAP7_75t_L g8543 ( 
.A(n_8383),
.B(n_6207),
.Y(n_8543)
);

NAND2xp5_ASAP7_75t_L g8544 ( 
.A(n_8401),
.B(n_5929),
.Y(n_8544)
);

OAI22xp5_ASAP7_75t_L g8545 ( 
.A1(n_8447),
.A2(n_6853),
.B1(n_5929),
.B2(n_6009),
.Y(n_8545)
);

AND2x2_ASAP7_75t_L g8546 ( 
.A(n_8379),
.B(n_8399),
.Y(n_8546)
);

O2A1O1Ixp33_ASAP7_75t_L g8547 ( 
.A1(n_8458),
.A2(n_6133),
.B(n_6139),
.C(n_6136),
.Y(n_8547)
);

OAI31xp33_ASAP7_75t_L g8548 ( 
.A1(n_8386),
.A2(n_6133),
.A3(n_6139),
.B(n_6136),
.Y(n_8548)
);

INVx1_ASAP7_75t_SL g8549 ( 
.A(n_8428),
.Y(n_8549)
);

AOI21xp33_ASAP7_75t_L g8550 ( 
.A1(n_8388),
.A2(n_6448),
.B(n_6490),
.Y(n_8550)
);

AOI22xp5_ASAP7_75t_L g8551 ( 
.A1(n_8432),
.A2(n_6448),
.B1(n_6490),
.B2(n_6137),
.Y(n_8551)
);

HB1xp67_ASAP7_75t_L g8552 ( 
.A(n_8397),
.Y(n_8552)
);

OR2x2_ASAP7_75t_L g8553 ( 
.A(n_8370),
.B(n_6137),
.Y(n_8553)
);

INVx1_ASAP7_75t_L g8554 ( 
.A(n_8430),
.Y(n_8554)
);

NAND2xp5_ASAP7_75t_L g8555 ( 
.A(n_8403),
.B(n_5929),
.Y(n_8555)
);

AOI21xp33_ASAP7_75t_L g8556 ( 
.A1(n_8462),
.A2(n_6448),
.B(n_6490),
.Y(n_8556)
);

NAND2xp5_ASAP7_75t_L g8557 ( 
.A(n_8426),
.B(n_8368),
.Y(n_8557)
);

INVx1_ASAP7_75t_L g8558 ( 
.A(n_8382),
.Y(n_8558)
);

AOI21xp5_ASAP7_75t_L g8559 ( 
.A1(n_8407),
.A2(n_6137),
.B(n_6047),
.Y(n_8559)
);

AND2x2_ASAP7_75t_L g8560 ( 
.A(n_8394),
.B(n_6220),
.Y(n_8560)
);

INVxp67_ASAP7_75t_L g8561 ( 
.A(n_8380),
.Y(n_8561)
);

O2A1O1Ixp33_ASAP7_75t_L g8562 ( 
.A1(n_8426),
.A2(n_6151),
.B(n_6161),
.C(n_6158),
.Y(n_8562)
);

XNOR2x2_ASAP7_75t_L g8563 ( 
.A(n_8407),
.B(n_6130),
.Y(n_8563)
);

NOR2xp33_ASAP7_75t_L g8564 ( 
.A(n_8500),
.B(n_8378),
.Y(n_8564)
);

NAND2xp5_ASAP7_75t_L g8565 ( 
.A(n_8396),
.B(n_5975),
.Y(n_8565)
);

OAI22xp5_ASAP7_75t_L g8566 ( 
.A1(n_8360),
.A2(n_6853),
.B1(n_6129),
.B2(n_6194),
.Y(n_8566)
);

BUFx3_ASAP7_75t_L g8567 ( 
.A(n_8358),
.Y(n_8567)
);

AOI21xp5_ASAP7_75t_L g8568 ( 
.A1(n_8431),
.A2(n_6413),
.B(n_6398),
.Y(n_8568)
);

OR2x2_ASAP7_75t_L g8569 ( 
.A(n_8423),
.B(n_6398),
.Y(n_8569)
);

AND2x2_ASAP7_75t_L g8570 ( 
.A(n_8473),
.B(n_6220),
.Y(n_8570)
);

NAND2xp5_ASAP7_75t_L g8571 ( 
.A(n_8361),
.B(n_6775),
.Y(n_8571)
);

AOI31xp33_ASAP7_75t_SL g8572 ( 
.A1(n_8492),
.A2(n_6208),
.A3(n_6242),
.B(n_6175),
.Y(n_8572)
);

HB1xp67_ASAP7_75t_L g8573 ( 
.A(n_8397),
.Y(n_8573)
);

AOI32xp33_ASAP7_75t_L g8574 ( 
.A1(n_8390),
.A2(n_6119),
.A3(n_6151),
.B1(n_6161),
.B2(n_6158),
.Y(n_8574)
);

AND2x2_ASAP7_75t_L g8575 ( 
.A(n_8356),
.B(n_6220),
.Y(n_8575)
);

INVx1_ASAP7_75t_L g8576 ( 
.A(n_8445),
.Y(n_8576)
);

NOR4xp25_ASAP7_75t_SL g8577 ( 
.A(n_8440),
.B(n_6775),
.C(n_6490),
.D(n_6354),
.Y(n_8577)
);

INVx1_ASAP7_75t_L g8578 ( 
.A(n_8442),
.Y(n_8578)
);

INVx2_ASAP7_75t_L g8579 ( 
.A(n_8497),
.Y(n_8579)
);

OR2x2_ASAP7_75t_L g8580 ( 
.A(n_8397),
.B(n_6475),
.Y(n_8580)
);

AND2x2_ASAP7_75t_L g8581 ( 
.A(n_8416),
.B(n_6309),
.Y(n_8581)
);

NAND2xp5_ASAP7_75t_SL g8582 ( 
.A(n_8414),
.B(n_6475),
.Y(n_8582)
);

AOI221xp5_ASAP7_75t_L g8583 ( 
.A1(n_8413),
.A2(n_6171),
.B1(n_6168),
.B2(n_6353),
.C(n_6348),
.Y(n_8583)
);

INVx1_ASAP7_75t_L g8584 ( 
.A(n_8494),
.Y(n_8584)
);

OR2x2_ASAP7_75t_L g8585 ( 
.A(n_8438),
.B(n_6451),
.Y(n_8585)
);

INVxp67_ASAP7_75t_L g8586 ( 
.A(n_8374),
.Y(n_8586)
);

NAND2xp5_ASAP7_75t_L g8587 ( 
.A(n_8499),
.B(n_6775),
.Y(n_8587)
);

NAND2xp5_ASAP7_75t_L g8588 ( 
.A(n_8489),
.B(n_8493),
.Y(n_8588)
);

AOI21xp5_ASAP7_75t_L g8589 ( 
.A1(n_8404),
.A2(n_6171),
.B(n_6168),
.Y(n_8589)
);

NAND2xp5_ASAP7_75t_L g8590 ( 
.A(n_8481),
.B(n_5931),
.Y(n_8590)
);

NAND2xp5_ASAP7_75t_L g8591 ( 
.A(n_8389),
.B(n_5931),
.Y(n_8591)
);

AOI21xp5_ASAP7_75t_SL g8592 ( 
.A1(n_8371),
.A2(n_6207),
.B(n_6119),
.Y(n_8592)
);

NAND2xp5_ASAP7_75t_L g8593 ( 
.A(n_8491),
.B(n_5931),
.Y(n_8593)
);

NAND2xp5_ASAP7_75t_L g8594 ( 
.A(n_8488),
.B(n_5931),
.Y(n_8594)
);

OR2x2_ASAP7_75t_L g8595 ( 
.A(n_8425),
.B(n_8406),
.Y(n_8595)
);

INVx1_ASAP7_75t_SL g8596 ( 
.A(n_8393),
.Y(n_8596)
);

NAND2xp5_ASAP7_75t_L g8597 ( 
.A(n_8482),
.B(n_6437),
.Y(n_8597)
);

INVx1_ASAP7_75t_L g8598 ( 
.A(n_8402),
.Y(n_8598)
);

AOI21xp5_ASAP7_75t_L g8599 ( 
.A1(n_8395),
.A2(n_6353),
.B(n_6348),
.Y(n_8599)
);

AOI22xp5_ASAP7_75t_L g8600 ( 
.A1(n_8464),
.A2(n_8436),
.B1(n_8415),
.B2(n_8498),
.Y(n_8600)
);

INVxp67_ASAP7_75t_L g8601 ( 
.A(n_8502),
.Y(n_8601)
);

INVx1_ASAP7_75t_SL g8602 ( 
.A(n_8484),
.Y(n_8602)
);

AND2x4_ASAP7_75t_L g8603 ( 
.A(n_8455),
.B(n_8490),
.Y(n_8603)
);

INVx1_ASAP7_75t_L g8604 ( 
.A(n_8474),
.Y(n_8604)
);

AOI22xp5_ASAP7_75t_L g8605 ( 
.A1(n_8387),
.A2(n_6060),
.B1(n_6515),
.B2(n_6487),
.Y(n_8605)
);

AND2x2_ASAP7_75t_L g8606 ( 
.A(n_8385),
.B(n_6309),
.Y(n_8606)
);

OR2x2_ASAP7_75t_L g8607 ( 
.A(n_8424),
.B(n_6451),
.Y(n_8607)
);

O2A1O1Ixp33_ASAP7_75t_L g8608 ( 
.A1(n_8398),
.A2(n_6357),
.B(n_6368),
.C(n_6355),
.Y(n_8608)
);

INVx1_ASAP7_75t_L g8609 ( 
.A(n_8419),
.Y(n_8609)
);

AOI221xp5_ASAP7_75t_SL g8610 ( 
.A1(n_8372),
.A2(n_6368),
.B1(n_6395),
.B2(n_6357),
.C(n_6355),
.Y(n_8610)
);

INVx1_ASAP7_75t_L g8611 ( 
.A(n_8495),
.Y(n_8611)
);

BUFx6f_ASAP7_75t_L g8612 ( 
.A(n_8463),
.Y(n_8612)
);

AOI21xp5_ASAP7_75t_L g8613 ( 
.A1(n_8467),
.A2(n_6417),
.B(n_6395),
.Y(n_8613)
);

OAI21xp33_ASAP7_75t_SL g8614 ( 
.A1(n_8457),
.A2(n_8412),
.B(n_8411),
.Y(n_8614)
);

OAI22xp5_ASAP7_75t_L g8615 ( 
.A1(n_8377),
.A2(n_6129),
.B1(n_6194),
.B2(n_6172),
.Y(n_8615)
);

OAI22xp5_ASAP7_75t_L g8616 ( 
.A1(n_8367),
.A2(n_8391),
.B1(n_8417),
.B2(n_8392),
.Y(n_8616)
);

INVxp67_ASAP7_75t_L g8617 ( 
.A(n_8477),
.Y(n_8617)
);

OAI21xp33_ASAP7_75t_L g8618 ( 
.A1(n_8446),
.A2(n_5900),
.B(n_5993),
.Y(n_8618)
);

AOI22xp5_ASAP7_75t_L g8619 ( 
.A1(n_8496),
.A2(n_6060),
.B1(n_6515),
.B2(n_6487),
.Y(n_8619)
);

INVx1_ASAP7_75t_L g8620 ( 
.A(n_8503),
.Y(n_8620)
);

O2A1O1Ixp33_ASAP7_75t_L g8621 ( 
.A1(n_8487),
.A2(n_6418),
.B(n_6417),
.C(n_6513),
.Y(n_8621)
);

AOI22xp5_ASAP7_75t_L g8622 ( 
.A1(n_8469),
.A2(n_8483),
.B1(n_8471),
.B2(n_8479),
.Y(n_8622)
);

AND3x2_ASAP7_75t_L g8623 ( 
.A(n_8449),
.B(n_6451),
.C(n_6119),
.Y(n_8623)
);

INVx2_ASAP7_75t_L g8624 ( 
.A(n_8475),
.Y(n_8624)
);

NAND2xp5_ASAP7_75t_L g8625 ( 
.A(n_8455),
.B(n_6437),
.Y(n_8625)
);

NAND3xp33_ASAP7_75t_L g8626 ( 
.A(n_8450),
.B(n_6179),
.C(n_6175),
.Y(n_8626)
);

A2O1A1Ixp33_ASAP7_75t_L g8627 ( 
.A1(n_8470),
.A2(n_6418),
.B(n_6513),
.C(n_6179),
.Y(n_8627)
);

INVx1_ASAP7_75t_L g8628 ( 
.A(n_8453),
.Y(n_8628)
);

INVxp67_ASAP7_75t_L g8629 ( 
.A(n_8504),
.Y(n_8629)
);

INVx1_ASAP7_75t_L g8630 ( 
.A(n_8468),
.Y(n_8630)
);

INVx2_ASAP7_75t_L g8631 ( 
.A(n_8465),
.Y(n_8631)
);

OR2x2_ASAP7_75t_L g8632 ( 
.A(n_8456),
.B(n_6286),
.Y(n_8632)
);

INVx1_ASAP7_75t_L g8633 ( 
.A(n_8454),
.Y(n_8633)
);

OAI211xp5_ASAP7_75t_SL g8634 ( 
.A1(n_8505),
.A2(n_8451),
.B(n_8452),
.C(n_8486),
.Y(n_8634)
);

AOI21xp33_ASAP7_75t_L g8635 ( 
.A1(n_8525),
.A2(n_8485),
.B(n_8480),
.Y(n_8635)
);

NAND2xp5_ASAP7_75t_SL g8636 ( 
.A(n_8612),
.B(n_8528),
.Y(n_8636)
);

INVx1_ASAP7_75t_L g8637 ( 
.A(n_8528),
.Y(n_8637)
);

INVx1_ASAP7_75t_L g8638 ( 
.A(n_8552),
.Y(n_8638)
);

INVx1_ASAP7_75t_L g8639 ( 
.A(n_8573),
.Y(n_8639)
);

NAND2xp5_ASAP7_75t_L g8640 ( 
.A(n_8596),
.B(n_8461),
.Y(n_8640)
);

INVx1_ASAP7_75t_L g8641 ( 
.A(n_8529),
.Y(n_8641)
);

NAND2xp5_ASAP7_75t_L g8642 ( 
.A(n_8549),
.B(n_8470),
.Y(n_8642)
);

NAND2xp5_ASAP7_75t_L g8643 ( 
.A(n_8511),
.B(n_8466),
.Y(n_8643)
);

AOI22xp5_ASAP7_75t_L g8644 ( 
.A1(n_8541),
.A2(n_8466),
.B1(n_8460),
.B2(n_8478),
.Y(n_8644)
);

INVxp67_ASAP7_75t_L g8645 ( 
.A(n_8567),
.Y(n_8645)
);

INVx1_ASAP7_75t_L g8646 ( 
.A(n_8520),
.Y(n_8646)
);

INVx2_ASAP7_75t_SL g8647 ( 
.A(n_8612),
.Y(n_8647)
);

INVx1_ASAP7_75t_L g8648 ( 
.A(n_8546),
.Y(n_8648)
);

NOR2xp67_ASAP7_75t_L g8649 ( 
.A(n_8614),
.B(n_8420),
.Y(n_8649)
);

OAI22xp5_ASAP7_75t_L g8650 ( 
.A1(n_8595),
.A2(n_8472),
.B1(n_8459),
.B2(n_8501),
.Y(n_8650)
);

AOI22xp33_ASAP7_75t_L g8651 ( 
.A1(n_8556),
.A2(n_6182),
.B1(n_6208),
.B2(n_6204),
.Y(n_8651)
);

INVx1_ASAP7_75t_L g8652 ( 
.A(n_8509),
.Y(n_8652)
);

AOI32xp33_ASAP7_75t_L g8653 ( 
.A1(n_8515),
.A2(n_8476),
.A3(n_6129),
.B1(n_6194),
.B2(n_6172),
.Y(n_8653)
);

AND2x2_ASAP7_75t_L g8654 ( 
.A(n_8513),
.B(n_6309),
.Y(n_8654)
);

OAI22xp5_ASAP7_75t_SL g8655 ( 
.A1(n_8533),
.A2(n_5965),
.B1(n_6207),
.B2(n_6172),
.Y(n_8655)
);

NAND2xp5_ASAP7_75t_SL g8656 ( 
.A(n_8612),
.B(n_6089),
.Y(n_8656)
);

INVx1_ASAP7_75t_L g8657 ( 
.A(n_8532),
.Y(n_8657)
);

AOI32xp33_ASAP7_75t_L g8658 ( 
.A1(n_8527),
.A2(n_6211),
.A3(n_6212),
.B1(n_6204),
.B2(n_6182),
.Y(n_8658)
);

INVx1_ASAP7_75t_L g8659 ( 
.A(n_8519),
.Y(n_8659)
);

INVx1_ASAP7_75t_L g8660 ( 
.A(n_8557),
.Y(n_8660)
);

OAI22xp5_ASAP7_75t_L g8661 ( 
.A1(n_8576),
.A2(n_6211),
.B1(n_6214),
.B2(n_6212),
.Y(n_8661)
);

INVx1_ASAP7_75t_L g8662 ( 
.A(n_8516),
.Y(n_8662)
);

AND2x2_ASAP7_75t_L g8663 ( 
.A(n_8570),
.B(n_6207),
.Y(n_8663)
);

INVx1_ASAP7_75t_L g8664 ( 
.A(n_8536),
.Y(n_8664)
);

NAND2xp5_ASAP7_75t_L g8665 ( 
.A(n_8540),
.B(n_6222),
.Y(n_8665)
);

AOI22xp5_ASAP7_75t_SL g8666 ( 
.A1(n_8517),
.A2(n_6060),
.B1(n_6061),
.B2(n_6044),
.Y(n_8666)
);

AOI221x1_ASAP7_75t_L g8667 ( 
.A1(n_8523),
.A2(n_6226),
.B1(n_6242),
.B2(n_6222),
.C(n_6214),
.Y(n_8667)
);

NAND2xp5_ASAP7_75t_L g8668 ( 
.A(n_8526),
.B(n_6271),
.Y(n_8668)
);

AND2x2_ASAP7_75t_L g8669 ( 
.A(n_8606),
.B(n_6060),
.Y(n_8669)
);

INVxp67_ASAP7_75t_L g8670 ( 
.A(n_8522),
.Y(n_8670)
);

INVx1_ASAP7_75t_L g8671 ( 
.A(n_8531),
.Y(n_8671)
);

INVx1_ASAP7_75t_L g8672 ( 
.A(n_8569),
.Y(n_8672)
);

NAND2xp5_ASAP7_75t_L g8673 ( 
.A(n_8539),
.B(n_6272),
.Y(n_8673)
);

OAI21xp5_ASAP7_75t_L g8674 ( 
.A1(n_8614),
.A2(n_8508),
.B(n_8564),
.Y(n_8674)
);

INVx1_ASAP7_75t_L g8675 ( 
.A(n_8514),
.Y(n_8675)
);

OAI31xp33_ASAP7_75t_L g8676 ( 
.A1(n_8507),
.A2(n_6241),
.A3(n_6251),
.B(n_6226),
.Y(n_8676)
);

CKINVDCx14_ASAP7_75t_R g8677 ( 
.A(n_8603),
.Y(n_8677)
);

INVx1_ASAP7_75t_L g8678 ( 
.A(n_8554),
.Y(n_8678)
);

INVx1_ASAP7_75t_L g8679 ( 
.A(n_8535),
.Y(n_8679)
);

INVx1_ASAP7_75t_L g8680 ( 
.A(n_8512),
.Y(n_8680)
);

AOI22xp5_ASAP7_75t_L g8681 ( 
.A1(n_8579),
.A2(n_6515),
.B1(n_6487),
.B2(n_6251),
.Y(n_8681)
);

INVx2_ASAP7_75t_L g8682 ( 
.A(n_8603),
.Y(n_8682)
);

OAI22xp33_ASAP7_75t_L g8683 ( 
.A1(n_8600),
.A2(n_6271),
.B1(n_6272),
.B2(n_6241),
.Y(n_8683)
);

O2A1O1Ixp5_ASAP7_75t_L g8684 ( 
.A1(n_8524),
.A2(n_6281),
.B(n_6289),
.C(n_6277),
.Y(n_8684)
);

INVxp33_ASAP7_75t_L g8685 ( 
.A(n_8543),
.Y(n_8685)
);

INVx1_ASAP7_75t_L g8686 ( 
.A(n_8506),
.Y(n_8686)
);

INVxp67_ASAP7_75t_SL g8687 ( 
.A(n_8510),
.Y(n_8687)
);

AOI22xp5_ASAP7_75t_L g8688 ( 
.A1(n_8631),
.A2(n_8571),
.B1(n_8620),
.B2(n_8611),
.Y(n_8688)
);

OAI22xp5_ASAP7_75t_L g8689 ( 
.A1(n_8558),
.A2(n_6281),
.B1(n_6289),
.B2(n_6277),
.Y(n_8689)
);

OAI21xp33_ASAP7_75t_SL g8690 ( 
.A1(n_8559),
.A2(n_6301),
.B(n_6291),
.Y(n_8690)
);

INVx1_ASAP7_75t_SL g8691 ( 
.A(n_8588),
.Y(n_8691)
);

NOR2x1_ASAP7_75t_L g8692 ( 
.A(n_8521),
.B(n_6419),
.Y(n_8692)
);

OAI21x1_ASAP7_75t_SL g8693 ( 
.A1(n_8563),
.A2(n_8530),
.B(n_8565),
.Y(n_8693)
);

INVx1_ASAP7_75t_L g8694 ( 
.A(n_8538),
.Y(n_8694)
);

AND2x4_ASAP7_75t_L g8695 ( 
.A(n_8578),
.B(n_6291),
.Y(n_8695)
);

INVx2_ASAP7_75t_L g8696 ( 
.A(n_8580),
.Y(n_8696)
);

INVx1_ASAP7_75t_L g8697 ( 
.A(n_8534),
.Y(n_8697)
);

AND2x2_ASAP7_75t_L g8698 ( 
.A(n_8581),
.B(n_5900),
.Y(n_8698)
);

INVx2_ASAP7_75t_L g8699 ( 
.A(n_8623),
.Y(n_8699)
);

NAND2xp5_ASAP7_75t_L g8700 ( 
.A(n_8560),
.B(n_6301),
.Y(n_8700)
);

INVx1_ASAP7_75t_L g8701 ( 
.A(n_8587),
.Y(n_8701)
);

INVx1_ASAP7_75t_L g8702 ( 
.A(n_8572),
.Y(n_8702)
);

AOI21xp5_ASAP7_75t_L g8703 ( 
.A1(n_8582),
.A2(n_6354),
.B(n_6419),
.Y(n_8703)
);

INVx1_ASAP7_75t_L g8704 ( 
.A(n_8555),
.Y(n_8704)
);

A2O1A1Ixp33_ASAP7_75t_L g8705 ( 
.A1(n_8568),
.A2(n_8553),
.B(n_8550),
.C(n_8551),
.Y(n_8705)
);

INVx1_ASAP7_75t_L g8706 ( 
.A(n_8625),
.Y(n_8706)
);

AND2x2_ASAP7_75t_L g8707 ( 
.A(n_8575),
.B(n_6354),
.Y(n_8707)
);

AOI322xp5_ASAP7_75t_L g8708 ( 
.A1(n_8604),
.A2(n_6303),
.A3(n_6324),
.B1(n_6347),
.B2(n_6316),
.C1(n_6330),
.C2(n_6109),
.Y(n_8708)
);

XNOR2x2_ASAP7_75t_L g8709 ( 
.A(n_8616),
.B(n_6286),
.Y(n_8709)
);

INVx2_ASAP7_75t_L g8710 ( 
.A(n_8585),
.Y(n_8710)
);

INVx1_ASAP7_75t_L g8711 ( 
.A(n_8624),
.Y(n_8711)
);

INVx1_ASAP7_75t_L g8712 ( 
.A(n_8544),
.Y(n_8712)
);

NAND2xp5_ASAP7_75t_L g8713 ( 
.A(n_8518),
.B(n_8628),
.Y(n_8713)
);

AOI221xp5_ASAP7_75t_L g8714 ( 
.A1(n_8545),
.A2(n_6316),
.B1(n_6347),
.B2(n_6324),
.C(n_6303),
.Y(n_8714)
);

NAND2xp5_ASAP7_75t_L g8715 ( 
.A(n_8586),
.B(n_6437),
.Y(n_8715)
);

OAI222xp33_ASAP7_75t_L g8716 ( 
.A1(n_8574),
.A2(n_5973),
.B1(n_5932),
.B2(n_5999),
.C1(n_5972),
.C2(n_5963),
.Y(n_8716)
);

INVx1_ASAP7_75t_L g8717 ( 
.A(n_8597),
.Y(n_8717)
);

INVx1_ASAP7_75t_L g8718 ( 
.A(n_8562),
.Y(n_8718)
);

AOI32xp33_ASAP7_75t_L g8719 ( 
.A1(n_8609),
.A2(n_6098),
.A3(n_6109),
.B1(n_6066),
.B2(n_6298),
.Y(n_8719)
);

INVx2_ASAP7_75t_L g8720 ( 
.A(n_8607),
.Y(n_8720)
);

AOI32xp33_ASAP7_75t_L g8721 ( 
.A1(n_8594),
.A2(n_6098),
.A3(n_6066),
.B1(n_6298),
.B2(n_5408),
.Y(n_8721)
);

AND2x2_ASAP7_75t_L g8722 ( 
.A(n_8561),
.B(n_6089),
.Y(n_8722)
);

AOI221xp5_ASAP7_75t_L g8723 ( 
.A1(n_8542),
.A2(n_6288),
.B1(n_6346),
.B2(n_6317),
.C(n_6365),
.Y(n_8723)
);

INVx1_ASAP7_75t_L g8724 ( 
.A(n_8622),
.Y(n_8724)
);

NOR2xp33_ASAP7_75t_L g8725 ( 
.A(n_8592),
.B(n_6288),
.Y(n_8725)
);

INVx1_ASAP7_75t_L g8726 ( 
.A(n_8602),
.Y(n_8726)
);

NOR2xp33_ASAP7_75t_L g8727 ( 
.A(n_8601),
.B(n_6288),
.Y(n_8727)
);

OAI22xp5_ASAP7_75t_SL g8728 ( 
.A1(n_8630),
.A2(n_6096),
.B1(n_6071),
.B2(n_6419),
.Y(n_8728)
);

INVx2_ASAP7_75t_SL g8729 ( 
.A(n_8593),
.Y(n_8729)
);

AND2x2_ASAP7_75t_L g8730 ( 
.A(n_8633),
.B(n_6437),
.Y(n_8730)
);

OR2x2_ASAP7_75t_L g8731 ( 
.A(n_8584),
.B(n_6440),
.Y(n_8731)
);

OAI22xp5_ASAP7_75t_SL g8732 ( 
.A1(n_8617),
.A2(n_6419),
.B1(n_5932),
.B2(n_5972),
.Y(n_8732)
);

INVx1_ASAP7_75t_L g8733 ( 
.A(n_8626),
.Y(n_8733)
);

INVx1_ASAP7_75t_L g8734 ( 
.A(n_8632),
.Y(n_8734)
);

INVx1_ASAP7_75t_L g8735 ( 
.A(n_8537),
.Y(n_8735)
);

INVx3_ASAP7_75t_L g8736 ( 
.A(n_8591),
.Y(n_8736)
);

INVx1_ASAP7_75t_L g8737 ( 
.A(n_8598),
.Y(n_8737)
);

INVx1_ASAP7_75t_L g8738 ( 
.A(n_8608),
.Y(n_8738)
);

AOI22xp5_ASAP7_75t_L g8739 ( 
.A1(n_8660),
.A2(n_8590),
.B1(n_8566),
.B2(n_8619),
.Y(n_8739)
);

OAI211xp5_ASAP7_75t_L g8740 ( 
.A1(n_8674),
.A2(n_8629),
.B(n_8618),
.C(n_8599),
.Y(n_8740)
);

AOI322xp5_ASAP7_75t_L g8741 ( 
.A1(n_8692),
.A2(n_8610),
.A3(n_8577),
.B1(n_8583),
.B2(n_8627),
.C1(n_8605),
.C2(n_8548),
.Y(n_8741)
);

OAI21xp33_ASAP7_75t_L g8742 ( 
.A1(n_8687),
.A2(n_8615),
.B(n_8613),
.Y(n_8742)
);

AOI322xp5_ASAP7_75t_L g8743 ( 
.A1(n_8638),
.A2(n_8639),
.A3(n_8718),
.B1(n_8690),
.B2(n_8737),
.C1(n_8677),
.C2(n_8702),
.Y(n_8743)
);

AOI22xp5_ASAP7_75t_L g8744 ( 
.A1(n_8672),
.A2(n_8589),
.B1(n_6440),
.B2(n_6285),
.Y(n_8744)
);

NAND2xp33_ASAP7_75t_L g8745 ( 
.A(n_8647),
.B(n_6000),
.Y(n_8745)
);

AO22x2_ASAP7_75t_L g8746 ( 
.A1(n_8682),
.A2(n_8547),
.B1(n_8621),
.B2(n_6492),
.Y(n_8746)
);

OAI21xp5_ASAP7_75t_L g8747 ( 
.A1(n_8649),
.A2(n_8642),
.B(n_8688),
.Y(n_8747)
);

NAND2xp5_ASAP7_75t_SL g8748 ( 
.A(n_8649),
.B(n_6084),
.Y(n_8748)
);

AOI22xp5_ASAP7_75t_L g8749 ( 
.A1(n_8701),
.A2(n_6440),
.B1(n_6285),
.B2(n_6278),
.Y(n_8749)
);

OAI22xp5_ASAP7_75t_L g8750 ( 
.A1(n_8670),
.A2(n_6440),
.B1(n_6285),
.B2(n_6278),
.Y(n_8750)
);

OAI322xp33_ASAP7_75t_L g8751 ( 
.A1(n_8636),
.A2(n_5297),
.A3(n_5564),
.B1(n_6312),
.B2(n_4832),
.C1(n_4804),
.C2(n_4809),
.Y(n_8751)
);

OAI21xp5_ASAP7_75t_L g8752 ( 
.A1(n_8688),
.A2(n_6285),
.B(n_6278),
.Y(n_8752)
);

AOI221xp5_ASAP7_75t_L g8753 ( 
.A1(n_8693),
.A2(n_6346),
.B1(n_6317),
.B2(n_6367),
.C(n_6365),
.Y(n_8753)
);

AOI22xp5_ASAP7_75t_L g8754 ( 
.A1(n_8717),
.A2(n_6278),
.B1(n_6492),
.B2(n_6488),
.Y(n_8754)
);

OAI221xp5_ASAP7_75t_SL g8755 ( 
.A1(n_8653),
.A2(n_5972),
.B1(n_5973),
.B2(n_5963),
.C(n_5932),
.Y(n_8755)
);

OAI321xp33_ASAP7_75t_L g8756 ( 
.A1(n_8658),
.A2(n_5963),
.A3(n_5999),
.B1(n_5973),
.B2(n_5874),
.C(n_5909),
.Y(n_8756)
);

AOI22xp33_ASAP7_75t_L g8757 ( 
.A1(n_8707),
.A2(n_6185),
.B1(n_6203),
.B2(n_6488),
.Y(n_8757)
);

INVx2_ASAP7_75t_L g8758 ( 
.A(n_8646),
.Y(n_8758)
);

AOI22xp33_ASAP7_75t_SL g8759 ( 
.A1(n_8637),
.A2(n_6185),
.B1(n_6203),
.B2(n_6337),
.Y(n_8759)
);

OAI22xp5_ASAP7_75t_L g8760 ( 
.A1(n_8680),
.A2(n_6492),
.B1(n_6499),
.B2(n_6488),
.Y(n_8760)
);

INVx1_ASAP7_75t_L g8761 ( 
.A(n_8709),
.Y(n_8761)
);

NAND2xp5_ASAP7_75t_L g8762 ( 
.A(n_8724),
.B(n_6185),
.Y(n_8762)
);

OR2x2_ASAP7_75t_L g8763 ( 
.A(n_8640),
.B(n_6365),
.Y(n_8763)
);

NAND2xp5_ASAP7_75t_SL g8764 ( 
.A(n_8659),
.B(n_6084),
.Y(n_8764)
);

OAI21xp5_ASAP7_75t_SL g8765 ( 
.A1(n_8644),
.A2(n_5506),
.B(n_5521),
.Y(n_8765)
);

OAI22xp33_ASAP7_75t_SL g8766 ( 
.A1(n_8715),
.A2(n_5999),
.B1(n_5874),
.B2(n_5909),
.Y(n_8766)
);

NOR3xp33_ASAP7_75t_L g8767 ( 
.A(n_8634),
.B(n_5464),
.C(n_5460),
.Y(n_8767)
);

OAI22xp5_ASAP7_75t_L g8768 ( 
.A1(n_8691),
.A2(n_6492),
.B1(n_6499),
.B2(n_6488),
.Y(n_8768)
);

INVx1_ASAP7_75t_L g8769 ( 
.A(n_8648),
.Y(n_8769)
);

AOI221xp5_ASAP7_75t_L g8770 ( 
.A1(n_8635),
.A2(n_6346),
.B1(n_6317),
.B2(n_6367),
.C(n_4737),
.Y(n_8770)
);

OAI22xp5_ASAP7_75t_L g8771 ( 
.A1(n_8678),
.A2(n_6499),
.B1(n_6185),
.B2(n_6203),
.Y(n_8771)
);

INVx2_ASAP7_75t_L g8772 ( 
.A(n_8731),
.Y(n_8772)
);

NOR2xp33_ASAP7_75t_L g8773 ( 
.A(n_8652),
.B(n_8641),
.Y(n_8773)
);

AOI22xp5_ASAP7_75t_L g8774 ( 
.A1(n_8696),
.A2(n_6499),
.B1(n_6203),
.B2(n_6337),
.Y(n_8774)
);

INVx1_ASAP7_75t_L g8775 ( 
.A(n_8643),
.Y(n_8775)
);

OAI221xp5_ASAP7_75t_L g8776 ( 
.A1(n_8644),
.A2(n_6337),
.B1(n_6312),
.B2(n_5538),
.C(n_5909),
.Y(n_8776)
);

AOI222xp33_ASAP7_75t_L g8777 ( 
.A1(n_8723),
.A2(n_6312),
.B1(n_6337),
.B2(n_5512),
.C1(n_5477),
.C2(n_5517),
.Y(n_8777)
);

AOI221xp5_ASAP7_75t_L g8778 ( 
.A1(n_8650),
.A2(n_6367),
.B1(n_4737),
.B2(n_4815),
.C(n_4809),
.Y(n_8778)
);

OAI211xp5_ASAP7_75t_L g8779 ( 
.A1(n_8645),
.A2(n_8713),
.B(n_8657),
.C(n_8726),
.Y(n_8779)
);

AOI322xp5_ASAP7_75t_L g8780 ( 
.A1(n_8690),
.A2(n_5408),
.A3(n_4804),
.B1(n_4832),
.B2(n_4809),
.C1(n_4874),
.C2(n_4815),
.Y(n_8780)
);

INVx1_ASAP7_75t_L g8781 ( 
.A(n_8662),
.Y(n_8781)
);

OAI22xp33_ASAP7_75t_L g8782 ( 
.A1(n_8733),
.A2(n_6312),
.B1(n_5874),
.B2(n_5564),
.Y(n_8782)
);

OAI31xp33_ASAP7_75t_L g8783 ( 
.A1(n_8705),
.A2(n_5408),
.A3(n_5565),
.B(n_5291),
.Y(n_8783)
);

O2A1O1Ixp33_ASAP7_75t_L g8784 ( 
.A1(n_8699),
.A2(n_5823),
.B(n_5296),
.C(n_5467),
.Y(n_8784)
);

AOI221xp5_ASAP7_75t_L g8785 ( 
.A1(n_8703),
.A2(n_4737),
.B1(n_4815),
.B2(n_4809),
.C(n_4804),
.Y(n_8785)
);

NAND3xp33_ASAP7_75t_L g8786 ( 
.A(n_8738),
.B(n_8735),
.C(n_8711),
.Y(n_8786)
);

AOI21xp33_ASAP7_75t_L g8787 ( 
.A1(n_8685),
.A2(n_5477),
.B(n_5464),
.Y(n_8787)
);

OA21x2_ASAP7_75t_L g8788 ( 
.A1(n_8665),
.A2(n_5428),
.B(n_5425),
.Y(n_8788)
);

AOI22xp33_ASAP7_75t_SL g8789 ( 
.A1(n_8734),
.A2(n_6000),
.B1(n_4737),
.B2(n_4809),
.Y(n_8789)
);

INVx1_ASAP7_75t_L g8790 ( 
.A(n_8730),
.Y(n_8790)
);

INVx2_ASAP7_75t_L g8791 ( 
.A(n_8695),
.Y(n_8791)
);

A2O1A1Ixp33_ASAP7_75t_L g8792 ( 
.A1(n_8706),
.A2(n_5512),
.B(n_5517),
.C(n_5496),
.Y(n_8792)
);

OAI21xp33_ASAP7_75t_L g8793 ( 
.A1(n_8686),
.A2(n_5029),
.B(n_5375),
.Y(n_8793)
);

NAND3xp33_ASAP7_75t_L g8794 ( 
.A(n_8694),
.B(n_5620),
.C(n_5519),
.Y(n_8794)
);

OAI221xp5_ASAP7_75t_L g8795 ( 
.A1(n_8656),
.A2(n_5378),
.B1(n_5175),
.B2(n_5482),
.C(n_5480),
.Y(n_8795)
);

INVx1_ASAP7_75t_L g8796 ( 
.A(n_8695),
.Y(n_8796)
);

OAI221xp5_ASAP7_75t_SL g8797 ( 
.A1(n_8679),
.A2(n_5593),
.B1(n_5449),
.B2(n_5397),
.C(n_5396),
.Y(n_8797)
);

OAI221xp5_ASAP7_75t_L g8798 ( 
.A1(n_8675),
.A2(n_5378),
.B1(n_5558),
.B2(n_5461),
.C(n_5422),
.Y(n_8798)
);

NOR2xp33_ASAP7_75t_L g8799 ( 
.A(n_8663),
.B(n_5574),
.Y(n_8799)
);

AND2x2_ASAP7_75t_L g8800 ( 
.A(n_8722),
.B(n_5565),
.Y(n_8800)
);

OAI21xp5_ASAP7_75t_L g8801 ( 
.A1(n_8654),
.A2(n_5519),
.B(n_5496),
.Y(n_8801)
);

OAI21x1_ASAP7_75t_L g8802 ( 
.A1(n_8668),
.A2(n_5557),
.B(n_5281),
.Y(n_8802)
);

AND2x2_ASAP7_75t_L g8803 ( 
.A(n_8698),
.B(n_8669),
.Y(n_8803)
);

OAI31xp33_ASAP7_75t_L g8804 ( 
.A1(n_8683),
.A2(n_5547),
.A3(n_5559),
.B(n_5543),
.Y(n_8804)
);

OAI21xp5_ASAP7_75t_L g8805 ( 
.A1(n_8671),
.A2(n_5547),
.B(n_5543),
.Y(n_8805)
);

AOI221xp5_ASAP7_75t_L g8806 ( 
.A1(n_8664),
.A2(n_4737),
.B1(n_4832),
.B2(n_4815),
.C(n_4804),
.Y(n_8806)
);

AOI21xp33_ASAP7_75t_L g8807 ( 
.A1(n_8725),
.A2(n_5580),
.B(n_5559),
.Y(n_8807)
);

OA33x2_ASAP7_75t_L g8808 ( 
.A1(n_8700),
.A2(n_5073),
.A3(n_5004),
.B1(n_5032),
.B2(n_5020),
.B3(n_5578),
.Y(n_8808)
);

NAND2xp5_ASAP7_75t_L g8809 ( 
.A(n_8697),
.B(n_6459),
.Y(n_8809)
);

INVx1_ASAP7_75t_L g8810 ( 
.A(n_8673),
.Y(n_8810)
);

AOI22xp5_ASAP7_75t_L g8811 ( 
.A1(n_8710),
.A2(n_5580),
.B1(n_5610),
.B2(n_5608),
.Y(n_8811)
);

AOI22xp33_ASAP7_75t_L g8812 ( 
.A1(n_8728),
.A2(n_5620),
.B1(n_4815),
.B2(n_4832),
.Y(n_8812)
);

AOI21xp5_ASAP7_75t_L g8813 ( 
.A1(n_8720),
.A2(n_8729),
.B(n_8704),
.Y(n_8813)
);

AOI32xp33_ASAP7_75t_L g8814 ( 
.A1(n_8736),
.A2(n_4659),
.A3(n_4588),
.B1(n_5591),
.B2(n_4832),
.Y(n_8814)
);

OAI21xp5_ASAP7_75t_L g8815 ( 
.A1(n_8712),
.A2(n_5610),
.B(n_5608),
.Y(n_8815)
);

INVx1_ASAP7_75t_L g8816 ( 
.A(n_8684),
.Y(n_8816)
);

AOI22xp5_ASAP7_75t_L g8817 ( 
.A1(n_8736),
.A2(n_5623),
.B1(n_5625),
.B2(n_5378),
.Y(n_8817)
);

INVx1_ASAP7_75t_L g8818 ( 
.A(n_8661),
.Y(n_8818)
);

O2A1O1Ixp5_ASAP7_75t_SL g8819 ( 
.A1(n_8689),
.A2(n_5428),
.B(n_5430),
.C(n_5425),
.Y(n_8819)
);

OAI21xp33_ASAP7_75t_L g8820 ( 
.A1(n_8708),
.A2(n_5433),
.B(n_5430),
.Y(n_8820)
);

NAND2xp5_ASAP7_75t_L g8821 ( 
.A(n_8676),
.B(n_6459),
.Y(n_8821)
);

INVx1_ASAP7_75t_L g8822 ( 
.A(n_8667),
.Y(n_8822)
);

AOI21xp5_ASAP7_75t_L g8823 ( 
.A1(n_8727),
.A2(n_8681),
.B(n_8655),
.Y(n_8823)
);

NOR2xp33_ASAP7_75t_L g8824 ( 
.A(n_8651),
.B(n_5623),
.Y(n_8824)
);

NOR3xp33_ASAP7_75t_SL g8825 ( 
.A(n_8716),
.B(n_5507),
.C(n_5486),
.Y(n_8825)
);

INVx1_ASAP7_75t_L g8826 ( 
.A(n_8714),
.Y(n_8826)
);

NAND2xp5_ASAP7_75t_L g8827 ( 
.A(n_8666),
.B(n_6459),
.Y(n_8827)
);

INVx1_ASAP7_75t_L g8828 ( 
.A(n_8732),
.Y(n_8828)
);

OAI222xp33_ASAP7_75t_L g8829 ( 
.A1(n_8719),
.A2(n_8721),
.B1(n_5593),
.B2(n_5558),
.C1(n_4874),
.C2(n_4804),
.Y(n_8829)
);

NAND2xp5_ASAP7_75t_L g8830 ( 
.A(n_8677),
.B(n_6459),
.Y(n_8830)
);

NAND2xp5_ASAP7_75t_L g8831 ( 
.A(n_8677),
.B(n_6459),
.Y(n_8831)
);

AOI311xp33_ASAP7_75t_L g8832 ( 
.A1(n_8674),
.A2(n_5448),
.A3(n_5450),
.B(n_5445),
.C(n_5433),
.Y(n_8832)
);

NAND2xp5_ASAP7_75t_L g8833 ( 
.A(n_8747),
.B(n_5708),
.Y(n_8833)
);

INVx1_ASAP7_75t_L g8834 ( 
.A(n_8746),
.Y(n_8834)
);

NOR2x1_ASAP7_75t_L g8835 ( 
.A(n_8786),
.B(n_8779),
.Y(n_8835)
);

OAI211xp5_ASAP7_75t_L g8836 ( 
.A1(n_8743),
.A2(n_5510),
.B(n_5271),
.C(n_5479),
.Y(n_8836)
);

AOI22xp5_ASAP7_75t_L g8837 ( 
.A1(n_8761),
.A2(n_5625),
.B1(n_5620),
.B2(n_4588),
.Y(n_8837)
);

INVx1_ASAP7_75t_L g8838 ( 
.A(n_8746),
.Y(n_8838)
);

NAND2xp5_ASAP7_75t_L g8839 ( 
.A(n_8752),
.B(n_5708),
.Y(n_8839)
);

INVx2_ASAP7_75t_L g8840 ( 
.A(n_8758),
.Y(n_8840)
);

INVx2_ASAP7_75t_L g8841 ( 
.A(n_8775),
.Y(n_8841)
);

NOR3xp33_ASAP7_75t_L g8842 ( 
.A(n_8740),
.B(n_5594),
.C(n_5002),
.Y(n_8842)
);

INVx1_ASAP7_75t_L g8843 ( 
.A(n_8773),
.Y(n_8843)
);

NOR2x1_ASAP7_75t_L g8844 ( 
.A(n_8769),
.B(n_5445),
.Y(n_8844)
);

INVx1_ASAP7_75t_L g8845 ( 
.A(n_8830),
.Y(n_8845)
);

AOI221xp5_ASAP7_75t_SL g8846 ( 
.A1(n_8745),
.A2(n_5448),
.B1(n_5456),
.B2(n_5455),
.C(n_5450),
.Y(n_8846)
);

INVx1_ASAP7_75t_L g8847 ( 
.A(n_8831),
.Y(n_8847)
);

AND2x2_ASAP7_75t_L g8848 ( 
.A(n_8781),
.B(n_8825),
.Y(n_8848)
);

AO21x1_ASAP7_75t_L g8849 ( 
.A1(n_8816),
.A2(n_5456),
.B(n_5455),
.Y(n_8849)
);

AOI221xp5_ASAP7_75t_L g8850 ( 
.A1(n_8822),
.A2(n_4874),
.B1(n_5002),
.B2(n_5003),
.C(n_4913),
.Y(n_8850)
);

INVx1_ASAP7_75t_L g8851 ( 
.A(n_8762),
.Y(n_8851)
);

OAI32xp33_ASAP7_75t_L g8852 ( 
.A1(n_8790),
.A2(n_5558),
.A3(n_4659),
.B1(n_4588),
.B2(n_5466),
.Y(n_8852)
);

INVx1_ASAP7_75t_L g8853 ( 
.A(n_8791),
.Y(n_8853)
);

OAI22xp33_ASAP7_75t_L g8854 ( 
.A1(n_8739),
.A2(n_8772),
.B1(n_8744),
.B2(n_8763),
.Y(n_8854)
);

OAI322xp33_ASAP7_75t_L g8855 ( 
.A1(n_8813),
.A2(n_4874),
.A3(n_5470),
.B1(n_5550),
.B2(n_5605),
.C1(n_5466),
.C2(n_5457),
.Y(n_8855)
);

OAI211xp5_ASAP7_75t_SL g8856 ( 
.A1(n_8742),
.A2(n_5474),
.B(n_5328),
.C(n_4588),
.Y(n_8856)
);

INVx2_ASAP7_75t_L g8857 ( 
.A(n_8788),
.Y(n_8857)
);

INVx1_ASAP7_75t_L g8858 ( 
.A(n_8796),
.Y(n_8858)
);

OAI221xp5_ASAP7_75t_L g8859 ( 
.A1(n_8748),
.A2(n_5552),
.B1(n_5534),
.B2(n_4659),
.C(n_5255),
.Y(n_8859)
);

INVx1_ASAP7_75t_L g8860 ( 
.A(n_8809),
.Y(n_8860)
);

OAI211xp5_ASAP7_75t_L g8861 ( 
.A1(n_8741),
.A2(n_4659),
.B(n_5583),
.C(n_5354),
.Y(n_8861)
);

OAI211xp5_ASAP7_75t_L g8862 ( 
.A1(n_8823),
.A2(n_5256),
.B(n_5470),
.C(n_5457),
.Y(n_8862)
);

O2A1O1Ixp33_ASAP7_75t_L g8863 ( 
.A1(n_8826),
.A2(n_8828),
.B(n_8810),
.C(n_8818),
.Y(n_8863)
);

AOI211xp5_ASAP7_75t_SL g8864 ( 
.A1(n_8803),
.A2(n_5581),
.B(n_5567),
.C(n_5589),
.Y(n_8864)
);

AOI22xp33_ASAP7_75t_L g8865 ( 
.A1(n_8759),
.A2(n_4874),
.B1(n_4792),
.B2(n_4799),
.Y(n_8865)
);

AOI221xp5_ASAP7_75t_L g8866 ( 
.A1(n_8753),
.A2(n_5003),
.B1(n_5036),
.B2(n_5002),
.C(n_4913),
.Y(n_8866)
);

AOI22xp5_ASAP7_75t_L g8867 ( 
.A1(n_8749),
.A2(n_5605),
.B1(n_5550),
.B2(n_5552),
.Y(n_8867)
);

AOI221xp5_ASAP7_75t_L g8868 ( 
.A1(n_8827),
.A2(n_8764),
.B1(n_8821),
.B2(n_8750),
.C(n_8824),
.Y(n_8868)
);

INVx1_ASAP7_75t_L g8869 ( 
.A(n_8788),
.Y(n_8869)
);

INVx1_ASAP7_75t_L g8870 ( 
.A(n_8767),
.Y(n_8870)
);

AOI21xp33_ASAP7_75t_L g8871 ( 
.A1(n_8777),
.A2(n_4792),
.B(n_4742),
.Y(n_8871)
);

AND2x2_ASAP7_75t_L g8872 ( 
.A(n_8800),
.B(n_5708),
.Y(n_8872)
);

AOI332xp33_ASAP7_75t_L g8873 ( 
.A1(n_8812),
.A2(n_5497),
.A3(n_5503),
.B1(n_5513),
.B2(n_5514),
.B3(n_5626),
.C1(n_5622),
.C2(n_5598),
.Y(n_8873)
);

AOI22xp33_ASAP7_75t_L g8874 ( 
.A1(n_8771),
.A2(n_4792),
.B1(n_4799),
.B2(n_4742),
.Y(n_8874)
);

NAND2xp5_ASAP7_75t_L g8875 ( 
.A(n_8799),
.B(n_5734),
.Y(n_8875)
);

NAND4xp75_ASAP7_75t_L g8876 ( 
.A(n_8804),
.B(n_8770),
.C(n_8787),
.D(n_8815),
.Y(n_8876)
);

OAI21xp33_ASAP7_75t_L g8877 ( 
.A1(n_8793),
.A2(n_5537),
.B(n_5522),
.Y(n_8877)
);

AOI22xp5_ASAP7_75t_L g8878 ( 
.A1(n_8765),
.A2(n_5552),
.B1(n_5586),
.B2(n_5555),
.Y(n_8878)
);

OAI31xp33_ASAP7_75t_L g8879 ( 
.A1(n_8829),
.A2(n_4580),
.A3(n_5002),
.B(n_4913),
.Y(n_8879)
);

OAI222xp33_ASAP7_75t_L g8880 ( 
.A1(n_8755),
.A2(n_5593),
.B1(n_5525),
.B2(n_4580),
.C1(n_5002),
.C2(n_5036),
.Y(n_8880)
);

AOI221xp5_ASAP7_75t_L g8881 ( 
.A1(n_8794),
.A2(n_5036),
.B1(n_5003),
.B2(n_4913),
.C(n_4799),
.Y(n_8881)
);

NAND2xp5_ASAP7_75t_L g8882 ( 
.A(n_8757),
.B(n_8754),
.Y(n_8882)
);

OAI211xp5_ASAP7_75t_L g8883 ( 
.A1(n_8832),
.A2(n_8820),
.B(n_8789),
.C(n_8783),
.Y(n_8883)
);

NOR2xp33_ASAP7_75t_SL g8884 ( 
.A(n_8784),
.B(n_5070),
.Y(n_8884)
);

NAND3xp33_ASAP7_75t_L g8885 ( 
.A(n_8774),
.B(n_5473),
.C(n_5444),
.Y(n_8885)
);

AOI221x1_ASAP7_75t_L g8886 ( 
.A1(n_8807),
.A2(n_5595),
.B1(n_4718),
.B2(n_4725),
.C(n_4722),
.Y(n_8886)
);

AND2x2_ASAP7_75t_L g8887 ( 
.A(n_8802),
.B(n_8819),
.Y(n_8887)
);

AOI22xp33_ASAP7_75t_L g8888 ( 
.A1(n_8768),
.A2(n_4792),
.B1(n_4799),
.B2(n_4742),
.Y(n_8888)
);

AOI221xp5_ASAP7_75t_L g8889 ( 
.A1(n_8805),
.A2(n_8760),
.B1(n_8776),
.B2(n_8778),
.C(n_8801),
.Y(n_8889)
);

AOI22xp33_ASAP7_75t_L g8890 ( 
.A1(n_8785),
.A2(n_4824),
.B1(n_4843),
.B2(n_4742),
.Y(n_8890)
);

AOI211x1_ASAP7_75t_SL g8891 ( 
.A1(n_8792),
.A2(n_5734),
.B(n_5774),
.C(n_5741),
.Y(n_8891)
);

AOI22xp5_ASAP7_75t_L g8892 ( 
.A1(n_8795),
.A2(n_8817),
.B1(n_8782),
.B2(n_8798),
.Y(n_8892)
);

OAI221xp5_ASAP7_75t_L g8893 ( 
.A1(n_8814),
.A2(n_5198),
.B1(n_5528),
.B2(n_4977),
.C(n_5195),
.Y(n_8893)
);

OAI21xp33_ASAP7_75t_L g8894 ( 
.A1(n_8780),
.A2(n_8766),
.B(n_8797),
.Y(n_8894)
);

AOI221xp5_ASAP7_75t_L g8895 ( 
.A1(n_8751),
.A2(n_5036),
.B1(n_5003),
.B2(n_4913),
.C(n_4845),
.Y(n_8895)
);

OAI211xp5_ASAP7_75t_L g8896 ( 
.A1(n_8806),
.A2(n_4863),
.B(n_4762),
.C(n_4836),
.Y(n_8896)
);

NAND2xp5_ASAP7_75t_L g8897 ( 
.A(n_8811),
.B(n_5734),
.Y(n_8897)
);

NAND3xp33_ASAP7_75t_L g8898 ( 
.A(n_8756),
.B(n_5473),
.C(n_5444),
.Y(n_8898)
);

INVx2_ASAP7_75t_SL g8899 ( 
.A(n_8808),
.Y(n_8899)
);

OAI21xp5_ASAP7_75t_L g8900 ( 
.A1(n_8747),
.A2(n_4843),
.B(n_4824),
.Y(n_8900)
);

AOI222xp33_ASAP7_75t_L g8901 ( 
.A1(n_8752),
.A2(n_5036),
.B1(n_5003),
.B2(n_4843),
.C1(n_4824),
.C2(n_4859),
.Y(n_8901)
);

OAI21xp33_ASAP7_75t_SL g8902 ( 
.A1(n_8819),
.A2(n_4958),
.B(n_4878),
.Y(n_8902)
);

AOI32xp33_ASAP7_75t_L g8903 ( 
.A1(n_8761),
.A2(n_4580),
.A3(n_4646),
.B1(n_4884),
.B2(n_4827),
.Y(n_8903)
);

NAND2xp5_ASAP7_75t_L g8904 ( 
.A(n_8747),
.B(n_5734),
.Y(n_8904)
);

OAI21xp33_ASAP7_75t_SL g8905 ( 
.A1(n_8819),
.A2(n_4958),
.B(n_4878),
.Y(n_8905)
);

OAI21xp5_ASAP7_75t_L g8906 ( 
.A1(n_8747),
.A2(n_4843),
.B(n_4824),
.Y(n_8906)
);

AOI22xp33_ASAP7_75t_L g8907 ( 
.A1(n_8790),
.A2(n_4850),
.B1(n_4859),
.B2(n_4845),
.Y(n_8907)
);

O2A1O1Ixp5_ASAP7_75t_L g8908 ( 
.A1(n_8748),
.A2(n_4706),
.B(n_4725),
.C(n_4722),
.Y(n_8908)
);

AOI311xp33_ASAP7_75t_L g8909 ( 
.A1(n_8779),
.A2(n_4722),
.A3(n_4764),
.B(n_4725),
.C(n_4706),
.Y(n_8909)
);

OAI22xp5_ASAP7_75t_L g8910 ( 
.A1(n_8786),
.A2(n_5072),
.B1(n_5152),
.B2(n_4850),
.Y(n_8910)
);

OAI22xp5_ASAP7_75t_L g8911 ( 
.A1(n_8786),
.A2(n_5072),
.B1(n_4850),
.B2(n_4859),
.Y(n_8911)
);

AOI22xp33_ASAP7_75t_L g8912 ( 
.A1(n_8790),
.A2(n_4850),
.B1(n_4859),
.B2(n_4845),
.Y(n_8912)
);

AOI222xp33_ASAP7_75t_L g8913 ( 
.A1(n_8752),
.A2(n_4845),
.B1(n_4866),
.B2(n_5741),
.C1(n_5774),
.C2(n_5959),
.Y(n_8913)
);

AOI221x1_ASAP7_75t_L g8914 ( 
.A1(n_8747),
.A2(n_4764),
.B1(n_4776),
.B2(n_4770),
.C(n_4768),
.Y(n_8914)
);

AND2x2_ASAP7_75t_SL g8915 ( 
.A(n_8773),
.B(n_4762),
.Y(n_8915)
);

INVx1_ASAP7_75t_L g8916 ( 
.A(n_8746),
.Y(n_8916)
);

O2A1O1Ixp33_ASAP7_75t_SL g8917 ( 
.A1(n_8779),
.A2(n_4958),
.B(n_5060),
.C(n_4878),
.Y(n_8917)
);

OAI221xp5_ASAP7_75t_L g8918 ( 
.A1(n_8747),
.A2(n_5528),
.B1(n_4977),
.B2(n_5473),
.C(n_5444),
.Y(n_8918)
);

NAND2xp5_ASAP7_75t_L g8919 ( 
.A(n_8747),
.B(n_5741),
.Y(n_8919)
);

OAI22xp5_ASAP7_75t_L g8920 ( 
.A1(n_8786),
.A2(n_5072),
.B1(n_4866),
.B2(n_4981),
.Y(n_8920)
);

INVx1_ASAP7_75t_L g8921 ( 
.A(n_8746),
.Y(n_8921)
);

NAND2xp5_ASAP7_75t_SL g8922 ( 
.A(n_8747),
.B(n_4820),
.Y(n_8922)
);

AOI21xp5_ASAP7_75t_L g8923 ( 
.A1(n_8748),
.A2(n_5528),
.B(n_4837),
.Y(n_8923)
);

INVx1_ASAP7_75t_L g8924 ( 
.A(n_8835),
.Y(n_8924)
);

INVx5_ASAP7_75t_L g8925 ( 
.A(n_8841),
.Y(n_8925)
);

NAND2xp5_ASAP7_75t_L g8926 ( 
.A(n_8899),
.B(n_8915),
.Y(n_8926)
);

NAND2xp5_ASAP7_75t_L g8927 ( 
.A(n_8840),
.B(n_5741),
.Y(n_8927)
);

OAI22xp5_ASAP7_75t_L g8928 ( 
.A1(n_8892),
.A2(n_5072),
.B1(n_4866),
.B2(n_4977),
.Y(n_8928)
);

INVx1_ASAP7_75t_L g8929 ( 
.A(n_8834),
.Y(n_8929)
);

NAND2x1_ASAP7_75t_L g8930 ( 
.A(n_8843),
.B(n_4708),
.Y(n_8930)
);

AND2x2_ASAP7_75t_L g8931 ( 
.A(n_8848),
.B(n_5774),
.Y(n_8931)
);

NAND2xp5_ASAP7_75t_L g8932 ( 
.A(n_8851),
.B(n_5774),
.Y(n_8932)
);

NAND2xp5_ASAP7_75t_L g8933 ( 
.A(n_8854),
.B(n_5959),
.Y(n_8933)
);

INVx1_ASAP7_75t_L g8934 ( 
.A(n_8838),
.Y(n_8934)
);

AND2x2_ASAP7_75t_L g8935 ( 
.A(n_8884),
.B(n_5959),
.Y(n_8935)
);

AND2x2_ASAP7_75t_L g8936 ( 
.A(n_8858),
.B(n_5959),
.Y(n_8936)
);

INVx1_ASAP7_75t_L g8937 ( 
.A(n_8916),
.Y(n_8937)
);

INVx1_ASAP7_75t_L g8938 ( 
.A(n_8921),
.Y(n_8938)
);

INVx1_ASAP7_75t_SL g8939 ( 
.A(n_8853),
.Y(n_8939)
);

NAND2xp33_ASAP7_75t_L g8940 ( 
.A(n_8894),
.B(n_5072),
.Y(n_8940)
);

INVx1_ASAP7_75t_L g8941 ( 
.A(n_8887),
.Y(n_8941)
);

OAI32xp33_ASAP7_75t_L g8942 ( 
.A1(n_8882),
.A2(n_4977),
.A3(n_4848),
.B1(n_4872),
.B2(n_4807),
.Y(n_8942)
);

INVx3_ASAP7_75t_L g8943 ( 
.A(n_8857),
.Y(n_8943)
);

NAND4xp25_ASAP7_75t_L g8944 ( 
.A(n_8863),
.B(n_8868),
.C(n_8870),
.D(n_8869),
.Y(n_8944)
);

NAND2xp5_ASAP7_75t_L g8945 ( 
.A(n_8872),
.B(n_5906),
.Y(n_8945)
);

INVx1_ASAP7_75t_L g8946 ( 
.A(n_8849),
.Y(n_8946)
);

INVx1_ASAP7_75t_L g8947 ( 
.A(n_8833),
.Y(n_8947)
);

NAND2xp5_ASAP7_75t_L g8948 ( 
.A(n_8904),
.B(n_5906),
.Y(n_8948)
);

AND2x2_ASAP7_75t_L g8949 ( 
.A(n_8922),
.B(n_4825),
.Y(n_8949)
);

NOR2xp33_ASAP7_75t_L g8950 ( 
.A(n_8919),
.B(n_4866),
.Y(n_8950)
);

NAND2xp5_ASAP7_75t_L g8951 ( 
.A(n_8860),
.B(n_5906),
.Y(n_8951)
);

OR2x2_ASAP7_75t_L g8952 ( 
.A(n_8839),
.B(n_5906),
.Y(n_8952)
);

NOR3xp33_ASAP7_75t_L g8953 ( 
.A(n_8845),
.B(n_5525),
.C(n_5624),
.Y(n_8953)
);

INVx1_ASAP7_75t_L g8954 ( 
.A(n_8844),
.Y(n_8954)
);

AND2x2_ASAP7_75t_L g8955 ( 
.A(n_8842),
.B(n_4825),
.Y(n_8955)
);

OAI22xp5_ASAP7_75t_L g8956 ( 
.A1(n_8878),
.A2(n_5072),
.B1(n_4984),
.B2(n_4981),
.Y(n_8956)
);

NAND2xp5_ASAP7_75t_SL g8957 ( 
.A(n_8889),
.B(n_5072),
.Y(n_8957)
);

AND2x2_ASAP7_75t_L g8958 ( 
.A(n_8909),
.B(n_4853),
.Y(n_8958)
);

INVx1_ASAP7_75t_L g8959 ( 
.A(n_8875),
.Y(n_8959)
);

INVx1_ASAP7_75t_L g8960 ( 
.A(n_8897),
.Y(n_8960)
);

INVx1_ASAP7_75t_SL g8961 ( 
.A(n_8876),
.Y(n_8961)
);

AND2x4_ASAP7_75t_L g8962 ( 
.A(n_8847),
.B(n_5930),
.Y(n_8962)
);

INVx1_ASAP7_75t_L g8963 ( 
.A(n_8883),
.Y(n_8963)
);

NAND4xp25_ASAP7_75t_L g8964 ( 
.A(n_8837),
.B(n_4884),
.C(n_4932),
.D(n_4827),
.Y(n_8964)
);

NAND2xp5_ASAP7_75t_SL g8965 ( 
.A(n_8900),
.B(n_5072),
.Y(n_8965)
);

HB1xp67_ASAP7_75t_L g8966 ( 
.A(n_8906),
.Y(n_8966)
);

NAND2xp5_ASAP7_75t_L g8967 ( 
.A(n_8846),
.B(n_5930),
.Y(n_8967)
);

AND2x2_ASAP7_75t_L g8968 ( 
.A(n_8836),
.B(n_4853),
.Y(n_8968)
);

NOR3xp33_ASAP7_75t_L g8969 ( 
.A(n_8920),
.B(n_5624),
.C(n_5404),
.Y(n_8969)
);

NAND2xp33_ASAP7_75t_L g8970 ( 
.A(n_8903),
.B(n_4820),
.Y(n_8970)
);

HB1xp67_ASAP7_75t_L g8971 ( 
.A(n_8902),
.Y(n_8971)
);

INVx2_ASAP7_75t_SL g8972 ( 
.A(n_8911),
.Y(n_8972)
);

NAND2xp33_ASAP7_75t_L g8973 ( 
.A(n_8877),
.B(n_4820),
.Y(n_8973)
);

OR2x2_ASAP7_75t_L g8974 ( 
.A(n_8910),
.B(n_5930),
.Y(n_8974)
);

NAND2xp5_ASAP7_75t_SL g8975 ( 
.A(n_8879),
.B(n_4820),
.Y(n_8975)
);

NAND2xp5_ASAP7_75t_L g8976 ( 
.A(n_8867),
.B(n_5930),
.Y(n_8976)
);

INVx1_ASAP7_75t_L g8977 ( 
.A(n_8862),
.Y(n_8977)
);

INVx1_ASAP7_75t_L g8978 ( 
.A(n_8914),
.Y(n_8978)
);

AND2x2_ASAP7_75t_L g8979 ( 
.A(n_8864),
.B(n_4853),
.Y(n_8979)
);

INVx1_ASAP7_75t_L g8980 ( 
.A(n_8908),
.Y(n_8980)
);

AOI21xp5_ASAP7_75t_L g8981 ( 
.A1(n_8861),
.A2(n_4837),
.B(n_4835),
.Y(n_8981)
);

NAND2xp5_ASAP7_75t_SL g8982 ( 
.A(n_8905),
.B(n_8850),
.Y(n_8982)
);

INVx1_ASAP7_75t_L g8983 ( 
.A(n_8917),
.Y(n_8983)
);

NOR2xp33_ASAP7_75t_L g8984 ( 
.A(n_8880),
.B(n_4915),
.Y(n_8984)
);

NOR2xp33_ASAP7_75t_L g8985 ( 
.A(n_8855),
.B(n_4915),
.Y(n_8985)
);

INVx1_ASAP7_75t_L g8986 ( 
.A(n_8886),
.Y(n_8986)
);

NOR2xp33_ASAP7_75t_L g8987 ( 
.A(n_8855),
.B(n_4915),
.Y(n_8987)
);

AND2x2_ASAP7_75t_L g8988 ( 
.A(n_8888),
.B(n_4853),
.Y(n_8988)
);

AND2x2_ASAP7_75t_L g8989 ( 
.A(n_8874),
.B(n_8865),
.Y(n_8989)
);

NAND2xp5_ASAP7_75t_L g8990 ( 
.A(n_8891),
.B(n_5935),
.Y(n_8990)
);

AND2x2_ASAP7_75t_L g8991 ( 
.A(n_8890),
.B(n_4853),
.Y(n_8991)
);

INVx1_ASAP7_75t_L g8992 ( 
.A(n_8891),
.Y(n_8992)
);

INVx1_ASAP7_75t_L g8993 ( 
.A(n_8898),
.Y(n_8993)
);

AOI322xp5_ASAP7_75t_L g8994 ( 
.A1(n_8961),
.A2(n_8871),
.A3(n_8907),
.B1(n_8912),
.B2(n_8866),
.C1(n_8895),
.C2(n_8881),
.Y(n_8994)
);

OAI211xp5_ASAP7_75t_SL g8995 ( 
.A1(n_8941),
.A2(n_8896),
.B(n_8913),
.C(n_8893),
.Y(n_8995)
);

NAND4xp25_ASAP7_75t_L g8996 ( 
.A(n_8924),
.B(n_8856),
.C(n_8859),
.D(n_8885),
.Y(n_8996)
);

AOI211xp5_ASAP7_75t_L g8997 ( 
.A1(n_8944),
.A2(n_8852),
.B(n_8918),
.C(n_8885),
.Y(n_8997)
);

NAND5xp2_ASAP7_75t_L g8998 ( 
.A(n_8963),
.B(n_8873),
.C(n_8923),
.D(n_8901),
.E(n_4848),
.Y(n_8998)
);

NOR3xp33_ASAP7_75t_L g8999 ( 
.A(n_8944),
.B(n_4948),
.C(n_4646),
.Y(n_8999)
);

A2O1A1Ixp33_ASAP7_75t_SL g9000 ( 
.A1(n_8943),
.A2(n_4764),
.B(n_4770),
.C(n_4768),
.Y(n_9000)
);

OA211x2_ASAP7_75t_L g9001 ( 
.A1(n_8926),
.A2(n_4984),
.B(n_5020),
.C(n_5004),
.Y(n_9001)
);

INVx1_ASAP7_75t_SL g9002 ( 
.A(n_8939),
.Y(n_9002)
);

NAND3xp33_ASAP7_75t_L g9003 ( 
.A(n_8925),
.B(n_4992),
.C(n_5032),
.Y(n_9003)
);

XNOR2x1_ASAP7_75t_L g9004 ( 
.A(n_8929),
.B(n_4677),
.Y(n_9004)
);

AOI211xp5_ASAP7_75t_L g9005 ( 
.A1(n_8971),
.A2(n_4836),
.B(n_4858),
.C(n_4820),
.Y(n_9005)
);

AOI21xp33_ASAP7_75t_SL g9006 ( 
.A1(n_8993),
.A2(n_4807),
.B(n_4788),
.Y(n_9006)
);

BUFx2_ASAP7_75t_L g9007 ( 
.A(n_8925),
.Y(n_9007)
);

OAI21xp5_ASAP7_75t_L g9008 ( 
.A1(n_8934),
.A2(n_5073),
.B(n_5386),
.Y(n_9008)
);

HB1xp67_ASAP7_75t_L g9009 ( 
.A(n_8925),
.Y(n_9009)
);

AOI22xp33_ASAP7_75t_L g9010 ( 
.A1(n_8937),
.A2(n_4915),
.B1(n_4701),
.B2(n_4884),
.Y(n_9010)
);

O2A1O1Ixp33_ASAP7_75t_SL g9011 ( 
.A1(n_8983),
.A2(n_5079),
.B(n_5060),
.C(n_4768),
.Y(n_9011)
);

NAND2xp5_ASAP7_75t_L g9012 ( 
.A(n_8943),
.B(n_5935),
.Y(n_9012)
);

AOI221xp5_ASAP7_75t_L g9013 ( 
.A1(n_8938),
.A2(n_8954),
.B1(n_8940),
.B2(n_8992),
.C(n_8986),
.Y(n_9013)
);

AOI221xp5_ASAP7_75t_L g9014 ( 
.A1(n_8946),
.A2(n_4992),
.B1(n_4770),
.B2(n_4781),
.C(n_4778),
.Y(n_9014)
);

INVx2_ASAP7_75t_SL g9015 ( 
.A(n_8966),
.Y(n_9015)
);

AOI221xp5_ASAP7_75t_L g9016 ( 
.A1(n_8980),
.A2(n_4776),
.B1(n_4782),
.B2(n_4781),
.C(n_4778),
.Y(n_9016)
);

NOR3xp33_ASAP7_75t_L g9017 ( 
.A(n_8947),
.B(n_4948),
.C(n_4646),
.Y(n_9017)
);

OAI221xp5_ASAP7_75t_L g9018 ( 
.A1(n_8978),
.A2(n_8977),
.B1(n_8970),
.B2(n_8957),
.C(n_8972),
.Y(n_9018)
);

NAND2xp5_ASAP7_75t_L g9019 ( 
.A(n_8931),
.B(n_5935),
.Y(n_9019)
);

HB1xp67_ASAP7_75t_L g9020 ( 
.A(n_8936),
.Y(n_9020)
);

OAI21xp33_ASAP7_75t_SL g9021 ( 
.A1(n_8965),
.A2(n_5079),
.B(n_5060),
.Y(n_9021)
);

AND2x2_ASAP7_75t_L g9022 ( 
.A(n_8949),
.B(n_5935),
.Y(n_9022)
);

OAI222xp33_ASAP7_75t_L g9023 ( 
.A1(n_8982),
.A2(n_4677),
.B1(n_4988),
.B2(n_4731),
.C1(n_4807),
.C2(n_4848),
.Y(n_9023)
);

AOI211xp5_ASAP7_75t_L g9024 ( 
.A1(n_8959),
.A2(n_8960),
.B(n_8989),
.C(n_8933),
.Y(n_9024)
);

O2A1O1Ixp33_ASAP7_75t_L g9025 ( 
.A1(n_8932),
.A2(n_4788),
.B(n_4848),
.C(n_4807),
.Y(n_9025)
);

AOI211x1_ASAP7_75t_SL g9026 ( 
.A1(n_8927),
.A2(n_4863),
.B(n_5600),
.C(n_5599),
.Y(n_9026)
);

AOI21xp33_ASAP7_75t_SL g9027 ( 
.A1(n_8951),
.A2(n_4872),
.B(n_4788),
.Y(n_9027)
);

AOI22xp5_ASAP7_75t_L g9028 ( 
.A1(n_8968),
.A2(n_4837),
.B1(n_4835),
.B2(n_4836),
.Y(n_9028)
);

AOI22xp5_ASAP7_75t_L g9029 ( 
.A1(n_8985),
.A2(n_4837),
.B1(n_4835),
.B2(n_4836),
.Y(n_9029)
);

AOI221xp5_ASAP7_75t_L g9030 ( 
.A1(n_8950),
.A2(n_4776),
.B1(n_4782),
.B2(n_4781),
.C(n_4778),
.Y(n_9030)
);

NAND4xp25_ASAP7_75t_L g9031 ( 
.A(n_8990),
.B(n_4932),
.C(n_5019),
.D(n_5001),
.Y(n_9031)
);

O2A1O1Ixp33_ASAP7_75t_SL g9032 ( 
.A1(n_8930),
.A2(n_5079),
.B(n_4782),
.C(n_4840),
.Y(n_9032)
);

OAI22xp5_ASAP7_75t_L g9033 ( 
.A1(n_8928),
.A2(n_8975),
.B1(n_8958),
.B2(n_8967),
.Y(n_9033)
);

NOR4xp25_ASAP7_75t_L g9034 ( 
.A(n_8948),
.B(n_8935),
.C(n_8945),
.D(n_8952),
.Y(n_9034)
);

AOI21xp5_ASAP7_75t_L g9035 ( 
.A1(n_8973),
.A2(n_8976),
.B(n_8987),
.Y(n_9035)
);

OAI21xp33_ASAP7_75t_L g9036 ( 
.A1(n_8955),
.A2(n_5001),
.B(n_4932),
.Y(n_9036)
);

OAI221xp5_ASAP7_75t_L g9037 ( 
.A1(n_8981),
.A2(n_4917),
.B1(n_4937),
.B2(n_4872),
.C(n_4788),
.Y(n_9037)
);

AOI211xp5_ASAP7_75t_L g9038 ( 
.A1(n_8956),
.A2(n_4820),
.B(n_4858),
.C(n_4836),
.Y(n_9038)
);

NAND2xp5_ASAP7_75t_L g9039 ( 
.A(n_8962),
.B(n_5206),
.Y(n_9039)
);

INVx1_ASAP7_75t_L g9040 ( 
.A(n_8962),
.Y(n_9040)
);

INVx1_ASAP7_75t_L g9041 ( 
.A(n_8974),
.Y(n_9041)
);

AOI221xp5_ASAP7_75t_L g9042 ( 
.A1(n_8984),
.A2(n_4834),
.B1(n_4847),
.B2(n_4841),
.C(n_4840),
.Y(n_9042)
);

AO22x2_ASAP7_75t_L g9043 ( 
.A1(n_8988),
.A2(n_4834),
.B1(n_4841),
.B2(n_4840),
.Y(n_9043)
);

AOI211xp5_ASAP7_75t_L g9044 ( 
.A1(n_8964),
.A2(n_4820),
.B(n_4858),
.C(n_4836),
.Y(n_9044)
);

O2A1O1Ixp33_ASAP7_75t_L g9045 ( 
.A1(n_8979),
.A2(n_4872),
.B(n_4937),
.C(n_4917),
.Y(n_9045)
);

OAI211xp5_ASAP7_75t_SL g9046 ( 
.A1(n_8969),
.A2(n_4841),
.B(n_4847),
.C(n_4834),
.Y(n_9046)
);

AOI21xp33_ASAP7_75t_L g9047 ( 
.A1(n_8991),
.A2(n_4915),
.B(n_5395),
.Y(n_9047)
);

AOI222xp33_ASAP7_75t_L g9048 ( 
.A1(n_8964),
.A2(n_5019),
.B1(n_5001),
.B2(n_4932),
.C1(n_4978),
.C2(n_4985),
.Y(n_9048)
);

O2A1O1Ixp5_ASAP7_75t_L g9049 ( 
.A1(n_8942),
.A2(n_4849),
.B(n_4976),
.C(n_4847),
.Y(n_9049)
);

INVxp67_ASAP7_75t_L g9050 ( 
.A(n_9009),
.Y(n_9050)
);

AOI22xp5_ASAP7_75t_L g9051 ( 
.A1(n_9002),
.A2(n_8953),
.B1(n_4835),
.B2(n_4837),
.Y(n_9051)
);

OAI22xp5_ASAP7_75t_L g9052 ( 
.A1(n_9018),
.A2(n_4976),
.B1(n_4978),
.B2(n_4849),
.Y(n_9052)
);

AND2x4_ASAP7_75t_L g9053 ( 
.A(n_9007),
.B(n_4820),
.Y(n_9053)
);

INVx1_ASAP7_75t_L g9054 ( 
.A(n_9015),
.Y(n_9054)
);

AND2x2_ASAP7_75t_L g9055 ( 
.A(n_9022),
.B(n_4853),
.Y(n_9055)
);

INVx1_ASAP7_75t_L g9056 ( 
.A(n_9020),
.Y(n_9056)
);

INVx1_ASAP7_75t_L g9057 ( 
.A(n_9012),
.Y(n_9057)
);

INVx1_ASAP7_75t_L g9058 ( 
.A(n_9004),
.Y(n_9058)
);

AND2x4_ASAP7_75t_L g9059 ( 
.A(n_9040),
.B(n_4836),
.Y(n_9059)
);

INVx1_ASAP7_75t_L g9060 ( 
.A(n_9043),
.Y(n_9060)
);

OAI21xp33_ASAP7_75t_L g9061 ( 
.A1(n_8998),
.A2(n_5019),
.B(n_5001),
.Y(n_9061)
);

OAI21xp5_ASAP7_75t_L g9062 ( 
.A1(n_9013),
.A2(n_5404),
.B(n_5386),
.Y(n_9062)
);

O2A1O1Ixp33_ASAP7_75t_L g9063 ( 
.A1(n_9041),
.A2(n_4917),
.B(n_4941),
.C(n_4937),
.Y(n_9063)
);

NOR2x1_ASAP7_75t_L g9064 ( 
.A(n_8995),
.B(n_8996),
.Y(n_9064)
);

BUFx3_ASAP7_75t_L g9065 ( 
.A(n_9033),
.Y(n_9065)
);

OAI211xp5_ASAP7_75t_SL g9066 ( 
.A1(n_9024),
.A2(n_4976),
.B(n_4978),
.C(n_4849),
.Y(n_9066)
);

AOI22xp33_ASAP7_75t_L g9067 ( 
.A1(n_9031),
.A2(n_4701),
.B1(n_5019),
.B2(n_4801),
.Y(n_9067)
);

INVx1_ASAP7_75t_L g9068 ( 
.A(n_9043),
.Y(n_9068)
);

AOI22xp33_ASAP7_75t_L g9069 ( 
.A1(n_9047),
.A2(n_4701),
.B1(n_4801),
.B2(n_4835),
.Y(n_9069)
);

AOI221xp5_ASAP7_75t_L g9070 ( 
.A1(n_9034),
.A2(n_5041),
.B1(n_4858),
.B2(n_4836),
.C(n_4985),
.Y(n_9070)
);

NAND2xp5_ASAP7_75t_L g9071 ( 
.A(n_8997),
.B(n_5516),
.Y(n_9071)
);

OAI21xp5_ASAP7_75t_L g9072 ( 
.A1(n_9035),
.A2(n_5417),
.B(n_5411),
.Y(n_9072)
);

AOI21xp5_ASAP7_75t_L g9073 ( 
.A1(n_9019),
.A2(n_9039),
.B(n_9042),
.Y(n_9073)
);

NAND3xp33_ASAP7_75t_L g9074 ( 
.A(n_8994),
.B(n_5041),
.C(n_4858),
.Y(n_9074)
);

INVx1_ASAP7_75t_L g9075 ( 
.A(n_9032),
.Y(n_9075)
);

O2A1O1Ixp33_ASAP7_75t_L g9076 ( 
.A1(n_9027),
.A2(n_4917),
.B(n_4941),
.C(n_4937),
.Y(n_9076)
);

BUFx3_ASAP7_75t_L g9077 ( 
.A(n_9037),
.Y(n_9077)
);

AOI221x1_ASAP7_75t_L g9078 ( 
.A1(n_9046),
.A2(n_4990),
.B1(n_5010),
.B2(n_4985),
.C(n_4982),
.Y(n_9078)
);

NAND2xp5_ASAP7_75t_SL g9079 ( 
.A(n_9005),
.B(n_4858),
.Y(n_9079)
);

INVx2_ASAP7_75t_L g9080 ( 
.A(n_9049),
.Y(n_9080)
);

AOI222xp33_ASAP7_75t_L g9081 ( 
.A1(n_9021),
.A2(n_5013),
.B1(n_5043),
.B2(n_5026),
.C1(n_5010),
.C2(n_4990),
.Y(n_9081)
);

INVxp67_ASAP7_75t_L g9082 ( 
.A(n_9008),
.Y(n_9082)
);

AOI21xp5_ASAP7_75t_L g9083 ( 
.A1(n_9045),
.A2(n_4701),
.B(n_4620),
.Y(n_9083)
);

INVx1_ASAP7_75t_L g9084 ( 
.A(n_9001),
.Y(n_9084)
);

NAND3xp33_ASAP7_75t_L g9085 ( 
.A(n_9044),
.B(n_5041),
.C(n_4858),
.Y(n_9085)
);

INVx1_ASAP7_75t_L g9086 ( 
.A(n_9011),
.Y(n_9086)
);

INVx1_ASAP7_75t_L g9087 ( 
.A(n_9026),
.Y(n_9087)
);

AOI21xp33_ASAP7_75t_SL g9088 ( 
.A1(n_9025),
.A2(n_4953),
.B(n_4941),
.Y(n_9088)
);

OAI22xp5_ASAP7_75t_L g9089 ( 
.A1(n_9038),
.A2(n_4990),
.B1(n_5010),
.B2(n_4982),
.Y(n_9089)
);

INVx1_ASAP7_75t_L g9090 ( 
.A(n_9029),
.Y(n_9090)
);

AOI22xp5_ASAP7_75t_L g9091 ( 
.A1(n_9036),
.A2(n_5041),
.B1(n_4858),
.B2(n_4950),
.Y(n_9091)
);

CKINVDCx20_ASAP7_75t_R g9092 ( 
.A(n_9003),
.Y(n_9092)
);

O2A1O1Ixp5_ASAP7_75t_SL g9093 ( 
.A1(n_9006),
.A2(n_5013),
.B(n_5026),
.C(n_4982),
.Y(n_9093)
);

OAI21xp33_ASAP7_75t_SL g9094 ( 
.A1(n_9016),
.A2(n_5052),
.B(n_4656),
.Y(n_9094)
);

NAND3xp33_ASAP7_75t_SL g9095 ( 
.A(n_9050),
.B(n_9014),
.C(n_9028),
.Y(n_9095)
);

A2O1A1Ixp33_ASAP7_75t_L g9096 ( 
.A1(n_9054),
.A2(n_9000),
.B(n_8999),
.C(n_9030),
.Y(n_9096)
);

NAND3xp33_ASAP7_75t_SL g9097 ( 
.A(n_9056),
.B(n_9017),
.C(n_9010),
.Y(n_9097)
);

OAI211xp5_ASAP7_75t_L g9098 ( 
.A1(n_9064),
.A2(n_9048),
.B(n_9023),
.C(n_5041),
.Y(n_9098)
);

NAND2xp5_ASAP7_75t_SL g9099 ( 
.A(n_9065),
.B(n_9053),
.Y(n_9099)
);

NOR2x1p5_ASAP7_75t_L g9100 ( 
.A(n_9087),
.B(n_5041),
.Y(n_9100)
);

NAND3xp33_ASAP7_75t_SL g9101 ( 
.A(n_9058),
.B(n_4953),
.C(n_4941),
.Y(n_9101)
);

OAI211xp5_ASAP7_75t_L g9102 ( 
.A1(n_9086),
.A2(n_5041),
.B(n_4986),
.C(n_5609),
.Y(n_9102)
);

AND2x2_ASAP7_75t_SL g9103 ( 
.A(n_9080),
.B(n_5041),
.Y(n_9103)
);

NAND3xp33_ASAP7_75t_L g9104 ( 
.A(n_9057),
.B(n_4974),
.C(n_4993),
.Y(n_9104)
);

AOI21xp5_ASAP7_75t_L g9105 ( 
.A1(n_9060),
.A2(n_4620),
.B(n_5411),
.Y(n_9105)
);

HB1xp67_ASAP7_75t_L g9106 ( 
.A(n_9053),
.Y(n_9106)
);

OAI211xp5_ASAP7_75t_SL g9107 ( 
.A1(n_9068),
.A2(n_9090),
.B(n_9073),
.C(n_9075),
.Y(n_9107)
);

A2O1A1Ixp33_ASAP7_75t_L g9108 ( 
.A1(n_9084),
.A2(n_4619),
.B(n_4668),
.C(n_4650),
.Y(n_9108)
);

INVx1_ASAP7_75t_L g9109 ( 
.A(n_9059),
.Y(n_9109)
);

AND4x1_ASAP7_75t_L g9110 ( 
.A(n_9071),
.B(n_5617),
.C(n_5627),
.D(n_5621),
.Y(n_9110)
);

OAI211xp5_ASAP7_75t_L g9111 ( 
.A1(n_9082),
.A2(n_4986),
.B(n_5026),
.C(n_5013),
.Y(n_9111)
);

AOI221xp5_ASAP7_75t_L g9112 ( 
.A1(n_9059),
.A2(n_5043),
.B1(n_4876),
.B2(n_4892),
.C(n_4888),
.Y(n_9112)
);

OR3x1_ASAP7_75t_L g9113 ( 
.A(n_9066),
.B(n_5043),
.C(n_4876),
.Y(n_9113)
);

OAI211xp5_ASAP7_75t_L g9114 ( 
.A1(n_9077),
.A2(n_4986),
.B(n_5426),
.C(n_5417),
.Y(n_9114)
);

A2O1A1Ixp33_ASAP7_75t_L g9115 ( 
.A1(n_9074),
.A2(n_4619),
.B(n_4668),
.C(n_4650),
.Y(n_9115)
);

AOI21xp5_ASAP7_75t_L g9116 ( 
.A1(n_9092),
.A2(n_4620),
.B(n_5426),
.Y(n_9116)
);

XNOR2x1_ASAP7_75t_L g9117 ( 
.A(n_9085),
.B(n_4953),
.Y(n_9117)
);

NAND5xp2_ASAP7_75t_L g9118 ( 
.A(n_9061),
.B(n_4954),
.C(n_4953),
.D(n_4720),
.E(n_4724),
.Y(n_9118)
);

NOR3xp33_ASAP7_75t_SL g9119 ( 
.A(n_9079),
.B(n_4888),
.C(n_4875),
.Y(n_9119)
);

AOI221xp5_ASAP7_75t_L g9120 ( 
.A1(n_9088),
.A2(n_4894),
.B1(n_4906),
.B2(n_4901),
.C(n_4892),
.Y(n_9120)
);

AOI22xp5_ASAP7_75t_L g9121 ( 
.A1(n_9062),
.A2(n_4950),
.B1(n_4952),
.B2(n_4986),
.Y(n_9121)
);

NOR3xp33_ASAP7_75t_SL g9122 ( 
.A(n_9052),
.B(n_9094),
.C(n_9070),
.Y(n_9122)
);

AOI211x1_ASAP7_75t_SL g9123 ( 
.A1(n_9083),
.A2(n_5516),
.B(n_4853),
.C(n_5138),
.Y(n_9123)
);

NOR2xp67_ASAP7_75t_L g9124 ( 
.A(n_9089),
.B(n_4780),
.Y(n_9124)
);

NOR4xp25_ASAP7_75t_L g9125 ( 
.A(n_9067),
.B(n_4894),
.C(n_4906),
.D(n_4901),
.Y(n_9125)
);

INVx1_ASAP7_75t_L g9126 ( 
.A(n_9078),
.Y(n_9126)
);

OAI211xp5_ASAP7_75t_L g9127 ( 
.A1(n_9081),
.A2(n_4986),
.B(n_4731),
.C(n_4922),
.Y(n_9127)
);

NAND2xp5_ASAP7_75t_L g9128 ( 
.A(n_9093),
.B(n_5516),
.Y(n_9128)
);

AOI221xp5_ASAP7_75t_L g9129 ( 
.A1(n_9072),
.A2(n_4922),
.B1(n_4933),
.B2(n_4927),
.C(n_4918),
.Y(n_9129)
);

OAI21xp33_ASAP7_75t_L g9130 ( 
.A1(n_9069),
.A2(n_4780),
.B(n_4954),
.Y(n_9130)
);

INVx1_ASAP7_75t_L g9131 ( 
.A(n_9051),
.Y(n_9131)
);

NAND2xp5_ASAP7_75t_L g9132 ( 
.A(n_9076),
.B(n_9091),
.Y(n_9132)
);

AOI221xp5_ASAP7_75t_L g9133 ( 
.A1(n_9063),
.A2(n_4927),
.B1(n_4935),
.B2(n_4933),
.C(n_4918),
.Y(n_9133)
);

AOI221xp5_ASAP7_75t_L g9134 ( 
.A1(n_9055),
.A2(n_4938),
.B1(n_5051),
.B2(n_4942),
.C(n_4935),
.Y(n_9134)
);

NAND4xp75_ASAP7_75t_L g9135 ( 
.A(n_9064),
.B(n_4828),
.C(n_4934),
.D(n_4795),
.Y(n_9135)
);

INVx1_ASAP7_75t_L g9136 ( 
.A(n_9106),
.Y(n_9136)
);

NAND2xp5_ASAP7_75t_L g9137 ( 
.A(n_9109),
.B(n_5516),
.Y(n_9137)
);

INVx1_ASAP7_75t_L g9138 ( 
.A(n_9103),
.Y(n_9138)
);

AND2x4_ASAP7_75t_L g9139 ( 
.A(n_9099),
.B(n_5516),
.Y(n_9139)
);

AND3x2_ASAP7_75t_L g9140 ( 
.A(n_9126),
.B(n_4942),
.C(n_4938),
.Y(n_9140)
);

NAND2x1p5_ASAP7_75t_L g9141 ( 
.A(n_9131),
.B(n_4967),
.Y(n_9141)
);

INVx1_ASAP7_75t_L g9142 ( 
.A(n_9098),
.Y(n_9142)
);

NAND4xp75_ASAP7_75t_L g9143 ( 
.A(n_9132),
.B(n_4828),
.C(n_4934),
.D(n_4795),
.Y(n_9143)
);

NOR2x1_ASAP7_75t_L g9144 ( 
.A(n_9107),
.B(n_4952),
.Y(n_9144)
);

OAI22xp5_ASAP7_75t_L g9145 ( 
.A1(n_9100),
.A2(n_4954),
.B1(n_5053),
.B2(n_5051),
.Y(n_9145)
);

INVx1_ASAP7_75t_L g9146 ( 
.A(n_9128),
.Y(n_9146)
);

XOR2xp5_ASAP7_75t_L g9147 ( 
.A(n_9097),
.B(n_4954),
.Y(n_9147)
);

NOR2xp33_ASAP7_75t_L g9148 ( 
.A(n_9095),
.B(n_4780),
.Y(n_9148)
);

NOR3xp33_ASAP7_75t_L g9149 ( 
.A(n_9096),
.B(n_5076),
.C(n_4619),
.Y(n_9149)
);

INVx2_ASAP7_75t_SL g9150 ( 
.A(n_9117),
.Y(n_9150)
);

INVx2_ASAP7_75t_SL g9151 ( 
.A(n_9110),
.Y(n_9151)
);

XNOR2x1_ASAP7_75t_L g9152 ( 
.A(n_9124),
.B(n_4677),
.Y(n_9152)
);

NAND4xp75_ASAP7_75t_L g9153 ( 
.A(n_9122),
.B(n_4828),
.C(n_4795),
.D(n_4896),
.Y(n_9153)
);

NAND3xp33_ASAP7_75t_SL g9154 ( 
.A(n_9130),
.B(n_4697),
.C(n_4694),
.Y(n_9154)
);

INVx1_ASAP7_75t_L g9155 ( 
.A(n_9113),
.Y(n_9155)
);

NOR2xp67_ASAP7_75t_L g9156 ( 
.A(n_9101),
.B(n_5053),
.Y(n_9156)
);

INVx1_ASAP7_75t_L g9157 ( 
.A(n_9119),
.Y(n_9157)
);

XNOR2xp5_ASAP7_75t_L g9158 ( 
.A(n_9125),
.B(n_9104),
.Y(n_9158)
);

INVx2_ASAP7_75t_L g9159 ( 
.A(n_9135),
.Y(n_9159)
);

INVx1_ASAP7_75t_L g9160 ( 
.A(n_9134),
.Y(n_9160)
);

INVx1_ASAP7_75t_L g9161 ( 
.A(n_9127),
.Y(n_9161)
);

AND2x2_ASAP7_75t_SL g9162 ( 
.A(n_9120),
.B(n_4828),
.Y(n_9162)
);

AND2x4_ASAP7_75t_L g9163 ( 
.A(n_9116),
.B(n_4868),
.Y(n_9163)
);

NOR3xp33_ASAP7_75t_L g9164 ( 
.A(n_9118),
.B(n_5076),
.C(n_4968),
.Y(n_9164)
);

INVxp33_ASAP7_75t_SL g9165 ( 
.A(n_9133),
.Y(n_9165)
);

INVx1_ASAP7_75t_L g9166 ( 
.A(n_9129),
.Y(n_9166)
);

INVx2_ASAP7_75t_L g9167 ( 
.A(n_9136),
.Y(n_9167)
);

NOR2x1_ASAP7_75t_L g9168 ( 
.A(n_9142),
.B(n_9111),
.Y(n_9168)
);

NOR2x1p5_ASAP7_75t_L g9169 ( 
.A(n_9155),
.B(n_9123),
.Y(n_9169)
);

NOR3xp33_ASAP7_75t_L g9170 ( 
.A(n_9146),
.B(n_9102),
.C(n_9114),
.Y(n_9170)
);

OAI221xp5_ASAP7_75t_L g9171 ( 
.A1(n_9138),
.A2(n_9150),
.B1(n_9147),
.B2(n_9158),
.C(n_9161),
.Y(n_9171)
);

INVx1_ASAP7_75t_L g9172 ( 
.A(n_9148),
.Y(n_9172)
);

AND2x4_ASAP7_75t_L g9173 ( 
.A(n_9151),
.B(n_9105),
.Y(n_9173)
);

INVx1_ASAP7_75t_L g9174 ( 
.A(n_9137),
.Y(n_9174)
);

AO211x2_ASAP7_75t_L g9175 ( 
.A1(n_9157),
.A2(n_9115),
.B(n_9121),
.C(n_9112),
.Y(n_9175)
);

OR5x1_ASAP7_75t_L g9176 ( 
.A(n_9154),
.B(n_9108),
.C(n_4853),
.D(n_5138),
.E(n_4652),
.Y(n_9176)
);

OAI22x1_ASAP7_75t_L g9177 ( 
.A1(n_9159),
.A2(n_9166),
.B1(n_9160),
.B2(n_9139),
.Y(n_9177)
);

NAND5xp2_ASAP7_75t_L g9178 ( 
.A(n_9165),
.B(n_4697),
.C(n_4720),
.D(n_4724),
.E(n_4751),
.Y(n_9178)
);

AND2x4_ASAP7_75t_L g9179 ( 
.A(n_9163),
.B(n_4868),
.Y(n_9179)
);

NOR4xp75_ASAP7_75t_SL g9180 ( 
.A(n_9145),
.B(n_9140),
.C(n_9156),
.D(n_9149),
.Y(n_9180)
);

OAI22xp5_ASAP7_75t_L g9181 ( 
.A1(n_9163),
.A2(n_9152),
.B1(n_9162),
.B2(n_9144),
.Y(n_9181)
);

NOR3xp33_ASAP7_75t_L g9182 ( 
.A(n_9139),
.B(n_5076),
.C(n_4968),
.Y(n_9182)
);

NAND5xp2_ASAP7_75t_L g9183 ( 
.A(n_9164),
.B(n_4694),
.C(n_4720),
.D(n_4697),
.E(n_4724),
.Y(n_9183)
);

NOR3xp33_ASAP7_75t_SL g9184 ( 
.A(n_9153),
.B(n_5061),
.C(n_5058),
.Y(n_9184)
);

NOR3xp33_ASAP7_75t_L g9185 ( 
.A(n_9143),
.B(n_4968),
.C(n_4967),
.Y(n_9185)
);

AND5x1_ASAP7_75t_L g9186 ( 
.A(n_9141),
.B(n_5138),
.C(n_4638),
.D(n_4887),
.E(n_4652),
.Y(n_9186)
);

NOR4xp25_ASAP7_75t_L g9187 ( 
.A(n_9136),
.B(n_5061),
.C(n_5065),
.D(n_5058),
.Y(n_9187)
);

OR2x2_ASAP7_75t_L g9188 ( 
.A(n_9167),
.B(n_5138),
.Y(n_9188)
);

HB1xp67_ASAP7_75t_L g9189 ( 
.A(n_9177),
.Y(n_9189)
);

CKINVDCx16_ASAP7_75t_R g9190 ( 
.A(n_9172),
.Y(n_9190)
);

BUFx2_ASAP7_75t_L g9191 ( 
.A(n_9168),
.Y(n_9191)
);

NAND2xp5_ASAP7_75t_L g9192 ( 
.A(n_9181),
.B(n_5138),
.Y(n_9192)
);

INVx2_ASAP7_75t_L g9193 ( 
.A(n_9169),
.Y(n_9193)
);

BUFx2_ASAP7_75t_L g9194 ( 
.A(n_9174),
.Y(n_9194)
);

OAI221xp5_ASAP7_75t_SL g9195 ( 
.A1(n_9171),
.A2(n_4677),
.B1(n_5000),
.B2(n_5008),
.C(n_4995),
.Y(n_9195)
);

BUFx2_ASAP7_75t_L g9196 ( 
.A(n_9173),
.Y(n_9196)
);

INVx1_ASAP7_75t_L g9197 ( 
.A(n_9170),
.Y(n_9197)
);

BUFx3_ASAP7_75t_L g9198 ( 
.A(n_9179),
.Y(n_9198)
);

HB1xp67_ASAP7_75t_L g9199 ( 
.A(n_9175),
.Y(n_9199)
);

INVx1_ASAP7_75t_SL g9200 ( 
.A(n_9180),
.Y(n_9200)
);

BUFx2_ASAP7_75t_L g9201 ( 
.A(n_9184),
.Y(n_9201)
);

CKINVDCx5p33_ASAP7_75t_R g9202 ( 
.A(n_9185),
.Y(n_9202)
);

BUFx2_ASAP7_75t_L g9203 ( 
.A(n_9183),
.Y(n_9203)
);

INVx2_ASAP7_75t_L g9204 ( 
.A(n_9176),
.Y(n_9204)
);

BUFx2_ASAP7_75t_L g9205 ( 
.A(n_9187),
.Y(n_9205)
);

NOR3xp33_ASAP7_75t_L g9206 ( 
.A(n_9182),
.B(n_4971),
.C(n_4967),
.Y(n_9206)
);

AOI22xp5_ASAP7_75t_L g9207 ( 
.A1(n_9191),
.A2(n_9186),
.B1(n_9178),
.B2(n_4952),
.Y(n_9207)
);

NOR4xp25_ASAP7_75t_L g9208 ( 
.A(n_9200),
.B(n_5068),
.C(n_5065),
.D(n_5007),
.Y(n_9208)
);

INVx2_ASAP7_75t_L g9209 ( 
.A(n_9199),
.Y(n_9209)
);

NOR4xp25_ASAP7_75t_L g9210 ( 
.A(n_9197),
.B(n_5068),
.C(n_5007),
.D(n_4993),
.Y(n_9210)
);

NAND4xp75_ASAP7_75t_L g9211 ( 
.A(n_9197),
.B(n_4896),
.C(n_4828),
.D(n_4795),
.Y(n_9211)
);

AOI22xp5_ASAP7_75t_L g9212 ( 
.A1(n_9189),
.A2(n_4952),
.B1(n_4950),
.B2(n_4959),
.Y(n_9212)
);

AND3x2_ASAP7_75t_L g9213 ( 
.A(n_9196),
.B(n_4904),
.C(n_4868),
.Y(n_9213)
);

INVx2_ASAP7_75t_L g9214 ( 
.A(n_9205),
.Y(n_9214)
);

AND2x2_ASAP7_75t_SL g9215 ( 
.A(n_9190),
.B(n_4896),
.Y(n_9215)
);

OR2x2_ASAP7_75t_L g9216 ( 
.A(n_9194),
.B(n_4887),
.Y(n_9216)
);

AND4x1_ASAP7_75t_L g9217 ( 
.A(n_9192),
.B(n_4887),
.C(n_4708),
.D(n_4652),
.Y(n_9217)
);

INVx1_ASAP7_75t_L g9218 ( 
.A(n_9203),
.Y(n_9218)
);

XNOR2xp5_ASAP7_75t_L g9219 ( 
.A(n_9193),
.B(n_4677),
.Y(n_9219)
);

NAND2xp5_ASAP7_75t_L g9220 ( 
.A(n_9198),
.B(n_4887),
.Y(n_9220)
);

AND3x4_ASAP7_75t_L g9221 ( 
.A(n_9204),
.B(n_4904),
.C(n_4868),
.Y(n_9221)
);

AND2x4_ASAP7_75t_L g9222 ( 
.A(n_9201),
.B(n_4868),
.Y(n_9222)
);

OR2x2_ASAP7_75t_L g9223 ( 
.A(n_9202),
.B(n_4887),
.Y(n_9223)
);

AND2x2_ASAP7_75t_L g9224 ( 
.A(n_9206),
.B(n_4904),
.Y(n_9224)
);

NAND2xp5_ASAP7_75t_L g9225 ( 
.A(n_9188),
.B(n_4887),
.Y(n_9225)
);

INVx2_ASAP7_75t_SL g9226 ( 
.A(n_9195),
.Y(n_9226)
);

INVx2_ASAP7_75t_L g9227 ( 
.A(n_9209),
.Y(n_9227)
);

NAND5xp2_ASAP7_75t_L g9228 ( 
.A(n_9218),
.B(n_4751),
.C(n_4697),
.D(n_4720),
.E(n_4724),
.Y(n_9228)
);

AND2x2_ASAP7_75t_SL g9229 ( 
.A(n_9214),
.B(n_4896),
.Y(n_9229)
);

OAI221xp5_ASAP7_75t_L g9230 ( 
.A1(n_9226),
.A2(n_4694),
.B1(n_4751),
.B2(n_4677),
.C(n_5000),
.Y(n_9230)
);

NOR2x1_ASAP7_75t_L g9231 ( 
.A(n_9222),
.B(n_4952),
.Y(n_9231)
);

AO22x2_ASAP7_75t_L g9232 ( 
.A1(n_9221),
.A2(n_4708),
.B1(n_4692),
.B2(n_5007),
.Y(n_9232)
);

NAND4xp25_ASAP7_75t_SL g9233 ( 
.A(n_9207),
.B(n_9225),
.C(n_9224),
.D(n_9220),
.Y(n_9233)
);

AOI22xp5_ASAP7_75t_L g9234 ( 
.A1(n_9219),
.A2(n_4950),
.B1(n_5017),
.B2(n_4959),
.Y(n_9234)
);

HB1xp67_ASAP7_75t_L g9235 ( 
.A(n_9208),
.Y(n_9235)
);

INVx1_ASAP7_75t_L g9236 ( 
.A(n_9213),
.Y(n_9236)
);

AND3x1_ASAP7_75t_L g9237 ( 
.A(n_9210),
.B(n_4887),
.C(n_4652),
.Y(n_9237)
);

INVx1_ASAP7_75t_L g9238 ( 
.A(n_9215),
.Y(n_9238)
);

OAI211xp5_ASAP7_75t_SL g9239 ( 
.A1(n_9212),
.A2(n_4931),
.B(n_4939),
.C(n_4826),
.Y(n_9239)
);

AOI22xp33_ASAP7_75t_SL g9240 ( 
.A1(n_9216),
.A2(n_9223),
.B1(n_9211),
.B2(n_9217),
.Y(n_9240)
);

OR4x2_ASAP7_75t_L g9241 ( 
.A(n_9209),
.B(n_4887),
.C(n_4652),
.D(n_4692),
.Y(n_9241)
);

OR2x2_ASAP7_75t_L g9242 ( 
.A(n_9227),
.B(n_9238),
.Y(n_9242)
);

INVx2_ASAP7_75t_L g9243 ( 
.A(n_9235),
.Y(n_9243)
);

AOI22xp5_ASAP7_75t_L g9244 ( 
.A1(n_9236),
.A2(n_4950),
.B1(n_5017),
.B2(n_4959),
.Y(n_9244)
);

AOI22xp5_ASAP7_75t_L g9245 ( 
.A1(n_9233),
.A2(n_4959),
.B1(n_5017),
.B2(n_4801),
.Y(n_9245)
);

OA22x2_ASAP7_75t_L g9246 ( 
.A1(n_9240),
.A2(n_4692),
.B1(n_4604),
.B2(n_4668),
.Y(n_9246)
);

OAI22x1_ASAP7_75t_L g9247 ( 
.A1(n_9231),
.A2(n_4751),
.B1(n_4694),
.B2(n_4896),
.Y(n_9247)
);

AND2x2_ASAP7_75t_SL g9248 ( 
.A(n_9229),
.B(n_4904),
.Y(n_9248)
);

XNOR2xp5_ASAP7_75t_L g9249 ( 
.A(n_9232),
.B(n_9237),
.Y(n_9249)
);

INVx1_ASAP7_75t_L g9250 ( 
.A(n_9239),
.Y(n_9250)
);

INVx1_ASAP7_75t_L g9251 ( 
.A(n_9234),
.Y(n_9251)
);

XNOR2xp5_ASAP7_75t_L g9252 ( 
.A(n_9230),
.B(n_9228),
.Y(n_9252)
);

INVx2_ASAP7_75t_L g9253 ( 
.A(n_9241),
.Y(n_9253)
);

AND2x4_ASAP7_75t_L g9254 ( 
.A(n_9243),
.B(n_4904),
.Y(n_9254)
);

XNOR2xp5_ASAP7_75t_L g9255 ( 
.A(n_9242),
.B(n_4983),
.Y(n_9255)
);

AOI22x1_ASAP7_75t_L g9256 ( 
.A1(n_9253),
.A2(n_2722),
.B1(n_2696),
.B2(n_2474),
.Y(n_9256)
);

NAND2xp5_ASAP7_75t_L g9257 ( 
.A(n_9249),
.B(n_4638),
.Y(n_9257)
);

INVx3_ASAP7_75t_SL g9258 ( 
.A(n_9251),
.Y(n_9258)
);

OAI22xp33_ASAP7_75t_L g9259 ( 
.A1(n_9250),
.A2(n_4931),
.B1(n_4939),
.B2(n_4826),
.Y(n_9259)
);

OAI22xp5_ASAP7_75t_L g9260 ( 
.A1(n_9252),
.A2(n_5000),
.B1(n_5008),
.B2(n_4995),
.Y(n_9260)
);

AOI22xp5_ASAP7_75t_L g9261 ( 
.A1(n_9258),
.A2(n_9248),
.B1(n_9247),
.B2(n_9245),
.Y(n_9261)
);

OAI22xp33_ASAP7_75t_L g9262 ( 
.A1(n_9254),
.A2(n_9246),
.B1(n_9244),
.B2(n_5000),
.Y(n_9262)
);

OAI22xp5_ASAP7_75t_L g9263 ( 
.A1(n_9255),
.A2(n_5000),
.B1(n_5008),
.B2(n_4995),
.Y(n_9263)
);

OAI22xp5_ASAP7_75t_SL g9264 ( 
.A1(n_9257),
.A2(n_5000),
.B1(n_5008),
.B2(n_4995),
.Y(n_9264)
);

INVx2_ASAP7_75t_L g9265 ( 
.A(n_9261),
.Y(n_9265)
);

INVx1_ASAP7_75t_L g9266 ( 
.A(n_9262),
.Y(n_9266)
);

AND3x1_ASAP7_75t_L g9267 ( 
.A(n_9264),
.B(n_9256),
.C(n_9260),
.Y(n_9267)
);

OAI21x1_ASAP7_75t_L g9268 ( 
.A1(n_9265),
.A2(n_9263),
.B(n_9259),
.Y(n_9268)
);

AOI21xp5_ASAP7_75t_L g9269 ( 
.A1(n_9268),
.A2(n_9266),
.B(n_9267),
.Y(n_9269)
);

AOI21xp33_ASAP7_75t_L g9270 ( 
.A1(n_9269),
.A2(n_2479),
.B(n_2371),
.Y(n_9270)
);

AOI22xp5_ASAP7_75t_L g9271 ( 
.A1(n_9270),
.A2(n_5000),
.B1(n_5008),
.B2(n_4995),
.Y(n_9271)
);

AO21x2_ASAP7_75t_L g9272 ( 
.A1(n_9271),
.A2(n_4656),
.B(n_4971),
.Y(n_9272)
);

OAI221xp5_ASAP7_75t_R g9273 ( 
.A1(n_9272),
.A2(n_4652),
.B1(n_4638),
.B2(n_4962),
.C(n_4928),
.Y(n_9273)
);

OAI221xp5_ASAP7_75t_R g9274 ( 
.A1(n_9272),
.A2(n_4652),
.B1(n_4638),
.B2(n_4962),
.C(n_4928),
.Y(n_9274)
);

AOI22xp5_ASAP7_75t_L g9275 ( 
.A1(n_9273),
.A2(n_4929),
.B1(n_5008),
.B2(n_4995),
.Y(n_9275)
);

AOI211xp5_ASAP7_75t_L g9276 ( 
.A1(n_9275),
.A2(n_9274),
.B(n_2474),
.C(n_2501),
.Y(n_9276)
);


endmodule