module fake_jpeg_25252_n_315 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_315);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_29),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_16),
.B1(n_20),
.B2(n_17),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_24),
.B1(n_27),
.B2(n_25),
.Y(n_59)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_50),
.B1(n_62),
.B2(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_16),
.B1(n_20),
.B2(n_33),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_33),
.B1(n_24),
.B2(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_61),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_25),
.B1(n_27),
.B2(n_11),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_25),
.B1(n_11),
.B2(n_15),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx2_ASAP7_75t_SL g82 ( 
.A(n_65),
.Y(n_82)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_36),
.B1(n_38),
.B2(n_37),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_77),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_58),
.B(n_50),
.C(n_62),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_22),
.B(n_29),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_57),
.B(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_30),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_38),
.B1(n_37),
.B2(n_46),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_66),
.B1(n_45),
.B2(n_42),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_60),
.B1(n_59),
.B2(n_56),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_94),
.B1(n_99),
.B2(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_90),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_28),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_91),
.B(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_48),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_101),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_0),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_65),
.B1(n_49),
.B2(n_64),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_53),
.B1(n_55),
.B2(n_42),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_107),
.B(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_55),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_77),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_69),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_31),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_84),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_69),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_58),
.B(n_1),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_111),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_83),
.C(n_76),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_126),
.C(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_116),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_70),
.B1(n_75),
.B2(n_79),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_115),
.A2(n_117),
.B(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_74),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_122),
.B(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_124),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_72),
.C(n_53),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_134),
.B1(n_138),
.B2(n_105),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_107),
.B(n_94),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_82),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_94),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_72),
.Y(n_133)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_87),
.A2(n_78),
.B1(n_72),
.B2(n_65),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_104),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_69),
.Y(n_136)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_15),
.B1(n_14),
.B2(n_26),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_87),
.A2(n_58),
.B1(n_69),
.B2(n_15),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_98),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_139),
.A2(n_153),
.B(n_131),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_111),
.B(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_140),
.B(n_163),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_146),
.B1(n_149),
.B2(n_156),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_126),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_99),
.B1(n_98),
.B2(n_101),
.Y(n_146)
);

OAI22x1_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_98),
.B1(n_94),
.B2(n_105),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_137),
.B1(n_135),
.B2(n_119),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_85),
.B1(n_98),
.B2(n_105),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_98),
.B1(n_94),
.B2(n_107),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_169),
.B1(n_119),
.B2(n_123),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_86),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_154),
.B(n_157),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_94),
.B1(n_86),
.B2(n_92),
.Y(n_156)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_117),
.B1(n_122),
.B2(n_108),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_179)
);

AOI32xp33_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_26),
.A3(n_32),
.B1(n_104),
.B2(n_68),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_123),
.C(n_124),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_68),
.B1(n_63),
.B2(n_13),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_67),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_63),
.B1(n_13),
.B2(n_21),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_114),
.A2(n_63),
.B1(n_13),
.B2(n_21),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_118),
.A2(n_63),
.B1(n_21),
.B2(n_14),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_118),
.A2(n_28),
.A3(n_18),
.B1(n_21),
.B2(n_23),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_110),
.A2(n_28),
.A3(n_18),
.B1(n_26),
.B2(n_32),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_131),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_110),
.Y(n_176)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_181),
.C(n_182),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_113),
.C(n_112),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_157),
.C(n_153),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_153),
.B(n_139),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_161),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_188),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_186),
.A2(n_199),
.B(n_200),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_195),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_132),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_112),
.C(n_132),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_190),
.B(n_155),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_128),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_192),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_196),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_63),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_67),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_67),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_139),
.A2(n_67),
.B(n_18),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_28),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_162),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_167),
.C(n_144),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_192),
.B1(n_189),
.B2(n_178),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_210),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_159),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_188),
.B(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_184),
.B(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_186),
.A2(n_142),
.B1(n_156),
.B2(n_149),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_173),
.B1(n_179),
.B2(n_195),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_144),
.B(n_152),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_219),
.A2(n_221),
.B(n_223),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_190),
.B(n_164),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_198),
.B(n_197),
.C(n_176),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_172),
.B(n_171),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_155),
.B(n_67),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_196),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_204),
.Y(n_244)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_229),
.A2(n_246),
.B1(n_218),
.B2(n_223),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_208),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_203),
.B(n_185),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_231),
.B(n_232),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_203),
.B(n_185),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_177),
.C(n_182),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_242),
.C(n_230),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_194),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_245),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_189),
.B1(n_178),
.B2(n_201),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_213),
.B1(n_207),
.B2(n_224),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_67),
.B1(n_28),
.B2(n_2),
.Y(n_240)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_28),
.C(n_1),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_214),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_0),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_259),
.B1(n_261),
.B2(n_245),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_250),
.B(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_253),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_212),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_260),
.C(n_3),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_221),
.B1(n_207),
.B2(n_222),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_262),
.B1(n_233),
.B2(n_246),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_206),
.B(n_219),
.Y(n_256)
);

OAI321xp33_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_209),
.B1(n_218),
.B2(n_204),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_209),
.B1(n_206),
.B2(n_205),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_237),
.C(n_238),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_274),
.C(n_275),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_265),
.B(n_272),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_232),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_271),
.Y(n_282)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_231),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_227),
.B1(n_235),
.B2(n_4),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_6),
.B(n_7),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_3),
.C(n_4),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_3),
.C(n_5),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_255),
.C(n_258),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_259),
.B1(n_261),
.B2(n_257),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_281),
.Y(n_292)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_258),
.C(n_6),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_284),
.C(n_276),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_5),
.C(n_6),
.Y(n_284)
);

OAI21x1_ASAP7_75t_SL g285 ( 
.A1(n_266),
.A2(n_5),
.B(n_6),
.Y(n_285)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_10),
.B(n_7),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_284),
.B(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_7),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_267),
.Y(n_290)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_268),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_282),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_295),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_271),
.B(n_8),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_298),
.C(n_287),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_302),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_278),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_293),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_289),
.B(n_294),
.Y(n_305)
);

O2A1O1Ixp33_ASAP7_75t_SL g308 ( 
.A1(n_305),
.A2(n_299),
.B(n_301),
.C(n_297),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_307),
.A2(n_306),
.B(n_300),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_309),
.B(n_8),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_310),
.A2(n_9),
.B(n_10),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_9),
.C(n_10),
.Y(n_312)
);

AND2x2_ASAP7_75t_SL g313 ( 
.A(n_312),
.B(n_9),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_9),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_10),
.C(n_212),
.Y(n_315)
);


endmodule