module real_aes_7960_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g242 ( .A1(n_0), .A2(n_243), .B(n_244), .C(n_247), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_1), .B(n_184), .Y(n_248) );
INVx1_ASAP7_75t_L g422 ( .A(n_2), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_3), .B(n_154), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_4), .A2(n_124), .B(n_127), .C(n_435), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_5), .A2(n_144), .B(n_475), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_6), .A2(n_144), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_7), .B(n_184), .Y(n_481) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_8), .A2(n_111), .B(n_164), .Y(n_163) );
AND2x6_ASAP7_75t_L g124 ( .A(n_9), .B(n_125), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g126 ( .A1(n_10), .A2(n_124), .B(n_127), .C(n_130), .Y(n_126) );
INVx1_ASAP7_75t_L g451 ( .A(n_11), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_12), .B(n_39), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_13), .B(n_134), .Y(n_437) );
INVx1_ASAP7_75t_L g116 ( .A(n_14), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_15), .B(n_154), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_16), .A2(n_132), .B(n_459), .C(n_461), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_17), .B(n_184), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_18), .B(n_208), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_19), .A2(n_127), .B(n_171), .C(n_204), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_20), .A2(n_136), .B(n_246), .C(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_21), .B(n_134), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_22), .B(n_134), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_23), .Y(n_509) );
INVx1_ASAP7_75t_L g501 ( .A(n_24), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_25), .A2(n_127), .B(n_167), .C(n_171), .Y(n_166) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_26), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_27), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_28), .Y(n_433) );
INVx1_ASAP7_75t_L g492 ( .A(n_29), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_30), .A2(n_144), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g122 ( .A(n_31), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_32), .A2(n_146), .B(n_157), .C(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_33), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_34), .A2(n_246), .B(n_478), .C(n_480), .Y(n_477) );
INVxp67_ASAP7_75t_L g493 ( .A(n_35), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_36), .B(n_169), .Y(n_168) );
CKINVDCx14_ASAP7_75t_R g476 ( .A(n_37), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_38), .A2(n_127), .B(n_171), .C(n_500), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_40), .A2(n_247), .B(n_449), .C(n_450), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_41), .B(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_42), .Y(n_139) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_43), .A2(n_68), .B1(n_101), .B2(n_694), .C1(n_699), .C2(n_700), .Y(n_100) );
INVx1_ASAP7_75t_L g699 ( .A(n_43), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_44), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_45), .B(n_144), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_46), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_47), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_48), .A2(n_146), .B(n_148), .C(n_157), .Y(n_145) );
INVx1_ASAP7_75t_L g245 ( .A(n_49), .Y(n_245) );
INVx1_ASAP7_75t_L g149 ( .A(n_50), .Y(n_149) );
INVx1_ASAP7_75t_L g466 ( .A(n_51), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_52), .B(n_144), .Y(n_143) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_53), .A2(n_99), .B1(n_704), .B2(n_713), .C1(n_726), .C2(n_732), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_53), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_53), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_54), .Y(n_211) );
CKINVDCx14_ASAP7_75t_R g447 ( .A(n_55), .Y(n_447) );
INVx1_ASAP7_75t_L g125 ( .A(n_56), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_57), .B(n_144), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_58), .B(n_184), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_59), .A2(n_178), .B(n_180), .C(n_182), .Y(n_177) );
INVx1_ASAP7_75t_L g115 ( .A(n_60), .Y(n_115) );
INVx1_ASAP7_75t_SL g479 ( .A(n_61), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_62), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_63), .B(n_154), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_64), .B(n_184), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_65), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g512 ( .A(n_66), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g241 ( .A(n_67), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_69), .B(n_151), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_70), .A2(n_127), .B(n_157), .C(n_218), .Y(n_217) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_71), .Y(n_176) );
INVx1_ASAP7_75t_L g708 ( .A(n_72), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_73), .A2(n_144), .B(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_74), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_75), .A2(n_144), .B(n_456), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_76), .A2(n_202), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g457 ( .A(n_77), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_78), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_79), .B(n_150), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_80), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_81), .A2(n_144), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g460 ( .A(n_82), .Y(n_460) );
INVx2_ASAP7_75t_L g113 ( .A(n_83), .Y(n_113) );
INVx1_ASAP7_75t_L g436 ( .A(n_84), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_85), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_86), .B(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g420 ( .A(n_87), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g693 ( .A(n_87), .Y(n_693) );
OR2x2_ASAP7_75t_L g712 ( .A(n_87), .B(n_703), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_88), .A2(n_127), .B(n_157), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_89), .B(n_144), .Y(n_190) );
INVx1_ASAP7_75t_L g193 ( .A(n_90), .Y(n_193) );
INVxp67_ASAP7_75t_L g181 ( .A(n_91), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_92), .B(n_111), .Y(n_452) );
INVx1_ASAP7_75t_L g118 ( .A(n_93), .Y(n_118) );
INVx1_ASAP7_75t_L g219 ( .A(n_94), .Y(n_219) );
INVx2_ASAP7_75t_L g469 ( .A(n_95), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_96), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g160 ( .A(n_97), .B(n_159), .Y(n_160) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_418), .B1(n_424), .B2(n_690), .Y(n_101) );
INVx2_ASAP7_75t_L g696 ( .A(n_102), .Y(n_696) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_102), .Y(n_717) );
OR3x1_ASAP7_75t_L g102 ( .A(n_103), .B(n_316), .C(n_381), .Y(n_102) );
NAND4xp25_ASAP7_75t_SL g103 ( .A(n_104), .B(n_257), .C(n_283), .D(n_306), .Y(n_103) );
AOI221xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_185), .B1(n_226), .B2(n_233), .C(n_249), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_106), .A2(n_250), .B1(n_274), .B2(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_161), .Y(n_106) );
INVx1_ASAP7_75t_SL g310 ( .A(n_107), .Y(n_310) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_141), .Y(n_107) );
OR2x2_ASAP7_75t_L g231 ( .A(n_108), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g252 ( .A(n_108), .B(n_162), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_108), .B(n_172), .Y(n_265) );
AND2x2_ASAP7_75t_L g282 ( .A(n_108), .B(n_141), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_108), .B(n_229), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_108), .B(n_281), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_108), .B(n_161), .Y(n_403) );
AOI211xp5_ASAP7_75t_SL g414 ( .A1(n_108), .A2(n_320), .B(n_415), .C(n_416), .Y(n_414) );
INVx5_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_109), .B(n_162), .Y(n_286) );
AND2x2_ASAP7_75t_L g289 ( .A(n_109), .B(n_163), .Y(n_289) );
OR2x2_ASAP7_75t_L g334 ( .A(n_109), .B(n_162), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_109), .B(n_172), .Y(n_343) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_117), .B(n_138), .Y(n_109) );
INVx3_ASAP7_75t_L g184 ( .A(n_110), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_110), .B(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_110), .A2(n_216), .B(n_224), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_110), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_110), .B(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_110), .B(n_504), .Y(n_503) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_110), .A2(n_508), .B(n_514), .Y(n_507) );
INVx4_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_111), .A2(n_165), .B(n_166), .Y(n_164) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_111), .Y(n_173) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g140 ( .A(n_112), .Y(n_140) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_113), .B(n_114), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_119), .B(n_126), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_119), .A2(n_433), .B(n_434), .Y(n_432) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_119), .A2(n_159), .B(n_498), .C(n_499), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_119), .A2(n_509), .B(n_510), .Y(n_508) );
NAND2x1p5_ASAP7_75t_L g119 ( .A(n_120), .B(n_124), .Y(n_119) );
AND2x4_ASAP7_75t_L g144 ( .A(n_120), .B(n_124), .Y(n_144) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_123), .Y(n_120) );
INVx1_ASAP7_75t_L g182 ( .A(n_121), .Y(n_182) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g128 ( .A(n_122), .Y(n_128) );
INVx1_ASAP7_75t_L g137 ( .A(n_122), .Y(n_137) );
INVx1_ASAP7_75t_L g129 ( .A(n_123), .Y(n_129) );
INVx3_ASAP7_75t_L g132 ( .A(n_123), .Y(n_132) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_123), .Y(n_134) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_123), .Y(n_152) );
INVx1_ASAP7_75t_L g169 ( .A(n_123), .Y(n_169) );
INVx4_ASAP7_75t_SL g158 ( .A(n_124), .Y(n_158) );
BUFx3_ASAP7_75t_L g171 ( .A(n_124), .Y(n_171) );
INVx5_ASAP7_75t_L g147 ( .A(n_127), .Y(n_147) );
AND2x6_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
BUFx3_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_128), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_133), .B(n_135), .Y(n_130) );
INVx5_ASAP7_75t_L g154 ( .A(n_132), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_132), .B(n_451), .Y(n_450) );
INVx4_ASAP7_75t_L g246 ( .A(n_134), .Y(n_246) );
INVx2_ASAP7_75t_L g449 ( .A(n_134), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_135), .A2(n_168), .B(n_170), .Y(n_167) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
INVx2_ASAP7_75t_L g486 ( .A(n_140), .Y(n_486) );
INVx5_ASAP7_75t_SL g232 ( .A(n_141), .Y(n_232) );
AND2x2_ASAP7_75t_L g251 ( .A(n_141), .B(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_141), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g337 ( .A(n_141), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g369 ( .A(n_141), .B(n_172), .Y(n_369) );
OR2x2_ASAP7_75t_L g375 ( .A(n_141), .B(n_265), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_141), .B(n_325), .Y(n_384) );
OR2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_160), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_145), .B(n_159), .Y(n_142) );
BUFx2_ASAP7_75t_L g202 ( .A(n_144), .Y(n_202) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_147), .A2(n_158), .B(n_176), .C(n_177), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g240 ( .A1(n_147), .A2(n_158), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g446 ( .A1(n_147), .A2(n_158), .B(n_447), .C(n_448), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_SL g456 ( .A1(n_147), .A2(n_158), .B(n_457), .C(n_458), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_147), .A2(n_158), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_147), .A2(n_158), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_147), .A2(n_158), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_153), .C(n_155), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_150), .A2(n_155), .B(n_193), .C(n_194), .Y(n_192) );
O2A1O1Ixp5_ASAP7_75t_L g435 ( .A1(n_150), .A2(n_436), .B(n_437), .C(n_438), .Y(n_435) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_150), .A2(n_438), .B(n_512), .C(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_154), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g243 ( .A(n_154), .Y(n_243) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_154), .A2(n_179), .B1(n_492), .B2(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_154), .A2(n_207), .B(n_501), .C(n_502), .Y(n_500) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g247 ( .A(n_156), .Y(n_247) );
INVx1_ASAP7_75t_L g461 ( .A(n_156), .Y(n_461) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_159), .A2(n_190), .B(n_191), .Y(n_189) );
INVx2_ASAP7_75t_L g209 ( .A(n_159), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_159), .Y(n_212) );
OA21x2_ASAP7_75t_L g444 ( .A1(n_159), .A2(n_445), .B(n_452), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_172), .Y(n_161) );
AND2x2_ASAP7_75t_L g266 ( .A(n_162), .B(n_232), .Y(n_266) );
INVx1_ASAP7_75t_SL g279 ( .A(n_162), .Y(n_279) );
OR2x2_ASAP7_75t_L g314 ( .A(n_162), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g320 ( .A(n_162), .B(n_172), .Y(n_320) );
AND2x2_ASAP7_75t_L g378 ( .A(n_162), .B(n_229), .Y(n_378) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_163), .B(n_232), .Y(n_305) );
INVx3_ASAP7_75t_L g229 ( .A(n_172), .Y(n_229) );
OR2x2_ASAP7_75t_L g271 ( .A(n_172), .B(n_232), .Y(n_271) );
AND2x2_ASAP7_75t_L g281 ( .A(n_172), .B(n_279), .Y(n_281) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_172), .Y(n_329) );
AND2x2_ASAP7_75t_L g338 ( .A(n_172), .B(n_252), .Y(n_338) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_183), .Y(n_172) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_173), .A2(n_455), .B(n_462), .Y(n_454) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_173), .A2(n_464), .B(n_470), .Y(n_463) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_173), .A2(n_474), .B(n_481), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_178), .A2(n_219), .B(n_220), .C(n_221), .Y(n_218) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_179), .B(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_179), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g207 ( .A(n_182), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_182), .B(n_491), .Y(n_490) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_184), .A2(n_239), .B(n_248), .Y(n_238) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_185), .A2(n_355), .B1(n_357), .B2(n_359), .C(n_362), .Y(n_354) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OR2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_197), .Y(n_186) );
AND2x2_ASAP7_75t_L g328 ( .A(n_187), .B(n_309), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_187), .B(n_387), .Y(n_391) );
OR2x2_ASAP7_75t_L g412 ( .A(n_187), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_187), .B(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx5_ASAP7_75t_L g259 ( .A(n_188), .Y(n_259) );
AND2x2_ASAP7_75t_L g336 ( .A(n_188), .B(n_199), .Y(n_336) );
AND2x2_ASAP7_75t_L g397 ( .A(n_188), .B(n_276), .Y(n_397) );
AND2x2_ASAP7_75t_L g410 ( .A(n_188), .B(n_229), .Y(n_410) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_195), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_213), .Y(n_197) );
AND2x4_ASAP7_75t_L g236 ( .A(n_198), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g255 ( .A(n_198), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g262 ( .A(n_198), .Y(n_262) );
AND2x2_ASAP7_75t_L g331 ( .A(n_198), .B(n_309), .Y(n_331) );
AND2x2_ASAP7_75t_L g341 ( .A(n_198), .B(n_259), .Y(n_341) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_198), .Y(n_349) );
AND2x2_ASAP7_75t_L g361 ( .A(n_198), .B(n_238), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_198), .B(n_293), .Y(n_365) );
AND2x2_ASAP7_75t_L g402 ( .A(n_198), .B(n_397), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_198), .B(n_276), .Y(n_413) );
OR2x2_ASAP7_75t_L g415 ( .A(n_198), .B(n_351), .Y(n_415) );
INVx5_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g301 ( .A(n_199), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g311 ( .A(n_199), .B(n_256), .Y(n_311) );
AND2x2_ASAP7_75t_L g323 ( .A(n_199), .B(n_238), .Y(n_323) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_199), .Y(n_353) );
AND2x4_ASAP7_75t_L g387 ( .A(n_199), .B(n_237), .Y(n_387) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_210), .Y(n_199) );
AOI21xp5_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_203), .B(n_208), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_209), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AO21x2_ASAP7_75t_L g431 ( .A1(n_212), .A2(n_432), .B(n_439), .Y(n_431) );
BUFx2_ASAP7_75t_L g235 ( .A(n_213), .Y(n_235) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g276 ( .A(n_214), .Y(n_276) );
AND2x2_ASAP7_75t_L g309 ( .A(n_214), .B(n_238), .Y(n_309) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g256 ( .A(n_215), .B(n_238), .Y(n_256) );
BUFx2_ASAP7_75t_L g302 ( .A(n_215), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_223), .Y(n_216) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx3_ASAP7_75t_L g480 ( .A(n_222), .Y(n_480) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_228), .B(n_310), .Y(n_389) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_229), .B(n_252), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_229), .B(n_232), .Y(n_291) );
AND2x2_ASAP7_75t_L g346 ( .A(n_229), .B(n_282), .Y(n_346) );
AOI221xp5_ASAP7_75t_SL g283 ( .A1(n_230), .A2(n_284), .B1(n_292), .B2(n_294), .C(n_298), .Y(n_283) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g278 ( .A(n_231), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g319 ( .A(n_231), .B(n_320), .Y(n_319) );
OAI321xp33_ASAP7_75t_L g326 ( .A1(n_231), .A2(n_285), .A3(n_327), .B1(n_329), .B2(n_330), .C(n_332), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_232), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_235), .B(n_387), .Y(n_405) );
AND2x2_ASAP7_75t_L g292 ( .A(n_236), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_236), .B(n_296), .Y(n_295) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_237), .Y(n_268) );
AND2x2_ASAP7_75t_L g275 ( .A(n_237), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_237), .B(n_350), .Y(n_380) );
INVx1_ASAP7_75t_L g417 ( .A(n_237), .Y(n_417) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_246), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g438 ( .A(n_247), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_253), .B(n_254), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_251), .A2(n_361), .B(n_410), .C(n_411), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_252), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_252), .B(n_290), .Y(n_356) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g299 ( .A(n_256), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_256), .B(n_259), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_256), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_256), .B(n_341), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_260), .B1(n_272), .B2(n_277), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g273 ( .A(n_259), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g296 ( .A(n_259), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g308 ( .A(n_259), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_259), .B(n_302), .Y(n_344) );
OR2x2_ASAP7_75t_L g351 ( .A(n_259), .B(n_276), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_259), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g401 ( .A(n_259), .B(n_387), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_263), .B1(n_267), .B2(n_269), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g307 ( .A(n_262), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_265), .A2(n_280), .B1(n_348), .B2(n_352), .Y(n_347) );
INVx1_ASAP7_75t_L g395 ( .A(n_266), .Y(n_395) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_270), .A2(n_307), .B1(n_310), .B2(n_311), .C(n_312), .Y(n_306) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g285 ( .A(n_271), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_275), .B(n_341), .Y(n_373) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_276), .Y(n_293) );
INVx1_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
NAND2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
AND2x2_ASAP7_75t_L g324 ( .A(n_282), .B(n_325), .Y(n_324) );
NAND2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx2_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AND2x2_ASAP7_75t_L g368 ( .A(n_289), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_292), .A2(n_318), .B1(n_321), .B2(n_324), .C(n_326), .Y(n_317) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_296), .B(n_353), .Y(n_352) );
AOI21xp33_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_300), .B(n_303), .Y(n_298) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g400 ( .A(n_303), .Y(n_400) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
OR2x2_ASAP7_75t_L g342 ( .A(n_305), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g363 ( .A(n_308), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_308), .B(n_368), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_311), .B(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND4xp25_ASAP7_75t_L g316 ( .A(n_317), .B(n_335), .C(n_354), .D(n_367), .Y(n_316) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_SL g325 ( .A(n_320), .Y(n_325) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g358 ( .A(n_329), .B(n_334), .Y(n_358) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B(n_339), .C(n_347), .Y(n_335) );
AOI211xp5_ASAP7_75t_L g406 ( .A1(n_337), .A2(n_379), .B(n_407), .C(n_414), .Y(n_406) );
INVx1_ASAP7_75t_SL g366 ( .A(n_338), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B1(n_344), .B2(n_345), .Y(n_339) );
INVx1_ASAP7_75t_L g370 ( .A(n_344), .Y(n_370) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_350), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_350), .B(n_361), .Y(n_394) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g371 ( .A(n_361), .Y(n_371) );
AOI21xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B(n_366), .Y(n_362) );
INVxp33_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI322xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .A3(n_371), .B1(n_372), .B2(n_374), .C1(n_376), .C2(n_379), .Y(n_367) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND3xp33_ASAP7_75t_SL g381 ( .A(n_382), .B(n_399), .C(n_406), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B1(n_388), .B2(n_390), .C(n_392), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g398 ( .A(n_387), .Y(n_398) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_395), .B2(n_396), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_402), .B2(n_403), .C(n_404), .Y(n_399) );
NAND2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g695 ( .A(n_419), .Y(n_695) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g692 ( .A(n_421), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g703 ( .A(n_421), .Y(n_703) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx2_ASAP7_75t_L g697 ( .A(n_424), .Y(n_697) );
OR2x2_ASAP7_75t_SL g424 ( .A(n_425), .B(n_645), .Y(n_424) );
NAND5xp2_ASAP7_75t_L g425 ( .A(n_426), .B(n_557), .C(n_595), .D(n_616), .E(n_633), .Y(n_425) );
NOR3xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_529), .C(n_550), .Y(n_426) );
OAI221xp5_ASAP7_75t_SL g427 ( .A1(n_428), .A2(n_471), .B1(n_495), .B2(n_516), .C(n_520), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_441), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_430), .B(n_518), .Y(n_537) );
OR2x2_ASAP7_75t_L g564 ( .A(n_430), .B(n_454), .Y(n_564) );
AND2x2_ASAP7_75t_L g578 ( .A(n_430), .B(n_454), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_430), .B(n_444), .Y(n_592) );
AND2x2_ASAP7_75t_L g630 ( .A(n_430), .B(n_594), .Y(n_630) );
AND2x2_ASAP7_75t_L g659 ( .A(n_430), .B(n_569), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_430), .B(n_541), .Y(n_676) );
INVx4_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g556 ( .A(n_431), .B(n_453), .Y(n_556) );
BUFx3_ASAP7_75t_L g581 ( .A(n_431), .Y(n_581) );
AND2x2_ASAP7_75t_L g610 ( .A(n_431), .B(n_454), .Y(n_610) );
AND3x2_ASAP7_75t_L g623 ( .A(n_431), .B(n_624), .C(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g546 ( .A(n_441), .Y(n_546) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_453), .Y(n_441) );
AOI32xp33_ASAP7_75t_L g601 ( .A1(n_442), .A2(n_553), .A3(n_602), .B1(n_605), .B2(n_606), .Y(n_601) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g528 ( .A(n_443), .B(n_453), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_443), .B(n_556), .Y(n_599) );
AND2x2_ASAP7_75t_L g606 ( .A(n_443), .B(n_578), .Y(n_606) );
OR2x2_ASAP7_75t_L g612 ( .A(n_443), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_443), .B(n_567), .Y(n_637) );
OR2x2_ASAP7_75t_L g655 ( .A(n_443), .B(n_483), .Y(n_655) );
BUFx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g519 ( .A(n_444), .B(n_463), .Y(n_519) );
INVx2_ASAP7_75t_L g541 ( .A(n_444), .Y(n_541) );
OR2x2_ASAP7_75t_L g563 ( .A(n_444), .B(n_463), .Y(n_563) );
AND2x2_ASAP7_75t_L g568 ( .A(n_444), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_444), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g624 ( .A(n_444), .B(n_518), .Y(n_624) );
INVx1_ASAP7_75t_SL g675 ( .A(n_453), .Y(n_675) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_463), .Y(n_453) );
INVx1_ASAP7_75t_SL g518 ( .A(n_454), .Y(n_518) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_454), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_454), .B(n_604), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_454), .B(n_541), .C(n_659), .Y(n_670) );
INVx2_ASAP7_75t_L g569 ( .A(n_463), .Y(n_569) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_463), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .Y(n_471) );
INVx1_ASAP7_75t_L g605 ( .A(n_472), .Y(n_605) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g523 ( .A(n_473), .B(n_506), .Y(n_523) );
INVx2_ASAP7_75t_L g540 ( .A(n_473), .Y(n_540) );
AND2x2_ASAP7_75t_L g545 ( .A(n_473), .B(n_507), .Y(n_545) );
AND2x2_ASAP7_75t_L g560 ( .A(n_473), .B(n_496), .Y(n_560) );
AND2x2_ASAP7_75t_L g572 ( .A(n_473), .B(n_544), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_482), .B(n_588), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g644 ( .A(n_482), .B(n_545), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_482), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_482), .B(n_539), .Y(n_667) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g505 ( .A(n_483), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_483), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g549 ( .A(n_483), .B(n_496), .Y(n_549) );
AND2x2_ASAP7_75t_L g575 ( .A(n_483), .B(n_506), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_483), .B(n_615), .Y(n_614) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_487), .B(n_494), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_485), .A2(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g534 ( .A(n_487), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_494), .Y(n_535) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_505), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_496), .B(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g539 ( .A(n_496), .B(n_540), .Y(n_539) );
INVx3_ASAP7_75t_SL g544 ( .A(n_496), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_496), .B(n_531), .Y(n_597) );
OR2x2_ASAP7_75t_L g607 ( .A(n_496), .B(n_533), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_496), .B(n_575), .Y(n_635) );
OR2x2_ASAP7_75t_L g665 ( .A(n_496), .B(n_506), .Y(n_665) );
AND2x2_ASAP7_75t_L g669 ( .A(n_496), .B(n_507), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_496), .B(n_545), .Y(n_682) );
AND2x2_ASAP7_75t_L g689 ( .A(n_496), .B(n_571), .Y(n_689) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
INVx1_ASAP7_75t_SL g632 ( .A(n_505), .Y(n_632) );
AND2x2_ASAP7_75t_L g571 ( .A(n_506), .B(n_533), .Y(n_571) );
AND2x2_ASAP7_75t_L g585 ( .A(n_506), .B(n_540), .Y(n_585) );
AND2x2_ASAP7_75t_L g588 ( .A(n_506), .B(n_544), .Y(n_588) );
INVx1_ASAP7_75t_L g615 ( .A(n_506), .Y(n_615) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g527 ( .A(n_507), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_519), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g686 ( .A1(n_517), .A2(n_563), .B(n_687), .C(n_688), .Y(n_686) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g593 ( .A(n_518), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_519), .B(n_536), .Y(n_551) );
AND2x2_ASAP7_75t_L g577 ( .A(n_519), .B(n_578), .Y(n_577) );
OAI21xp5_ASAP7_75t_SL g520 ( .A1(n_521), .A2(n_524), .B(n_528), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_522), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g548 ( .A(n_523), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_523), .B(n_544), .Y(n_589) );
AND2x2_ASAP7_75t_L g680 ( .A(n_523), .B(n_531), .Y(n_680) );
INVxp67_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g553 ( .A(n_527), .B(n_540), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_527), .B(n_538), .Y(n_554) );
OAI322xp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_537), .A3(n_538), .B1(n_541), .B2(n_542), .C1(n_546), .C2(n_547), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
AND2x2_ASAP7_75t_L g641 ( .A(n_531), .B(n_553), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_531), .B(n_605), .Y(n_687) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g584 ( .A(n_533), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g650 ( .A(n_537), .B(n_563), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_538), .B(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_539), .B(n_571), .Y(n_628) );
AND2x2_ASAP7_75t_L g574 ( .A(n_540), .B(n_544), .Y(n_574) );
AND2x2_ASAP7_75t_L g582 ( .A(n_541), .B(n_583), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_541), .A2(n_620), .B(n_680), .C(n_681), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g652 ( .A1(n_542), .A2(n_555), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_544), .B(n_571), .Y(n_611) );
AND2x2_ASAP7_75t_L g617 ( .A(n_544), .B(n_585), .Y(n_617) );
AND2x2_ASAP7_75t_L g651 ( .A(n_544), .B(n_553), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_545), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_SL g661 ( .A(n_545), .Y(n_661) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_549), .A2(n_577), .B1(n_579), .B2(n_584), .Y(n_576) );
OAI22xp5_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_552), .B1(n_554), .B2(n_555), .Y(n_550) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_551), .A2(n_587), .B1(n_589), .B2(n_590), .Y(n_586) );
INVxp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_556), .A2(n_658), .B1(n_660), .B2(n_662), .C(n_666), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B(n_565), .C(n_586), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
OR2x2_ASAP7_75t_L g627 ( .A(n_563), .B(n_580), .Y(n_627) );
INVx1_ASAP7_75t_L g678 ( .A(n_563), .Y(n_678) );
OAI221xp5_ASAP7_75t_L g565 ( .A1(n_564), .A2(n_566), .B1(n_570), .B2(n_573), .C(n_576), .Y(n_565) );
INVx2_ASAP7_75t_SL g620 ( .A(n_564), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g685 ( .A(n_567), .Y(n_685) );
AND2x2_ASAP7_75t_L g609 ( .A(n_568), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g594 ( .A(n_569), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g656 ( .A(n_572), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_580), .B(n_682), .Y(n_681) );
CKINVDCx16_ASAP7_75t_R g580 ( .A(n_581), .Y(n_580) );
INVxp67_ASAP7_75t_L g625 ( .A(n_583), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g595 ( .A1(n_584), .A2(n_596), .B(n_598), .C(n_600), .Y(n_595) );
INVx1_ASAP7_75t_L g673 ( .A(n_587), .Y(n_673) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_591), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx2_ASAP7_75t_L g604 ( .A(n_594), .Y(n_604) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI222xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_607), .B1(n_608), .B2(n_611), .C1(n_612), .C2(n_614), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_SL g640 ( .A(n_604), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_607), .B(n_661), .Y(n_660) );
NAND2xp33_ASAP7_75t_SL g638 ( .A(n_608), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g613 ( .A(n_610), .Y(n_613) );
AND2x2_ASAP7_75t_L g677 ( .A(n_610), .B(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g643 ( .A(n_613), .B(n_640), .Y(n_643) );
INVx1_ASAP7_75t_L g672 ( .A(n_614), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_621), .C(n_626), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_620), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
AOI322xp5_ASAP7_75t_L g671 ( .A1(n_623), .A2(n_651), .A3(n_656), .B1(n_672), .B2(n_673), .C1(n_674), .C2(n_677), .Y(n_671) );
AND2x2_ASAP7_75t_L g658 ( .A(n_624), .B(n_659), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_629), .B2(n_631), .Y(n_626) );
INVxp33_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B1(n_638), .B2(n_641), .C(n_642), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NAND5xp2_ASAP7_75t_L g645 ( .A(n_646), .B(n_657), .C(n_671), .D(n_679), .E(n_683), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_651), .B(n_652), .Y(n_646) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVxp33_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_659), .A2(n_684), .B(n_685), .C(n_686), .Y(n_683) );
AOI31xp33_ASAP7_75t_L g666 ( .A1(n_661), .A2(n_667), .A3(n_668), .B(n_670), .Y(n_666) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g684 ( .A(n_682), .Y(n_684) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g698 ( .A(n_691), .Y(n_698) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NOR2x2_ASAP7_75t_L g702 ( .A(n_693), .B(n_703), .Y(n_702) );
OAI22x1_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_694) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_710), .Y(n_705) );
NOR2xp33_ASAP7_75t_SL g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx1_ASAP7_75t_SL g731 ( .A(n_707), .Y(n_731) );
INVx1_ASAP7_75t_L g730 ( .A(n_709), .Y(n_730) );
OA21x2_ASAP7_75t_L g733 ( .A1(n_709), .A2(n_731), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_712), .Y(n_721) );
INVx2_ASAP7_75t_L g725 ( .A(n_712), .Y(n_725) );
BUFx2_ASAP7_75t_L g734 ( .A(n_712), .Y(n_734) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_719), .B(n_722), .Y(n_714) );
INVx1_ASAP7_75t_L g718 ( .A(n_717), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
endmodule