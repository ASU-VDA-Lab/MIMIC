module fake_netlist_5_1473_n_770 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_770);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_770;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_501;
wire n_245;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_718;
wire n_671;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_443;
wire n_372;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_150;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_519;
wire n_406;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_432;
wire n_164;
wire n_553;
wire n_395;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_679;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_82),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_36),
.Y(n_150)
);

BUFx10_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_75),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_55),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_50),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_78),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_57),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_44),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_4),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_119),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_25),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_94),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_45),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_25),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_16),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_72),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_39),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_35),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_70),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_37),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_115),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_65),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_18),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_69),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_60),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_61),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_24),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_47),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_0),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_52),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_21),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_97),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_141),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_13),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_14),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_96),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_77),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_16),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_139),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_62),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_19),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_144),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_183),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_152),
.B(n_26),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_151),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

BUFx8_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_151),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_0),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_27),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_157),
.B(n_197),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_1),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_147),
.B(n_1),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_154),
.B(n_161),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_164),
.B(n_2),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_151),
.B(n_2),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_3),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_3),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_4),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_5),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_160),
.B(n_167),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_169),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_158),
.B(n_5),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_6),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_176),
.B1(n_153),
.B2(n_155),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_223),
.B(n_210),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g242 ( 
.A(n_223),
.B(n_153),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_176),
.B1(n_155),
.B2(n_195),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_216),
.A2(n_226),
.B1(n_208),
.B2(n_201),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_226),
.A2(n_208),
.B1(n_201),
.B2(n_220),
.Y(n_245)
);

OR2x6_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_150),
.Y(n_246)
);

NAND3x1_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_225),
.C(n_222),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_189),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_201),
.A2(n_185),
.B1(n_179),
.B2(n_168),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_198),
.B1(n_187),
.B2(n_194),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_202),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_189),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_190),
.B1(n_194),
.B2(n_184),
.Y(n_254)
);

AO22x2_ASAP7_75t_L g255 ( 
.A1(n_201),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_202),
.B(n_190),
.Y(n_257)
);

AO22x2_ASAP7_75t_L g258 ( 
.A1(n_208),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_174),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_196),
.B1(n_186),
.B2(n_182),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_180),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_207),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_204),
.B(n_175),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_208),
.B(n_28),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_206),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_209),
.B(n_29),
.Y(n_268)
);

AO22x2_ASAP7_75t_L g269 ( 
.A1(n_217),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_230),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_215),
.B(n_12),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_207),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_234),
.Y(n_274)
);

AO22x2_ASAP7_75t_L g275 ( 
.A1(n_217),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_211),
.B(n_231),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_200),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_236),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_215),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_200),
.B(n_212),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_207),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_200),
.B(n_30),
.Y(n_282)
);

INVx8_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_235),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_212),
.B(n_31),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_212),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_266),
.B(n_217),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_235),
.Y(n_290)
);

AND2x4_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_217),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_250),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_240),
.B(n_238),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_262),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

XNOR2x2_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_22),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_205),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_268),
.Y(n_306)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_265),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_248),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_253),
.Y(n_314)
);

NAND2x1p5_ASAP7_75t_L g315 ( 
.A(n_241),
.B(n_228),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_224),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_261),
.Y(n_317)
);

INVx4_ASAP7_75t_SL g318 ( 
.A(n_246),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_261),
.Y(n_319)
);

INVx4_ASAP7_75t_SL g320 ( 
.A(n_246),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

XNOR2x2_ASAP7_75t_L g322 ( 
.A(n_258),
.B(n_23),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_257),
.B(n_235),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_269),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_254),
.B(n_237),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

INVx4_ASAP7_75t_SL g327 ( 
.A(n_246),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_275),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_260),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_275),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_R g331 ( 
.A(n_267),
.B(n_24),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_275),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

BUFx6f_ASAP7_75t_SL g334 ( 
.A(n_283),
.Y(n_334)
);

AND2x6_ASAP7_75t_L g335 ( 
.A(n_278),
.B(n_209),
.Y(n_335)
);

NAND2x1p5_ASAP7_75t_L g336 ( 
.A(n_272),
.B(n_199),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_245),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_245),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_244),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_249),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_283),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_249),
.B(n_237),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_244),
.B(n_214),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_271),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_255),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_283),
.B(n_237),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_276),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_242),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_255),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_255),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_287),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_329),
.B(n_271),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_209),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_298),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_214),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_303),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_305),
.B(n_284),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_333),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_308),
.B(n_214),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_298),
.B(n_251),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_316),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_286),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_289),
.B(n_339),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_214),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_214),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_348),
.Y(n_366)
);

AND2x2_ASAP7_75t_SL g367 ( 
.A(n_313),
.B(n_279),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_291),
.B(n_214),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_343),
.A2(n_199),
.B(n_224),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_32),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_300),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_211),
.B(n_199),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_291),
.B(n_203),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_304),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_302),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_312),
.B(n_314),
.Y(n_379)
);

AND2x2_ASAP7_75t_SL g380 ( 
.A(n_313),
.B(n_224),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_292),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_311),
.B(n_199),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_297),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_315),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_299),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_290),
.B(n_203),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_315),
.B(n_224),
.Y(n_388)
);

INVx6_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_309),
.B(n_224),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_321),
.B(n_324),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_310),
.B(n_224),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_293),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_301),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_295),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_296),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_328),
.B(n_229),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_203),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_330),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_332),
.B(n_345),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_349),
.Y(n_404)
);

AND2x2_ASAP7_75t_SL g405 ( 
.A(n_342),
.B(n_229),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_336),
.B(n_229),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_335),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_SL g408 ( 
.A(n_294),
.B(n_229),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_340),
.B(n_203),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_335),
.B(n_213),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_290),
.B(n_213),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_322),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_318),
.B(n_33),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_323),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_362),
.B(n_318),
.Y(n_417)
);

CKINVDCx6p67_ASAP7_75t_R g418 ( 
.A(n_354),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_353),
.B(n_323),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_353),
.B(n_325),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_307),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_354),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_346),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_382),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_378),
.B(n_366),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_382),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_378),
.B(n_341),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_382),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_362),
.B(n_318),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_382),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_358),
.B(n_334),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_397),
.Y(n_434)
);

BUFx8_ASAP7_75t_SL g435 ( 
.A(n_396),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_362),
.B(n_320),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_397),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_370),
.B(n_213),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_390),
.B(n_320),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_376),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_361),
.B(n_213),
.Y(n_441)
);

BUFx4f_ASAP7_75t_L g442 ( 
.A(n_415),
.Y(n_442)
);

CKINVDCx6p67_ASAP7_75t_R g443 ( 
.A(n_367),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_408),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_320),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_360),
.B(n_229),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_361),
.B(n_327),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_407),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_403),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_379),
.B(n_327),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_379),
.B(n_327),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_356),
.Y(n_453)
);

OR2x6_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_334),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_403),
.B(n_211),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_360),
.B(n_229),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_383),
.B(n_211),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_376),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_371),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_413),
.B(n_211),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_416),
.B(n_211),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_356),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_376),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_415),
.B(n_34),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_416),
.B(n_385),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_397),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_356),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_383),
.B(n_38),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_413),
.B(n_396),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_403),
.B(n_40),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_422),
.Y(n_473)
);

INVx3_ASAP7_75t_SL g474 ( 
.A(n_418),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_453),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

BUFx2_ASAP7_75t_SL g477 ( 
.A(n_445),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_385),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_471),
.Y(n_479)
);

NAND2x1p5_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_393),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_463),
.Y(n_481)
);

CKINVDCx11_ASAP7_75t_R g482 ( 
.A(n_454),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_434),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_425),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_452),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_375),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_443),
.A2(n_393),
.B1(n_409),
.B2(n_367),
.Y(n_487)
);

INVx3_ASAP7_75t_SL g488 ( 
.A(n_454),
.Y(n_488)
);

BUFx12f_ASAP7_75t_L g489 ( 
.A(n_454),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_419),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_425),
.Y(n_491)
);

BUFx12f_ASAP7_75t_L g492 ( 
.A(n_445),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_425),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_437),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_425),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_417),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_421),
.B(n_404),
.Y(n_498)
);

BUFx4_ASAP7_75t_SL g499 ( 
.A(n_444),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_420),
.B(n_404),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_446),
.B(n_413),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_435),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_467),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_393),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_430),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_423),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_435),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_430),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_430),
.Y(n_509)
);

BUFx2_ASAP7_75t_R g510 ( 
.A(n_444),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_459),
.Y(n_511)
);

INVx3_ASAP7_75t_SL g512 ( 
.A(n_417),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_450),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_451),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_452),
.B(n_404),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

INVx6_ASAP7_75t_L g517 ( 
.A(n_417),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_470),
.Y(n_518)
);

BUFx8_ASAP7_75t_L g519 ( 
.A(n_431),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_465),
.A2(n_352),
.B1(n_405),
.B2(n_367),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_474),
.Y(n_521)
);

INVx6_ASAP7_75t_L g522 ( 
.A(n_519),
.Y(n_522)
);

OAI22xp33_ASAP7_75t_L g523 ( 
.A1(n_501),
.A2(n_352),
.B1(n_461),
.B2(n_416),
.Y(n_523)
);

INVx6_ASAP7_75t_L g524 ( 
.A(n_519),
.Y(n_524)
);

BUFx12f_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

AOI21xp33_ASAP7_75t_SL g526 ( 
.A1(n_474),
.A2(n_429),
.B(n_426),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_492),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_520),
.A2(n_460),
.B1(n_452),
.B2(n_464),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_475),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_479),
.Y(n_530)
);

INVx6_ASAP7_75t_L g531 ( 
.A(n_517),
.Y(n_531)
);

CKINVDCx11_ASAP7_75t_R g532 ( 
.A(n_482),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_520),
.A2(n_429),
.B(n_426),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_490),
.A2(n_460),
.B1(n_440),
.B2(n_464),
.Y(n_534)
);

BUFx4f_ASAP7_75t_SL g535 ( 
.A(n_489),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_476),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_499),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_518),
.A2(n_357),
.B1(n_405),
.B2(n_514),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_SL g539 ( 
.A1(n_490),
.A2(n_405),
.B1(n_465),
.B2(n_380),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_511),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_478),
.A2(n_460),
.B1(n_440),
.B2(n_389),
.Y(n_541)
);

INVx3_ASAP7_75t_SL g542 ( 
.A(n_488),
.Y(n_542)
);

AO22x1_ASAP7_75t_L g543 ( 
.A1(n_502),
.A2(n_439),
.B1(n_412),
.B2(n_465),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_483),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_481),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_494),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_478),
.A2(n_460),
.B1(n_389),
.B2(n_403),
.Y(n_547)
);

CKINVDCx11_ASAP7_75t_R g548 ( 
.A(n_507),
.Y(n_548)
);

OAI22xp33_ASAP7_75t_L g549 ( 
.A1(n_487),
.A2(n_456),
.B1(n_375),
.B2(n_412),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_503),
.Y(n_550)
);

CKINVDCx11_ASAP7_75t_R g551 ( 
.A(n_488),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_513),
.A2(n_357),
.B(n_387),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_506),
.A2(n_433),
.B1(n_375),
.B2(n_441),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_498),
.Y(n_554)
);

CKINVDCx11_ASAP7_75t_R g555 ( 
.A(n_473),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_499),
.Y(n_556)
);

BUFx4f_ASAP7_75t_L g557 ( 
.A(n_512),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_486),
.A2(n_357),
.B1(n_448),
.B2(n_458),
.Y(n_558)
);

CKINVDCx11_ASAP7_75t_R g559 ( 
.A(n_512),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_517),
.Y(n_560)
);

NAND2x1p5_ASAP7_75t_L g561 ( 
.A(n_505),
.B(n_431),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_554),
.B(n_498),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_555),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_539),
.A2(n_439),
.B1(n_389),
.B2(n_486),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_539),
.A2(n_533),
.B1(n_538),
.B2(n_558),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_523),
.B(n_500),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_540),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_552),
.A2(n_447),
.B1(n_357),
.B2(n_410),
.Y(n_568)
);

OAI222xp33_ASAP7_75t_L g569 ( 
.A1(n_523),
.A2(n_500),
.B1(n_515),
.B2(n_363),
.C1(n_410),
.C2(n_480),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_540),
.B(n_350),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_526),
.A2(n_389),
.B1(n_447),
.B2(n_480),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_537),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_553),
.A2(n_389),
.B1(n_504),
.B2(n_380),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_546),
.B(n_529),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_543),
.A2(n_469),
.B1(n_374),
.B2(n_400),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_556),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_531),
.B(n_510),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_536),
.B(n_545),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_530),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_549),
.A2(n_363),
.B1(n_384),
.B2(n_386),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_549),
.A2(n_386),
.B1(n_384),
.B2(n_438),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_551),
.A2(n_386),
.B1(n_414),
.B2(n_394),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_522),
.A2(n_380),
.B1(n_350),
.B2(n_504),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_528),
.B(n_400),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_544),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_550),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_534),
.B(n_391),
.C(n_394),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_522),
.A2(n_373),
.B1(n_462),
.B2(n_436),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_525),
.A2(n_414),
.B1(n_391),
.B2(n_398),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_561),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_521),
.A2(n_374),
.B1(n_431),
.B2(n_436),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_560),
.B(n_401),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_561),
.Y(n_593)
);

OAI21xp33_ASAP7_75t_L g594 ( 
.A1(n_541),
.A2(n_510),
.B(n_515),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_547),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_531),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_531),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_557),
.A2(n_517),
.B1(n_497),
.B2(n_477),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_557),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_559),
.A2(n_414),
.B1(n_398),
.B2(n_497),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_527),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_535),
.A2(n_388),
.B1(n_406),
.B2(n_485),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_542),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_522),
.A2(n_388),
.B1(n_406),
.B2(n_485),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_548),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_542),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_532),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_L g608 ( 
.A(n_524),
.B(n_516),
.C(n_472),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_524),
.A2(n_527),
.B1(n_399),
.B2(n_516),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_565),
.A2(n_524),
.B1(n_527),
.B2(n_436),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_600),
.A2(n_462),
.B1(n_449),
.B2(n_432),
.Y(n_611)
);

OAI211xp5_ASAP7_75t_L g612 ( 
.A1(n_575),
.A2(n_401),
.B(n_402),
.C(n_373),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_574),
.B(n_364),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_594),
.A2(n_377),
.B1(n_372),
.B2(n_399),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_583),
.A2(n_509),
.B1(n_505),
.B2(n_392),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_574),
.B(n_364),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_589),
.A2(n_427),
.B1(n_395),
.B2(n_505),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_584),
.A2(n_587),
.B(n_569),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_567),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_562),
.B(n_365),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_584),
.A2(n_372),
.B1(n_377),
.B2(n_365),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_566),
.A2(n_371),
.B1(n_509),
.B2(n_505),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_568),
.A2(n_372),
.B1(n_377),
.B2(n_368),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_608),
.A2(n_368),
.B1(n_371),
.B2(n_395),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_578),
.B(n_369),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_SL g626 ( 
.A1(n_564),
.A2(n_509),
.B1(n_491),
.B2(n_495),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_603),
.A2(n_606),
.B1(n_591),
.B2(n_582),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_585),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_573),
.A2(n_509),
.B1(n_491),
.B2(n_495),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_578),
.B(n_369),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_603),
.A2(n_424),
.B1(n_428),
.B2(n_381),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_606),
.A2(n_424),
.B1(n_428),
.B2(n_381),
.Y(n_632)
);

OAI221xp5_ASAP7_75t_L g633 ( 
.A1(n_609),
.A2(n_588),
.B1(n_602),
.B2(n_604),
.C(n_581),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_595),
.A2(n_381),
.B1(n_457),
.B2(n_359),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_599),
.A2(n_381),
.B1(n_355),
.B2(n_359),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_570),
.A2(n_392),
.B1(n_355),
.B2(n_468),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_596),
.A2(n_351),
.B1(n_468),
.B2(n_463),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_585),
.B(n_579),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_597),
.A2(n_351),
.B1(n_496),
.B2(n_484),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_586),
.B(n_592),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_577),
.A2(n_351),
.B1(n_496),
.B2(n_484),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_571),
.A2(n_351),
.B1(n_508),
.B2(n_493),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_563),
.A2(n_508),
.B1(n_493),
.B2(n_495),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_572),
.B(n_392),
.Y(n_644)
);

OAI221xp5_ASAP7_75t_L g645 ( 
.A1(n_580),
.A2(n_402),
.B1(n_455),
.B2(n_491),
.C(n_495),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_601),
.A2(n_392),
.B1(n_491),
.B2(n_43),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_628),
.B(n_590),
.Y(n_647)
);

NAND3xp33_ASAP7_75t_L g648 ( 
.A(n_627),
.B(n_598),
.C(n_601),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_619),
.B(n_590),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_618),
.B(n_601),
.C(n_593),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_619),
.B(n_593),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_610),
.A2(n_601),
.B1(n_605),
.B2(n_607),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_633),
.A2(n_605),
.B1(n_607),
.B2(n_576),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_640),
.B(n_572),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_638),
.B(n_628),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_618),
.A2(n_626),
.B1(n_646),
.B2(n_645),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_646),
.A2(n_576),
.B1(n_42),
.B2(n_46),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_629),
.B(n_625),
.Y(n_658)
);

OA21x2_ASAP7_75t_L g659 ( 
.A1(n_612),
.A2(n_41),
.B(n_48),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_630),
.B(n_49),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_613),
.B(n_51),
.Y(n_661)
);

AND4x1_ASAP7_75t_L g662 ( 
.A(n_643),
.B(n_641),
.C(n_624),
.D(n_644),
.Y(n_662)
);

OAI21xp33_ASAP7_75t_L g663 ( 
.A1(n_614),
.A2(n_53),
.B(n_54),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_636),
.B(n_56),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_636),
.B(n_58),
.C(n_63),
.Y(n_665)
);

OAI221xp5_ASAP7_75t_SL g666 ( 
.A1(n_622),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.C(n_68),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_616),
.B(n_71),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_615),
.B(n_73),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_L g669 ( 
.A(n_617),
.B(n_74),
.C(n_76),
.Y(n_669)
);

OAI221xp5_ASAP7_75t_L g670 ( 
.A1(n_615),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.C(n_83),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_642),
.B(n_84),
.C(n_85),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_620),
.B(n_87),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_634),
.B(n_88),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_611),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_623),
.A2(n_92),
.B(n_93),
.Y(n_675)
);

OAI211xp5_ASAP7_75t_L g676 ( 
.A1(n_631),
.A2(n_95),
.B(n_98),
.C(n_99),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_621),
.B(n_100),
.Y(n_677)
);

AO21x2_ASAP7_75t_L g678 ( 
.A1(n_650),
.A2(n_651),
.B(n_649),
.Y(n_678)
);

NAND4xp75_ASAP7_75t_L g679 ( 
.A(n_659),
.B(n_101),
.C(n_102),
.D(n_103),
.Y(n_679)
);

NAND4xp25_ASAP7_75t_L g680 ( 
.A(n_656),
.B(n_653),
.C(n_663),
.D(n_654),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_SL g681 ( 
.A(n_648),
.B(n_639),
.C(n_632),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_647),
.B(n_635),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_655),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_647),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_658),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_658),
.B(n_637),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_659),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_672),
.B(n_142),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_664),
.B(n_104),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_659),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_664),
.B(n_105),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_668),
.B(n_110),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_660),
.B(n_111),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_L g694 ( 
.A(n_685),
.B(n_665),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_684),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_684),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_683),
.Y(n_697)
);

NAND4xp75_ASAP7_75t_L g698 ( 
.A(n_689),
.B(n_668),
.C(n_673),
.D(n_660),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_683),
.Y(n_699)
);

XNOR2xp5_ASAP7_75t_L g700 ( 
.A(n_680),
.B(n_652),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_682),
.B(n_667),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_678),
.B(n_673),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_678),
.Y(n_703)
);

XOR2x2_ASAP7_75t_L g704 ( 
.A(n_700),
.B(n_662),
.Y(n_704)
);

XNOR2x1_ASAP7_75t_L g705 ( 
.A(n_700),
.B(n_691),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_701),
.B(n_678),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_702),
.B(n_682),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_702),
.B(n_686),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_704),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_707),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_708),
.Y(n_711)
);

XNOR2x1_ASAP7_75t_L g712 ( 
.A(n_705),
.B(n_698),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_706),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_704),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_709),
.A2(n_680),
.B1(n_694),
.B2(n_692),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_711),
.Y(n_716)
);

OAI322xp33_ASAP7_75t_L g717 ( 
.A1(n_712),
.A2(n_703),
.A3(n_699),
.B1(n_697),
.B2(n_687),
.C1(n_690),
.C2(n_696),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_709),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_711),
.Y(n_719)
);

AND4x1_ASAP7_75t_L g720 ( 
.A(n_715),
.B(n_714),
.C(n_709),
.D(n_657),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_716),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_719),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_SL g723 ( 
.A1(n_721),
.A2(n_709),
.B(n_714),
.C(n_718),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_722),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_720),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_721),
.A2(n_712),
.B1(n_714),
.B2(n_710),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_724),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_725),
.B(n_714),
.Y(n_728)
);

NOR2x1_ASAP7_75t_L g729 ( 
.A(n_726),
.B(n_717),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_723),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_726),
.B(n_710),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_726),
.A2(n_713),
.B1(n_692),
.B2(n_679),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_727),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_729),
.A2(n_713),
.B1(n_692),
.B2(n_679),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_728),
.A2(n_692),
.B1(n_691),
.B2(n_689),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_732),
.A2(n_730),
.B1(n_731),
.B2(n_688),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_730),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_730),
.Y(n_738)
);

NOR2xp67_ASAP7_75t_L g739 ( 
.A(n_730),
.B(n_696),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_734),
.A2(n_693),
.B1(n_687),
.B2(n_686),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_736),
.A2(n_687),
.B1(n_695),
.B2(n_690),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_737),
.A2(n_693),
.B1(n_675),
.B2(n_663),
.Y(n_742)
);

OAI211xp5_ASAP7_75t_L g743 ( 
.A1(n_738),
.A2(n_674),
.B(n_670),
.C(n_666),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_739),
.A2(n_681),
.B1(n_661),
.B2(n_669),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_733),
.A2(n_671),
.B1(n_676),
.B2(n_677),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_735),
.Y(n_746)
);

AND4x1_ASAP7_75t_L g747 ( 
.A(n_734),
.B(n_662),
.C(n_113),
.D(n_114),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_737),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_748),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_746),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_740),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_744),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_747),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_742),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_745),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_741),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_750),
.A2(n_743),
.B1(n_121),
.B2(n_123),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_749),
.A2(n_120),
.B1(n_124),
.B2(n_125),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_751),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_753),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_754),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_761)
);

INVxp67_ASAP7_75t_SL g762 ( 
.A(n_760),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_759),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_762),
.A2(n_755),
.B1(n_756),
.B2(n_757),
.Y(n_764)
);

AOI31xp33_ASAP7_75t_L g765 ( 
.A1(n_763),
.A2(n_756),
.A3(n_752),
.B(n_761),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_765),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_L g767 ( 
.A1(n_766),
.A2(n_758),
.B1(n_764),
.B2(n_131),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_767),
.Y(n_768)
);

AOI221xp5_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.C(n_135),
.Y(n_769)
);

AOI211xp5_ASAP7_75t_L g770 ( 
.A1(n_769),
.A2(n_136),
.B(n_137),
.C(n_138),
.Y(n_770)
);


endmodule