module fake_netlist_6_1446_n_1013 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1013);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1013;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_720;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_940;
wire n_770;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_886;
wire n_1004;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_217;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_262;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_956;
wire n_841;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_133),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_171),
.Y(n_215)
);

INVxp33_ASAP7_75t_SL g216 ( 
.A(n_124),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_140),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_42),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_138),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_13),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_185),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_105),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_136),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_77),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_47),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_95),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_92),
.Y(n_229)
);

BUFx8_ASAP7_75t_SL g230 ( 
.A(n_127),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_189),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_45),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_204),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_192),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_26),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_74),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_18),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_102),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_169),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_165),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_134),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_120),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_106),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_205),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_180),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_18),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_132),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_43),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_198),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_14),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_16),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_206),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_79),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_25),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_10),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_178),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_72),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_210),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_82),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_30),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_110),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_139),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_150),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_93),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_119),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_55),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_104),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_62),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_142),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_144),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_17),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_80),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_23),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_187),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_69),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_114),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_125),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_158),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_89),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_85),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_61),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_51),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_76),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_174),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_31),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_108),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_181),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_57),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_160),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_67),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_145),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_195),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_149),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_121),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_137),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_12),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_9),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_162),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_301),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_252),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_222),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_225),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_237),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_263),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_275),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_302),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_0),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_230),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_252),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_215),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_254),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_216),
.B(n_0),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_256),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_252),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_252),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_258),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_219),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_277),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_289),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_246),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_220),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_223),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_246),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_254),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_230),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_288),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_288),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_299),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_218),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_299),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_213),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_287),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_221),
.B(n_1),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_297),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_214),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_233),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_240),
.Y(n_348)
);

INVxp33_ASAP7_75t_L g349 ( 
.A(n_242),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_221),
.B(n_226),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_294),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_224),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_227),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_251),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_298),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_267),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_306),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_322),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_315),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_323),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_308),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_326),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_317),
.B(n_226),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_324),
.B(n_282),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_342),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_315),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_332),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_332),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_331),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_305),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_320),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_328),
.B(n_282),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_307),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_347),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_329),
.B(n_303),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_343),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_350),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_327),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_318),
.B(n_228),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

NAND2xp33_ASAP7_75t_L g398 ( 
.A(n_309),
.B(n_229),
.Y(n_398)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_340),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_313),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_345),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_267),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_314),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_353),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_309),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_353),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_354),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_354),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_310),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_310),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_330),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_335),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_311),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_311),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_337),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_312),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_402),
.Y(n_417)
);

BUFx4f_ASAP7_75t_L g418 ( 
.A(n_399),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_393),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_365),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_383),
.Y(n_422)
);

AND2x6_ASAP7_75t_L g423 ( 
.A(n_397),
.B(n_229),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_400),
.B(n_312),
.C(n_357),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_378),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_379),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_371),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_358),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_397),
.B(n_217),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_R g435 ( 
.A(n_362),
.B(n_335),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_236),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_359),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_375),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_382),
.B(n_339),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_R g441 ( 
.A(n_362),
.B(n_339),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_375),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_397),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_392),
.B(n_270),
.Y(n_444)
);

INVx8_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_360),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_392),
.B(n_272),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_388),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_380),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_387),
.B(n_276),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_367),
.B(n_231),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_377),
.B(n_229),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_402),
.Y(n_453)
);

INVx4_ASAP7_75t_SL g454 ( 
.A(n_399),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_395),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_363),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_361),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_371),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_364),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_376),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_368),
.B(n_232),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_381),
.B(n_234),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_413),
.A2(n_266),
.B1(n_300),
.B2(n_296),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_377),
.Y(n_466)
);

AND2x6_ASAP7_75t_L g467 ( 
.A(n_404),
.B(n_229),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_364),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_376),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_394),
.B(n_403),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_394),
.A2(n_273),
.B1(n_235),
.B2(n_267),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_412),
.Y(n_472)
);

INVx6_ASAP7_75t_L g473 ( 
.A(n_399),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_377),
.B(n_273),
.Y(n_474)
);

AO22x2_ASAP7_75t_L g475 ( 
.A1(n_413),
.A2(n_235),
.B1(n_2),
.B2(n_3),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_366),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_366),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_410),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_410),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_404),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_414),
.B(n_273),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_414),
.A2(n_273),
.B1(n_281),
.B2(n_293),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_406),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_406),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_398),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_405),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_389),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_391),
.B(n_341),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_409),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_396),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_480),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_480),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_407),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_480),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_488),
.A2(n_417),
.B1(n_453),
.B2(n_455),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_443),
.A2(n_239),
.B(n_238),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_443),
.B(n_407),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_443),
.B(n_444),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_440),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_480),
.B(n_408),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_444),
.B(n_408),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_416),
.A2(n_341),
.B1(n_241),
.B2(n_274),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_483),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_434),
.B(n_437),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_489),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_463),
.B(n_396),
.Y(n_508)
);

A2O1A1Ixp33_ASAP7_75t_L g509 ( 
.A1(n_463),
.A2(n_243),
.B(n_244),
.C(n_245),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_427),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_429),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_430),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_464),
.B(n_248),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_464),
.B(n_249),
.Y(n_514)
);

NOR3xp33_ASAP7_75t_L g515 ( 
.A(n_483),
.B(n_412),
.C(n_411),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_250),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_421),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_427),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_477),
.B(n_253),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_470),
.B(n_390),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_370),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_481),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_433),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_481),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_484),
.B(n_373),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_427),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_477),
.B(n_484),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_471),
.B(n_373),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_471),
.B(n_374),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_421),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_484),
.B(n_374),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_447),
.B(n_255),
.Y(n_532)
);

AND2x4_ASAP7_75t_SL g533 ( 
.A(n_485),
.B(n_281),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_478),
.B(n_259),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_422),
.Y(n_535)
);

NOR2xp67_ASAP7_75t_L g536 ( 
.A(n_485),
.B(n_390),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_449),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_485),
.B(n_260),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_486),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_418),
.B(n_262),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_487),
.B(n_268),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_479),
.B(n_269),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_457),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_487),
.B(n_271),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_482),
.A2(n_281),
.B1(n_278),
.B2(n_284),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_424),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_418),
.B(n_280),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_482),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_548)
);

A2O1A1Ixp33_ASAP7_75t_L g549 ( 
.A1(n_436),
.A2(n_283),
.B(n_295),
.C(n_401),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_451),
.B(n_1),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_439),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_481),
.B(n_40),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_475),
.A2(n_401),
.B1(n_386),
.B2(n_415),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_445),
.B(n_386),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_466),
.B(n_41),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_466),
.B(n_44),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_459),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_466),
.B(n_46),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_449),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_450),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_442),
.B(n_48),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_450),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_491),
.B(n_4),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_456),
.B(n_49),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_460),
.B(n_50),
.Y(n_565)
);

AO22x1_ASAP7_75t_L g566 ( 
.A1(n_491),
.A2(n_492),
.B1(n_450),
.B2(n_490),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_492),
.B(n_5),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_461),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_468),
.B(n_52),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_476),
.B(n_53),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_459),
.B(n_54),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_472),
.B(n_5),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_459),
.B(n_58),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_425),
.A2(n_103),
.B1(n_212),
.B2(n_209),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_459),
.B(n_59),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_422),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_426),
.Y(n_577)
);

A2O1A1Ixp33_ASAP7_75t_L g578 ( 
.A1(n_469),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_SL g579 ( 
.A(n_503),
.B(n_441),
.C(n_435),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_530),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_494),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_535),
.B(n_454),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_520),
.B(n_473),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_505),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_505),
.Y(n_585)
);

AND3x1_ASAP7_75t_SL g586 ( 
.A(n_559),
.B(n_475),
.C(n_441),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_510),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_511),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_506),
.B(n_469),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_SL g590 ( 
.A(n_508),
.B(n_435),
.C(n_420),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_495),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_494),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_512),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_493),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_500),
.B(n_419),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_560),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_535),
.B(n_576),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_545),
.B(n_465),
.C(n_448),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_518),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_501),
.B(n_562),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_535),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_535),
.B(n_454),
.Y(n_602)
);

INVx6_ASAP7_75t_L g603 ( 
.A(n_554),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_543),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_513),
.B(n_462),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_517),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_521),
.B(n_419),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_537),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_554),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_SL g610 ( 
.A(n_528),
.B(n_475),
.C(n_445),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_SL g611 ( 
.A(n_499),
.B(n_428),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_577),
.B(n_454),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_523),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_522),
.Y(n_614)
);

CKINVDCx16_ASAP7_75t_R g615 ( 
.A(n_554),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_507),
.B(n_431),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_521),
.B(n_419),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_550),
.A2(n_419),
.B1(n_428),
.B2(n_432),
.Y(n_618)
);

BUFx4f_ASAP7_75t_L g619 ( 
.A(n_572),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_R g620 ( 
.A(n_525),
.B(n_445),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_563),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_497),
.B(n_473),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_551),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_527),
.A2(n_423),
.B(n_432),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_514),
.B(n_525),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_550),
.A2(n_448),
.B1(n_431),
.B2(n_446),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_568),
.B(n_438),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_526),
.Y(n_628)
);

INVx6_ASAP7_75t_L g629 ( 
.A(n_493),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_SL g630 ( 
.A(n_529),
.B(n_504),
.C(n_502),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_496),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_502),
.B(n_438),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_496),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_SL g634 ( 
.A(n_545),
.B(n_446),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_531),
.B(n_473),
.Y(n_635)
);

AND2x2_ASAP7_75t_SL g636 ( 
.A(n_553),
.B(n_452),
.Y(n_636)
);

NOR3xp33_ASAP7_75t_SL g637 ( 
.A(n_549),
.B(n_6),
.C(n_7),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_524),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_R g639 ( 
.A(n_531),
.B(n_462),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_L g640 ( 
.A(n_546),
.B(n_458),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_557),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_561),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_552),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_557),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_567),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_541),
.Y(n_646)
);

OAI21xp33_ASAP7_75t_L g647 ( 
.A1(n_645),
.A2(n_591),
.B(n_548),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_625),
.B(n_567),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_624),
.A2(n_556),
.B(n_555),
.Y(n_649)
);

CKINVDCx11_ASAP7_75t_R g650 ( 
.A(n_606),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_589),
.A2(n_605),
.B(n_594),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_594),
.A2(n_558),
.B(n_538),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_631),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_581),
.A2(n_592),
.B(n_595),
.Y(n_654)
);

CKINVDCx6p67_ASAP7_75t_R g655 ( 
.A(n_580),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_619),
.A2(n_548),
.B1(n_536),
.B2(n_516),
.Y(n_656)
);

NAND2x1_ASAP7_75t_L g657 ( 
.A(n_629),
.B(n_594),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_604),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_581),
.A2(n_573),
.B(n_571),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_582),
.Y(n_660)
);

A2O1A1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_630),
.A2(n_544),
.B(n_541),
.C(n_515),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_584),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_607),
.A2(n_575),
.B(n_519),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_598),
.A2(n_634),
.B(n_643),
.C(n_640),
.Y(n_664)
);

OA22x2_ASAP7_75t_L g665 ( 
.A1(n_586),
.A2(n_553),
.B1(n_533),
.B2(n_544),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_634),
.A2(n_515),
.B(n_509),
.C(n_532),
.Y(n_666)
);

OA22x2_ASAP7_75t_L g667 ( 
.A1(n_600),
.A2(n_574),
.B1(n_566),
.B2(n_539),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_607),
.A2(n_565),
.B(n_564),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_581),
.A2(n_570),
.B(n_569),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_585),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_580),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_616),
.B(n_534),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_SL g673 ( 
.A(n_620),
.B(n_578),
.C(n_542),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_588),
.Y(n_674)
);

BUFx8_ASAP7_75t_SL g675 ( 
.A(n_606),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_617),
.A2(n_547),
.B(n_540),
.Y(n_676)
);

BUFx2_ASAP7_75t_SL g677 ( 
.A(n_583),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_L g678 ( 
.A(n_626),
.B(n_498),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_593),
.Y(n_679)
);

AOI211x1_ASAP7_75t_L g680 ( 
.A1(n_613),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_617),
.A2(n_474),
.B(n_452),
.Y(n_681)
);

AO31x2_ASAP7_75t_L g682 ( 
.A1(n_587),
.A2(n_628),
.A3(n_599),
.B(n_641),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_635),
.B(n_462),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_619),
.B(n_458),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_620),
.B(n_597),
.Y(n_685)
);

INVx4_ASAP7_75t_SL g686 ( 
.A(n_603),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_601),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_595),
.A2(n_423),
.B(n_452),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_592),
.A2(n_599),
.B(n_587),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_623),
.Y(n_690)
);

OAI21x1_ASAP7_75t_L g691 ( 
.A1(n_592),
.A2(n_423),
.B(n_467),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_616),
.B(n_474),
.Y(n_692)
);

AOI21x1_ASAP7_75t_L g693 ( 
.A1(n_628),
.A2(n_474),
.B(n_423),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_601),
.B(n_423),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_618),
.A2(n_467),
.B(n_111),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_636),
.A2(n_467),
.B1(n_112),
.B2(n_113),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_608),
.B(n_11),
.Y(n_697)
);

AO31x2_ASAP7_75t_L g698 ( 
.A1(n_641),
.A2(n_467),
.A3(n_12),
.B(n_13),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_627),
.Y(n_699)
);

AOI21x1_ASAP7_75t_L g700 ( 
.A1(n_644),
.A2(n_109),
.B(n_208),
.Y(n_700)
);

OAI21xp33_ASAP7_75t_L g701 ( 
.A1(n_610),
.A2(n_11),
.B(n_14),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_631),
.A2(n_115),
.B(n_202),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_582),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_597),
.B(n_60),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_682),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_660),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_672),
.B(n_579),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_682),
.Y(n_708)
);

BUFx5_ASAP7_75t_L g709 ( 
.A(n_699),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_689),
.A2(n_632),
.B(n_644),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_674),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_701),
.A2(n_636),
.B1(n_621),
.B2(n_590),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_659),
.A2(n_638),
.B(n_622),
.Y(n_713)
);

OAI21x1_ASAP7_75t_L g714 ( 
.A1(n_654),
.A2(n_638),
.B(n_611),
.Y(n_714)
);

OAI21x1_ASAP7_75t_L g715 ( 
.A1(n_652),
.A2(n_669),
.B(n_663),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_648),
.B(n_646),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_647),
.B(n_684),
.Y(n_717)
);

AO31x2_ASAP7_75t_L g718 ( 
.A1(n_664),
.A2(n_611),
.A3(n_637),
.B(n_639),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_R g719 ( 
.A1(n_665),
.A2(n_615),
.B1(n_603),
.B2(n_609),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_693),
.A2(n_596),
.B(n_642),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_679),
.Y(n_721)
);

AOI221xp5_ASAP7_75t_L g722 ( 
.A1(n_647),
.A2(n_627),
.B1(n_609),
.B2(n_614),
.C(n_597),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_692),
.B(n_627),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_687),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_661),
.A2(n_651),
.B(n_666),
.Y(n_725)
);

INVx8_ASAP7_75t_L g726 ( 
.A(n_687),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_695),
.A2(n_642),
.B(n_639),
.Y(n_727)
);

AO21x2_ASAP7_75t_L g728 ( 
.A1(n_649),
.A2(n_582),
.B(n_602),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_690),
.Y(n_729)
);

AO21x2_ASAP7_75t_L g730 ( 
.A1(n_649),
.A2(n_602),
.B(n_612),
.Y(n_730)
);

OAI21x1_ASAP7_75t_L g731 ( 
.A1(n_668),
.A2(n_629),
.B(n_631),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_662),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_682),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_700),
.A2(n_629),
.B(n_633),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_670),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_660),
.B(n_614),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_658),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_703),
.B(n_602),
.Y(n_738)
);

CKINVDCx6p67_ASAP7_75t_R g739 ( 
.A(n_650),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_683),
.B(n_612),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_681),
.A2(n_633),
.B(n_603),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_676),
.A2(n_633),
.B(n_612),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_701),
.A2(n_633),
.B1(n_16),
.B2(n_17),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_703),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_677),
.B(n_15),
.Y(n_745)
);

OAI21x1_ASAP7_75t_L g746 ( 
.A1(n_691),
.A2(n_116),
.B(n_201),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_685),
.A2(n_15),
.B1(n_19),
.B2(n_20),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_678),
.A2(n_117),
.B(n_200),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_687),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_686),
.B(n_63),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_653),
.B(n_19),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_686),
.B(n_64),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_L g753 ( 
.A(n_696),
.B(n_65),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_657),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_671),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_724),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_717),
.B(n_698),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_SL g758 ( 
.A(n_743),
.B(n_656),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_716),
.B(n_697),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_706),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_SL g761 ( 
.A1(n_753),
.A2(n_667),
.B1(n_702),
.B2(n_688),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_732),
.B(n_655),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_L g763 ( 
.A1(n_707),
.A2(n_678),
.B1(n_673),
.B2(n_704),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_737),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_726),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_753),
.A2(n_719),
.B1(n_712),
.B2(n_725),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_705),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_726),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_723),
.A2(n_722),
.B1(n_721),
.B2(n_711),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_724),
.Y(n_770)
);

NAND3xp33_ASAP7_75t_SL g771 ( 
.A(n_748),
.B(n_675),
.C(n_694),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_735),
.B(n_698),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_738),
.B(n_698),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_755),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_726),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_719),
.A2(n_680),
.B1(n_21),
.B2(n_22),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_745),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_729),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_751),
.B(n_24),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_744),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_708),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_736),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_736),
.B(n_26),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_738),
.B(n_66),
.Y(n_784)
);

CKINVDCx11_ASAP7_75t_R g785 ( 
.A(n_739),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_708),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_747),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_733),
.Y(n_788)
);

CKINVDCx14_ASAP7_75t_R g789 ( 
.A(n_739),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_755),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_706),
.B(n_68),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_733),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_724),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_740),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_749),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_726),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_724),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_738),
.B(n_30),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_706),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_740),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_750),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_730),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_710),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_728),
.B(n_32),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_728),
.B(n_33),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_754),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_750),
.B(n_34),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_709),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_730),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_709),
.B(n_37),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_709),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_728),
.B(n_70),
.Y(n_812)
);

OAI221xp5_ASAP7_75t_L g813 ( 
.A1(n_758),
.A2(n_777),
.B1(n_766),
.B2(n_787),
.C(n_761),
.Y(n_813)
);

AOI221xp5_ASAP7_75t_L g814 ( 
.A1(n_758),
.A2(n_752),
.B1(n_750),
.B2(n_730),
.C(n_754),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_771),
.A2(n_752),
.B1(n_709),
.B2(n_754),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_801),
.B(n_752),
.Y(n_816)
);

OAI221xp5_ASAP7_75t_L g817 ( 
.A1(n_802),
.A2(n_718),
.B1(n_709),
.B2(n_741),
.C(n_742),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_763),
.A2(n_709),
.B1(n_741),
.B2(n_727),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_SL g819 ( 
.A1(n_804),
.A2(n_709),
.B1(n_727),
.B2(n_742),
.Y(n_819)
);

OAI221xp5_ASAP7_75t_L g820 ( 
.A1(n_809),
.A2(n_718),
.B1(n_713),
.B2(n_715),
.C(n_38),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_804),
.B(n_718),
.C(n_713),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_772),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_786),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_807),
.B(n_718),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_805),
.A2(n_720),
.B1(n_731),
.B2(n_714),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_759),
.B(n_71),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_805),
.A2(n_720),
.B1(n_731),
.B2(n_714),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_800),
.B(n_718),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_SL g829 ( 
.A1(n_794),
.A2(n_746),
.B1(n_710),
.B2(n_734),
.Y(n_829)
);

OAI22xp33_ASAP7_75t_L g830 ( 
.A1(n_762),
.A2(n_38),
.B1(n_39),
.B2(n_734),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_780),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_776),
.A2(n_746),
.B1(n_39),
.B2(n_75),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_810),
.A2(n_779),
.B1(n_778),
.B2(n_806),
.Y(n_833)
);

OAI22xp33_ASAP7_75t_L g834 ( 
.A1(n_810),
.A2(n_73),
.B1(n_78),
.B2(n_81),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_782),
.B(n_83),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_756),
.Y(n_836)
);

OAI211xp5_ASAP7_75t_L g837 ( 
.A1(n_783),
.A2(n_84),
.B(n_86),
.C(n_87),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_798),
.B(n_88),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_764),
.B(n_90),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_793),
.B(n_91),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_790),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_841)
);

AOI221xp5_ASAP7_75t_L g842 ( 
.A1(n_769),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.C(n_101),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_L g843 ( 
.A(n_790),
.B(n_107),
.Y(n_843)
);

AOI221xp5_ASAP7_75t_L g844 ( 
.A1(n_812),
.A2(n_118),
.B1(n_122),
.B2(n_123),
.C(n_126),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_788),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_767),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_SL g847 ( 
.A1(n_812),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_784),
.A2(n_131),
.B1(n_135),
.B2(n_141),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_801),
.A2(n_143),
.B(n_146),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_774),
.A2(n_147),
.B1(n_148),
.B2(n_151),
.Y(n_850)
);

OAI22xp33_ASAP7_75t_L g851 ( 
.A1(n_801),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_851)
);

OAI21x1_ASAP7_75t_L g852 ( 
.A1(n_803),
.A2(n_155),
.B(n_156),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_767),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_789),
.A2(n_157),
.B1(n_159),
.B2(n_161),
.Y(n_854)
);

OAI22xp33_ASAP7_75t_L g855 ( 
.A1(n_784),
.A2(n_163),
.B1(n_164),
.B2(n_167),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_795),
.B(n_168),
.Y(n_856)
);

AOI221xp5_ASAP7_75t_L g857 ( 
.A1(n_757),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.C(n_175),
.Y(n_857)
);

NAND3xp33_ASAP7_75t_L g858 ( 
.A(n_784),
.B(n_176),
.C(n_177),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_773),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_824),
.B(n_757),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_822),
.B(n_773),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_853),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_846),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_846),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_R g865 ( 
.A(n_843),
.B(n_789),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_828),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_813),
.A2(n_768),
.B1(n_765),
.B2(n_796),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_823),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_845),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_833),
.A2(n_768),
.B1(n_765),
.B2(n_796),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_831),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_836),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_821),
.B(n_773),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_819),
.B(n_792),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_817),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_852),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_819),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_825),
.B(n_792),
.Y(n_878)
);

NOR2x1_ASAP7_75t_L g879 ( 
.A(n_834),
.B(n_811),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_827),
.B(n_781),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_836),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_818),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_820),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_814),
.B(n_781),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_836),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_836),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_829),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_856),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_835),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_815),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_R g891 ( 
.A(n_872),
.B(n_785),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_868),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_868),
.Y(n_893)
);

OAI31xp33_ASAP7_75t_L g894 ( 
.A1(n_883),
.A2(n_834),
.A3(n_830),
.B(n_832),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_868),
.Y(n_895)
);

OAI222xp33_ASAP7_75t_L g896 ( 
.A1(n_890),
.A2(n_883),
.B1(n_887),
.B2(n_877),
.C1(n_867),
.C2(n_847),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_SL g897 ( 
.A1(n_865),
.A2(n_858),
.B1(n_837),
.B2(n_826),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_885),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_860),
.B(n_803),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_860),
.B(n_873),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_869),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_869),
.Y(n_902)
);

NOR2x1_ASAP7_75t_L g903 ( 
.A(n_879),
.B(n_808),
.Y(n_903)
);

OAI21xp33_ASAP7_75t_L g904 ( 
.A1(n_875),
.A2(n_847),
.B(n_842),
.Y(n_904)
);

NAND2xp33_ASAP7_75t_R g905 ( 
.A(n_877),
.B(n_839),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_869),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_L g907 ( 
.A(n_870),
.B(n_844),
.C(n_854),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_866),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_871),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_SL g910 ( 
.A1(n_890),
.A2(n_829),
.B1(n_859),
.B2(n_848),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_900),
.B(n_873),
.Y(n_911)
);

AOI32xp33_ASAP7_75t_L g912 ( 
.A1(n_903),
.A2(n_887),
.A3(n_875),
.B1(n_879),
.B2(n_851),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_900),
.B(n_875),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_908),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_901),
.Y(n_915)
);

INVxp67_ASAP7_75t_SL g916 ( 
.A(n_903),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_906),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_908),
.B(n_866),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_901),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_899),
.B(n_874),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_899),
.B(n_874),
.Y(n_921)
);

OR2x6_ASAP7_75t_L g922 ( 
.A(n_910),
.B(n_884),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_898),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_898),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_906),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_906),
.B(n_861),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_911),
.B(n_909),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_913),
.B(n_918),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_911),
.B(n_906),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_920),
.B(n_909),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_915),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_915),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_920),
.B(n_893),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_921),
.B(n_901),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_932),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_928),
.Y(n_936)
);

OAI211xp5_ASAP7_75t_SL g937 ( 
.A1(n_930),
.A2(n_912),
.B(n_894),
.C(n_904),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_932),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_927),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_934),
.B(n_918),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_929),
.B(n_914),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_937),
.A2(n_922),
.B(n_896),
.C(n_904),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_936),
.A2(n_922),
.B(n_916),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_935),
.B(n_922),
.C(n_894),
.Y(n_944)
);

OAI21xp33_ASAP7_75t_L g945 ( 
.A1(n_936),
.A2(n_922),
.B(n_897),
.Y(n_945)
);

AOI31xp33_ASAP7_75t_L g946 ( 
.A1(n_945),
.A2(n_905),
.A3(n_785),
.B(n_938),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_942),
.A2(n_907),
.B(n_941),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_944),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_948),
.Y(n_949)
);

NAND2x1p5_ASAP7_75t_L g950 ( 
.A(n_946),
.B(n_943),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_947),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_948),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_951),
.B(n_939),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_950),
.B(n_941),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_950),
.Y(n_955)
);

AOI21xp33_ASAP7_75t_SL g956 ( 
.A1(n_949),
.A2(n_940),
.B(n_891),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_952),
.A2(n_849),
.B(n_851),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_951),
.B(n_929),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_951),
.A2(n_850),
.B(n_857),
.Y(n_959)
);

AOI221xp5_ASAP7_75t_L g960 ( 
.A1(n_955),
.A2(n_910),
.B1(n_914),
.B2(n_855),
.C(n_882),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_954),
.A2(n_882),
.B1(n_888),
.B2(n_889),
.Y(n_961)
);

OAI221xp5_ASAP7_75t_SL g962 ( 
.A1(n_953),
.A2(n_838),
.B1(n_934),
.B2(n_931),
.C(n_933),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_958),
.A2(n_886),
.B1(n_885),
.B2(n_816),
.Y(n_963)
);

AOI221xp5_ASAP7_75t_L g964 ( 
.A1(n_956),
.A2(n_841),
.B1(n_924),
.B2(n_923),
.C(n_886),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_959),
.A2(n_919),
.B(n_871),
.Y(n_965)
);

NAND4xp25_ASAP7_75t_L g966 ( 
.A(n_957),
.B(n_840),
.C(n_816),
.D(n_881),
.Y(n_966)
);

NAND3x2_ASAP7_75t_L g967 ( 
.A(n_962),
.B(n_921),
.C(n_884),
.Y(n_967)
);

AO22x2_ASAP7_75t_L g968 ( 
.A1(n_965),
.A2(n_925),
.B1(n_917),
.B2(n_919),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_960),
.B(n_926),
.Y(n_969)
);

NOR3xp33_ASAP7_75t_L g970 ( 
.A(n_966),
.B(n_791),
.C(n_775),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_SL g971 ( 
.A1(n_963),
.A2(n_888),
.B(n_885),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_964),
.A2(n_881),
.B1(n_888),
.B2(n_889),
.Y(n_972)
);

NAND4xp75_ASAP7_75t_L g973 ( 
.A(n_961),
.B(n_775),
.C(n_791),
.D(n_926),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_969),
.B(n_925),
.Y(n_974)
);

NAND4xp75_ASAP7_75t_L g975 ( 
.A(n_972),
.B(n_893),
.C(n_917),
.D(n_880),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_968),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_970),
.B(n_797),
.C(n_770),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_967),
.B(n_797),
.Y(n_978)
);

AND3x2_ASAP7_75t_L g979 ( 
.A(n_973),
.B(n_889),
.C(n_876),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_971),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_970),
.A2(n_881),
.B1(n_876),
.B2(n_902),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_L g982 ( 
.A(n_972),
.B(n_797),
.C(n_770),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_969),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_983),
.B(n_902),
.Y(n_984)
);

AOI221xp5_ASAP7_75t_SL g985 ( 
.A1(n_978),
.A2(n_797),
.B1(n_770),
.B2(n_756),
.C(n_876),
.Y(n_985)
);

AOI221xp5_ASAP7_75t_L g986 ( 
.A1(n_980),
.A2(n_770),
.B1(n_756),
.B2(n_863),
.C(n_864),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_976),
.Y(n_987)
);

NAND3xp33_ASAP7_75t_L g988 ( 
.A(n_982),
.B(n_756),
.C(n_799),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_974),
.B(n_895),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_977),
.A2(n_880),
.B1(n_878),
.B2(n_861),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_975),
.Y(n_991)
);

NAND4xp25_ASAP7_75t_L g992 ( 
.A(n_981),
.B(n_878),
.C(n_864),
.D(n_863),
.Y(n_992)
);

NOR4xp25_ASAP7_75t_L g993 ( 
.A(n_979),
.B(n_895),
.C(n_892),
.D(n_862),
.Y(n_993)
);

INVxp67_ASAP7_75t_SL g994 ( 
.A(n_976),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_994),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_987),
.B(n_892),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_991),
.B(n_862),
.Y(n_997)
);

INVx8_ASAP7_75t_L g998 ( 
.A(n_985),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_SL g999 ( 
.A(n_984),
.B(n_760),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_986),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_995),
.B(n_989),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_996),
.Y(n_1002)
);

OAI22x1_ASAP7_75t_L g1003 ( 
.A1(n_1000),
.A2(n_988),
.B1(n_993),
.B2(n_992),
.Y(n_1003)
);

AOI21xp33_ASAP7_75t_SL g1004 ( 
.A1(n_1003),
.A2(n_998),
.B(n_997),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_1002),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_1005),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_1004),
.B(n_1001),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_1007),
.A2(n_998),
.B(n_999),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_1006),
.B(n_990),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_1009),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_1010),
.A2(n_1008),
.B1(n_862),
.B2(n_760),
.Y(n_1011)
);

OAI221xp5_ASAP7_75t_R g1012 ( 
.A1(n_1011),
.A2(n_184),
.B1(n_186),
.B2(n_191),
.C(n_193),
.Y(n_1012)
);

AOI211xp5_ASAP7_75t_L g1013 ( 
.A1(n_1012),
.A2(n_194),
.B(n_196),
.C(n_197),
.Y(n_1013)
);


endmodule