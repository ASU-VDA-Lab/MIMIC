module fake_jpeg_4516_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_12),
.Y(n_69)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_52),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_19),
.B1(n_16),
.B2(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_64),
.B1(n_71),
.B2(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_27),
.B1(n_18),
.B2(n_31),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_53),
.B1(n_30),
.B2(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_27),
.B1(n_31),
.B2(n_24),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_55),
.Y(n_89)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_28),
.B(n_29),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_25),
.B(n_32),
.C(n_30),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_28),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_23),
.Y(n_88)
);

CKINVDCx12_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_29),
.B1(n_33),
.B2(n_23),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_33),
.B1(n_25),
.B2(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_33),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_57),
.B1(n_55),
.B2(n_68),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_23),
.B1(n_25),
.B2(n_13),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_0),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_30),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_62),
.CI(n_46),
.CON(n_102),
.SN(n_102)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_50),
.B1(n_62),
.B2(n_58),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_103),
.B1(n_108),
.B2(n_117),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_102),
.B(n_61),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_58),
.B1(n_67),
.B2(n_56),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_54),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_25),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_47),
.C(n_66),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_117),
.C(n_109),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_55),
.B1(n_57),
.B2(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_56),
.B1(n_63),
.B2(n_47),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_110),
.B1(n_119),
.B2(n_94),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_43),
.B1(n_39),
.B2(n_45),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_83),
.B(n_93),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_74),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_118),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_43),
.B1(n_65),
.B2(n_45),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_74),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_45),
.B1(n_65),
.B2(n_70),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_87),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_128),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_93),
.B1(n_88),
.B2(n_87),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_131),
.B1(n_119),
.B2(n_101),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_121),
.B1(n_98),
.B2(n_103),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_78),
.B1(n_86),
.B2(n_83),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_102),
.Y(n_163)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_145),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_102),
.B(n_112),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_136),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_73),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_73),
.B(n_80),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_141),
.B(n_120),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_72),
.B(n_81),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_149),
.C(n_151),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_143),
.B(n_144),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_107),
.B(n_69),
.CI(n_94),
.CON(n_144),
.SN(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_102),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_80),
.C(n_95),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_150),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_96),
.C(n_86),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_154),
.Y(n_192)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_169),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_158),
.A2(n_116),
.B(n_82),
.Y(n_197)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_161),
.B(n_162),
.Y(n_182)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_174),
.B(n_175),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_149),
.C(n_127),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_177),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_101),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_147),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_108),
.B1(n_78),
.B2(n_94),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_151),
.B1(n_124),
.B2(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_126),
.A2(n_145),
.B1(n_136),
.B2(n_135),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_140),
.A2(n_146),
.B1(n_144),
.B2(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_140),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_128),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_198),
.Y(n_217)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_188),
.B1(n_205),
.B2(n_152),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_142),
.B1(n_125),
.B2(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_191),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_133),
.C(n_141),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_171),
.B1(n_173),
.B2(n_159),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_193),
.A2(n_156),
.B1(n_179),
.B2(n_177),
.Y(n_213)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_196),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_162),
.B(n_169),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_105),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_105),
.C(n_116),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_202),
.Y(n_227)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_165),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_204),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_65),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_154),
.A2(n_78),
.B1(n_97),
.B2(n_26),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_0),
.B(n_1),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_1),
.B(n_3),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_207),
.A2(n_220),
.B(n_232),
.Y(n_247)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_208),
.A2(n_3),
.B(n_4),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_152),
.B1(n_163),
.B2(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_221),
.B1(n_184),
.B2(n_181),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_226),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_205),
.B1(n_188),
.B2(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_160),
.B1(n_157),
.B2(n_26),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_160),
.B1(n_153),
.B2(n_20),
.Y(n_221)
);

XOR2x2_ASAP7_75t_SL g222 ( 
.A(n_203),
.B(n_15),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_206),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_225),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_182),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_0),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_181),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_231),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_180),
.C(n_191),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_242),
.C(n_254),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_190),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_248),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_187),
.B1(n_204),
.B2(n_194),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_198),
.C(n_187),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_231),
.B1(n_220),
.B2(n_223),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_14),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_225),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_14),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_253),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_14),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_13),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_240),
.B(n_222),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_259),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_213),
.B1(n_208),
.B2(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_212),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_270),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_SL g287 ( 
.A(n_258),
.B(n_262),
.C(n_12),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_219),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_215),
.B(n_228),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_265),
.B(n_245),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_247),
.B1(n_242),
.B2(n_229),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_251),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_210),
.B(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_248),
.B(n_250),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_272),
.C(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_233),
.B(n_223),
.C(n_218),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_275),
.B(n_282),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_283),
.C(n_263),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_252),
.B1(n_247),
.B2(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_229),
.B1(n_239),
.B2(n_7),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_281),
.B(n_289),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_5),
.C(n_6),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_262),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_258),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_10),
.C(n_6),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_265),
.Y(n_289)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_291),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_5),
.B(n_6),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_267),
.C(n_259),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_294),
.A2(n_299),
.B(n_8),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_273),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_297),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_273),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_275),
.B(n_264),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_255),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_282),
.B1(n_286),
.B2(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_8),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_271),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_8),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_298),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_305),
.B(n_308),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_310),
.C(n_312),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_SL g307 ( 
.A1(n_291),
.A2(n_277),
.B(n_283),
.C(n_7),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_307),
.A2(n_314),
.B(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_10),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_295),
.B1(n_9),
.B2(n_296),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_9),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_290),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_321),
.B(n_314),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_320),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_300),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_307),
.Y(n_324)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_318),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_297),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_324),
.A2(n_327),
.B(n_328),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_325),
.A2(n_322),
.B(n_9),
.Y(n_329)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_319),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_326),
.Y(n_331)
);

AOI21x1_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_330),
.B(n_323),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);


endmodule