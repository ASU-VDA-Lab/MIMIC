module fake_jpeg_6542_n_308 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_308);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_13),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_49),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx9p33_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_22),
.B1(n_27),
.B2(n_24),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_27),
.B1(n_36),
.B2(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_13),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_16),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_34),
.B(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_65),
.B1(n_27),
.B2(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_35),
.B1(n_16),
.B2(n_27),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_71),
.Y(n_90)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_76),
.B(n_78),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_83),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_93),
.B1(n_96),
.B2(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_41),
.C(n_42),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_95),
.C(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_89),
.Y(n_101)
);

AOI22x1_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_51),
.B1(n_36),
.B2(n_16),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_39),
.B1(n_71),
.B2(n_70),
.Y(n_107)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_92),
.Y(n_116)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_19),
.Y(n_115)
);

XOR2x2_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_45),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_64),
.B1(n_74),
.B2(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_20),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_104),
.Y(n_138)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_100),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_65),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_113),
.C(n_80),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_109),
.B(n_24),
.Y(n_139)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_108),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_118),
.B1(n_88),
.B2(n_46),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_92),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_112),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_54),
.B1(n_44),
.B2(n_45),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_93),
.B1(n_79),
.B2(n_89),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_77),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_72),
.C(n_56),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_17),
.B(n_20),
.Y(n_142)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_44),
.B1(n_70),
.B2(n_56),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_17),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_79),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_129),
.B1(n_143),
.B2(n_118),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_130),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_112),
.B1(n_109),
.B2(n_69),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_141),
.B(n_25),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_88),
.B1(n_55),
.B2(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_133),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_137),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_139),
.A2(n_142),
.B(n_114),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_15),
.B1(n_26),
.B2(n_17),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_100),
.A2(n_46),
.B1(n_53),
.B2(n_20),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_156),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_138),
.A2(n_115),
.B(n_104),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_167),
.B(n_168),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_151),
.C(n_29),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_104),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_132),
.B1(n_130),
.B2(n_125),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_100),
.B(n_105),
.C(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_163),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_137),
.B(n_117),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_124),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_134),
.B1(n_144),
.B2(n_140),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_18),
.B1(n_19),
.B2(n_32),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_113),
.B(n_105),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_25),
.B(n_26),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_117),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_108),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_162),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_136),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_53),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

AO32x1_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_16),
.A3(n_14),
.B1(n_108),
.B2(n_75),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_46),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_126),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_187),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_190),
.B1(n_192),
.B2(n_158),
.Y(n_200)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_180),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_195),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_145),
.B(n_99),
.Y(n_180)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_183),
.Y(n_212)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_149),
.C(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_25),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_19),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_196),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_152),
.B1(n_148),
.B2(n_156),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_201),
.C(n_204),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_172),
.B(n_147),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_202),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_182),
.B1(n_183),
.B2(n_179),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_196),
.B1(n_195),
.B2(n_193),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_200),
.A2(n_214),
.B1(n_18),
.B2(n_53),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_171),
.C(n_153),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_155),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_177),
.A2(n_171),
.B1(n_169),
.B2(n_158),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_170),
.B1(n_150),
.B2(n_176),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_163),
.C(n_146),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_146),
.C(n_159),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_208),
.C(n_188),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_164),
.C(n_168),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_170),
.B1(n_150),
.B2(n_91),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_194),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_185),
.B(n_175),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_235),
.B1(n_211),
.B2(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_223),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_150),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_215),
.B1(n_210),
.B2(n_216),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_170),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_228),
.Y(n_245)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_236),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_185),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_234),
.B(n_14),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_201),
.C(n_197),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_187),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_SL g255 ( 
.A(n_232),
.B(n_237),
.C(n_32),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_190),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_217),
.Y(n_241)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_205),
.B(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_32),
.Y(n_251)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_14),
.C(n_23),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_234),
.A2(n_18),
.B1(n_81),
.B2(n_91),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_253),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_81),
.B1(n_75),
.B2(n_23),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_247),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_270)
);

BUFx12f_ASAP7_75t_SL g250 ( 
.A(n_237),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_250),
.A2(n_231),
.B(n_226),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_230),
.Y(n_252)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_23),
.B1(n_31),
.B2(n_29),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_219),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_269),
.B(n_245),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_SL g259 ( 
.A(n_250),
.B(n_226),
.C(n_232),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_239),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_219),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_263),
.C(n_266),
.Y(n_274)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_31),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_31),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_268),
.C(n_265),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_262),
.A2(n_252),
.B1(n_254),
.B2(n_248),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_268),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_4),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_277),
.B(n_279),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_282),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_247),
.B(n_1),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_256),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_4),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_0),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_1),
.Y(n_281)
);

AOI31xp67_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_261),
.A3(n_2),
.B(n_3),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_257),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_289),
.B(n_292),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_284),
.B(n_291),
.Y(n_294)
);

AOI31xp67_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_277),
.A3(n_282),
.B(n_274),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_5),
.Y(n_298)
);

AOI31xp67_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_263),
.A3(n_267),
.B(n_3),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_280),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_296),
.B(n_297),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_290),
.B(n_5),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_11),
.Y(n_297)
);

OAI21xp33_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_5),
.B(n_6),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_294),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_6),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.C(n_300),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_285),
.C2(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_8),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_8),
.B(n_10),
.Y(n_308)
);


endmodule