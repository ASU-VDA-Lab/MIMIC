module fake_jpeg_27591_n_172 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx6p67_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_34),
.Y(n_38)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_2),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_21),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_16),
.C(n_26),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_46),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_23),
.B(n_28),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_19),
.B(n_24),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_17),
.C(n_26),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_14),
.B1(n_24),
.B2(n_17),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_22),
.B1(n_25),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_34),
.B1(n_31),
.B2(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_54),
.B(n_20),
.Y(n_86)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_33),
.B(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_23),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_19),
.B1(n_32),
.B2(n_18),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_42),
.B1(n_20),
.B2(n_4),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_65),
.B1(n_67),
.B2(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_63),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_46),
.B1(n_34),
.B2(n_31),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_70),
.Y(n_83)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_34),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_45),
.C(n_3),
.Y(n_90)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_92),
.Y(n_95)
);

BUFx24_ASAP7_75t_SL g78 ( 
.A(n_66),
.Y(n_78)
);

BUFx24_ASAP7_75t_SL g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_70),
.B1(n_59),
.B2(n_6),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_85),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_63),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_89),
.B1(n_64),
.B2(n_53),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_93),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_20),
.B1(n_45),
.B2(n_4),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_99),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_67),
.B(n_62),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

OAI221xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_109),
.B1(n_12),
.B2(n_11),
.C(n_6),
.Y(n_126)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_108),
.B(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_58),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_2),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_89),
.B1(n_80),
.B2(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_115),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_92),
.C(n_76),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_116),
.C(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_74),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_111),
.A2(n_81),
.B1(n_91),
.B2(n_85),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_123),
.B(n_126),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_121),
.B1(n_107),
.B2(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_127),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_90),
.B1(n_79),
.B2(n_75),
.Y(n_121)
);

NOR2x1_ASAP7_75t_R g123 ( 
.A(n_100),
.B(n_110),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_79),
.C(n_13),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_132),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_137),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_105),
.Y(n_132)
);

OAI321xp33_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_119),
.A3(n_122),
.B1(n_118),
.B2(n_109),
.C(n_117),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_135),
.A2(n_12),
.B(n_79),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_104),
.C(n_99),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_96),
.C(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_5),
.C(n_7),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_129),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_148),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_106),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

AO221x1_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_129),
.B1(n_139),
.B2(n_132),
.C(n_9),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_153),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_154),
.C(n_155),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_136),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_144),
.B1(n_145),
.B2(n_142),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_8),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g160 ( 
.A(n_152),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_155),
.B(n_143),
.Y(n_161)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_8),
.CI(n_9),
.CON(n_163),
.SN(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_9),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_8),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_168),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_166),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_163),
.B(n_169),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_163),
.Y(n_172)
);


endmodule