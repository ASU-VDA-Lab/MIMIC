module fake_netlist_6_3859_n_1856 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1856);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1856;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_131),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_15),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_109),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_91),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_20),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_83),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_5),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_73),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_72),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_33),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_124),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_108),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_16),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_71),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_140),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_153),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_36),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_139),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_86),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_38),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_34),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_49),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_50),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_77),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_10),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_80),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_15),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_84),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_146),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_134),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_113),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_10),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_54),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_128),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_13),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_27),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_47),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_52),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_121),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_81),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_106),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_47),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_110),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_44),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_63),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_45),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_96),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_12),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_23),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_32),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_142),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_103),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_62),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_67),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_129),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_119),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_18),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_1),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_115),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_169),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_166),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_59),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_41),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_90),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_1),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_23),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_18),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_14),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_118),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_42),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_75),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_92),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_31),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_101),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_29),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_85),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_20),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_97),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_8),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_70),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_126),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_163),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_94),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_14),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_82),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_167),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_159),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_62),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_148),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_2),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_74),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_53),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_13),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_104),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_32),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_105),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_44),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_28),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_164),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_58),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_78),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_123),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_144),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_39),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_93),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_69),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_61),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_165),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_7),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_88),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_162),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_149),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_87),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_51),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_36),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_59),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_114),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_63),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_5),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_52),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_37),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_61),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_48),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_89),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_117),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_3),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_33),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_40),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_46),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_4),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_25),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_12),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_31),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_116),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_112),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_99),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_100),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_98),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_51),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_19),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_95),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_21),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_21),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_35),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_111),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_53),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_58),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_40),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_22),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_9),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_155),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_251),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_170),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_251),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_176),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_174),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_175),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_209),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_177),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_199),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_310),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_242),
.B(n_0),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_178),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_180),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_240),
.B(n_2),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_212),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_173),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_182),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_242),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_187),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_209),
.B(n_4),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_310),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_310),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_174),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_238),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_238),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_309),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_203),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_258),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_188),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_190),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_191),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_240),
.B(n_6),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_258),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_192),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_218),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_232),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_173),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_235),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_302),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_292),
.B(n_6),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_302),
.B(n_8),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_194),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_171),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_250),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_181),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_171),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_260),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_292),
.B(n_9),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_321),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_181),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_189),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_189),
.Y(n_388)
);

INVxp33_ASAP7_75t_SL g389 ( 
.A(n_172),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_193),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_173),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_193),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_239),
.B(n_11),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_195),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_210),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_205),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_210),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_206),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_211),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_211),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_233),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_208),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_233),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_256),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_256),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_219),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_220),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_246),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_314),
.B(n_16),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_183),
.B(n_17),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_246),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_247),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_247),
.B(n_17),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_231),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_248),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_234),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_248),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_179),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_236),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_260),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_249),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_241),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_249),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_244),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_254),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_351),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_340),
.B(n_345),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_351),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_183),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_351),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_349),
.B(n_200),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_373),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_373),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_356),
.B(n_260),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_391),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_346),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_357),
.B(n_239),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_358),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_358),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_334),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_413),
.B(n_264),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_393),
.B(n_264),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_360),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_360),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_349),
.B(n_267),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_361),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_361),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_364),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_369),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_369),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_375),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_375),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_418),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_393),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_381),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_328),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_404),
.B(n_314),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_381),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_386),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_346),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_410),
.B(n_328),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_335),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_383),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

AND3x2_ASAP7_75t_L g479 ( 
.A(n_368),
.B(n_186),
.C(n_184),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_390),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_354),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_354),
.Y(n_484)
);

CKINVDCx6p67_ASAP7_75t_R g485 ( 
.A(n_363),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_379),
.B(n_334),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_347),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_425),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_396),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_382),
.B(n_184),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_392),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_392),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_397),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_399),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_376),
.B(n_299),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_399),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_401),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

OA21x2_ASAP7_75t_L g503 ( 
.A1(n_403),
.A2(n_259),
.B(n_254),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_350),
.A2(n_213),
.B1(n_277),
.B2(n_197),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_503),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_464),
.B(n_173),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_503),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_503),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_503),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_464),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_496),
.B(n_389),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_467),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_405),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_429),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_429),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_433),
.B(n_336),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_342),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_503),
.Y(n_518)
);

INVxp33_ASAP7_75t_SL g519 ( 
.A(n_482),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_429),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_482),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_429),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_429),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_429),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_496),
.B(n_433),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_L g526 ( 
.A(n_464),
.B(n_173),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_431),
.B(n_186),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_503),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_503),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_446),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_465),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_454),
.B(n_384),
.C(n_341),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_464),
.Y(n_533)
);

OR2x6_ASAP7_75t_L g534 ( 
.A(n_467),
.B(n_395),
.Y(n_534)
);

OAI22xp33_ASAP7_75t_L g535 ( 
.A1(n_439),
.A2(n_473),
.B1(n_454),
.B2(n_451),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_439),
.B(n_363),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_463),
.B(n_338),
.Y(n_537)
);

AND3x2_ASAP7_75t_L g538 ( 
.A(n_442),
.B(n_337),
.C(n_207),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_464),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

AND2x6_ASAP7_75t_L g541 ( 
.A(n_464),
.B(n_201),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_446),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_463),
.B(n_343),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_464),
.B(n_348),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_473),
.A2(n_337),
.B1(n_377),
.B2(n_274),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_464),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_467),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_468),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_473),
.A2(n_377),
.B1(n_274),
.B2(n_297),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_468),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_442),
.B(n_352),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_435),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_446),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_435),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_468),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_464),
.B(n_355),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_464),
.B(n_365),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_485),
.B(n_402),
.Y(n_560)
);

AND2x6_ASAP7_75t_L g561 ( 
.A(n_431),
.B(n_449),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_476),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_469),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_446),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_486),
.B(n_366),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_486),
.B(n_490),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_476),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_476),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_469),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_467),
.B(n_383),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_447),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_484),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_469),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_471),
.B(n_367),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_445),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_471),
.B(n_370),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_490),
.B(n_378),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_490),
.B(n_394),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_470),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_447),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_490),
.B(n_398),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_435),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_487),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_451),
.B(n_406),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_445),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_451),
.B(n_407),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_431),
.B(n_419),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_470),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_475),
.B(n_383),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_447),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_470),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_431),
.B(n_424),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_472),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_435),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_472),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_449),
.B(n_414),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_447),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_476),
.Y(n_598)
);

INVxp67_ASAP7_75t_SL g599 ( 
.A(n_445),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_485),
.B(n_416),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_420),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_427),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_435),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_472),
.Y(n_604)
);

INVx11_ASAP7_75t_L g605 ( 
.A(n_485),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_479),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_435),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_484),
.B(n_420),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_476),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_435),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_427),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_449),
.B(n_420),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_449),
.A2(n_303),
.B1(n_259),
.B2(n_300),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_477),
.Y(n_614)
);

INVxp67_ASAP7_75t_SL g615 ( 
.A(n_435),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_435),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_477),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_479),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_435),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_SL g620 ( 
.A(n_450),
.B(n_282),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_428),
.B(n_339),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_428),
.B(n_422),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_477),
.B(n_362),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_427),
.Y(n_624)
);

OR2x6_ASAP7_75t_L g625 ( 
.A(n_450),
.B(n_297),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_497),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_450),
.A2(n_300),
.B1(n_303),
.B2(n_313),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_434),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_R g629 ( 
.A(n_489),
.B(n_185),
.Y(n_629)
);

INVx4_ASAP7_75t_SL g630 ( 
.A(n_450),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_450),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_497),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_478),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_450),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_478),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_476),
.B(n_466),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_476),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_466),
.B(n_260),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_478),
.Y(n_639)
);

AND3x1_ASAP7_75t_L g640 ( 
.A(n_483),
.B(n_315),
.C(n_313),
.Y(n_640)
);

AND2x6_ASAP7_75t_L g641 ( 
.A(n_466),
.B(n_201),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_440),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_440),
.Y(n_643)
);

INVx6_ASAP7_75t_L g644 ( 
.A(n_476),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_466),
.B(n_315),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_434),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_466),
.B(n_207),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_434),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_436),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_480),
.A2(n_322),
.B1(n_326),
.B2(n_224),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_436),
.Y(n_651)
);

CKINVDCx11_ASAP7_75t_R g652 ( 
.A(n_487),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_489),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_440),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_483),
.B(n_408),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_483),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_652),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_508),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_521),
.Y(n_659)
);

NOR3xp33_ASAP7_75t_L g660 ( 
.A(n_511),
.B(n_504),
.C(n_198),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_561),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_575),
.B(n_480),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_535),
.A2(n_372),
.B1(n_374),
.B2(n_371),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_585),
.B(n_480),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_655),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_599),
.B(n_480),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_508),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_655),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_510),
.B(n_476),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_584),
.B(n_480),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_605),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_514),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_586),
.B(n_480),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_514),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_533),
.B(n_488),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_510),
.B(n_476),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_520),
.Y(n_677)
);

OAI22x1_ASAP7_75t_SL g678 ( 
.A1(n_583),
.A2(n_323),
.B1(n_289),
.B2(n_286),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_631),
.B(n_488),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_508),
.Y(n_680)
);

OAI221xp5_ASAP7_75t_L g681 ( 
.A1(n_525),
.A2(n_226),
.B1(n_322),
.B2(n_326),
.C(n_276),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_561),
.B(n_215),
.Y(n_682)
);

AND2x2_ASAP7_75t_SL g683 ( 
.A(n_544),
.B(n_558),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_631),
.B(n_634),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_560),
.B(n_485),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_510),
.B(n_306),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_520),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_539),
.B(n_306),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_561),
.A2(n_581),
.B1(n_577),
.B2(n_513),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_516),
.B(n_380),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_508),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_634),
.B(n_488),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_566),
.A2(n_512),
.B1(n_547),
.B2(n_565),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_561),
.B(n_488),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_521),
.B(n_359),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_519),
.B(n_385),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_508),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_523),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_572),
.B(n_309),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_513),
.B(n_309),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_512),
.B(n_547),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_519),
.B(n_504),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_570),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_570),
.Y(n_704)
);

AOI211xp5_ASAP7_75t_L g705 ( 
.A1(n_532),
.A2(n_504),
.B(n_621),
.C(n_596),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_612),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_539),
.B(n_306),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_621),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_523),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_561),
.B(n_488),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_539),
.B(n_306),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_561),
.B(n_488),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_592),
.B(n_491),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_543),
.B(n_196),
.Y(n_714)
);

OAI221xp5_ASAP7_75t_L g715 ( 
.A1(n_551),
.A2(n_294),
.B1(n_281),
.B2(n_253),
.C(n_252),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_518),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_630),
.B(n_306),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_546),
.B(n_491),
.Y(n_718)
);

BUFx5_ASAP7_75t_L g719 ( 
.A(n_546),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_518),
.A2(n_491),
.B1(n_494),
.B2(n_223),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_515),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_630),
.B(n_491),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_559),
.B(n_491),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_517),
.B(n_309),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_531),
.B(n_491),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_630),
.B(n_494),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_647),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_518),
.A2(n_494),
.B1(n_285),
.B2(n_290),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_R g729 ( 
.A(n_629),
.B(n_620),
.Y(n_729)
);

AND2x2_ASAP7_75t_SL g730 ( 
.A(n_506),
.B(n_215),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_630),
.B(n_518),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_518),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_550),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_524),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_550),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_531),
.B(n_494),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_534),
.B(n_589),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_552),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_540),
.B(n_494),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_515),
.B(n_494),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_552),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_515),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_647),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_524),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_534),
.B(n_499),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_522),
.B(n_497),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_625),
.B(n_222),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_522),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_522),
.B(n_497),
.Y(n_749)
);

CKINVDCx14_ASAP7_75t_R g750 ( 
.A(n_622),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_536),
.B(n_204),
.C(n_202),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_578),
.B(n_497),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_505),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_587),
.A2(n_534),
.B1(n_527),
.B2(n_507),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_557),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_563),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_589),
.B(n_408),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_553),
.B(n_214),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_589),
.Y(n_759)
);

NOR2x1p5_ASAP7_75t_L g760 ( 
.A(n_605),
.B(n_216),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_540),
.B(n_548),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_527),
.A2(n_276),
.B1(n_222),
.B2(n_223),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_638),
.A2(n_278),
.B1(n_255),
.B2(n_257),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_505),
.A2(n_507),
.B(n_528),
.C(n_509),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_527),
.A2(n_285),
.B1(n_245),
.B2(n_252),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_563),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_574),
.B(n_217),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_569),
.Y(n_768)
);

OAI21xp33_ASAP7_75t_L g769 ( 
.A1(n_545),
.A2(n_412),
.B(n_411),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_548),
.B(n_497),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_SL g771 ( 
.A(n_600),
.B(n_265),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_549),
.B(n_497),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_549),
.B(n_497),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_589),
.B(n_601),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_647),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_569),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_509),
.B(n_497),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_641),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_573),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_528),
.B(n_497),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_541),
.A2(n_319),
.B1(n_245),
.B2(n_253),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_529),
.B(n_281),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_573),
.B(n_474),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_576),
.B(n_221),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_588),
.B(n_474),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_529),
.B(n_227),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_588),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_591),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_623),
.A2(n_284),
.B1(n_263),
.B2(n_268),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_601),
.B(n_499),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_591),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_595),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_595),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_604),
.B(n_262),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_604),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_614),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_614),
.B(n_474),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_606),
.A2(n_287),
.B1(n_290),
.B2(n_294),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_608),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_601),
.B(n_411),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_601),
.B(n_500),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_617),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_617),
.B(n_474),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_633),
.B(n_481),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_633),
.B(n_481),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_537),
.B(n_225),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_635),
.B(n_481),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_541),
.B(n_287),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_506),
.A2(n_500),
.B(n_501),
.C(n_502),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_625),
.B(n_308),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_635),
.B(n_481),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_606),
.A2(n_295),
.B1(n_283),
.B2(n_273),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_639),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_626),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_639),
.B(n_492),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_656),
.B(n_492),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_618),
.B(n_500),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_656),
.B(n_269),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_579),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_593),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_618),
.B(n_228),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_636),
.B(n_271),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_602),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_657),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_689),
.A2(n_627),
.B1(n_613),
.B2(n_625),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_672),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_714),
.A2(n_641),
.B1(n_541),
.B2(n_625),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_690),
.B(n_653),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_708),
.B(n_645),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_684),
.A2(n_526),
.B(n_615),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_706),
.B(n_645),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_723),
.A2(n_526),
.B(n_645),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_706),
.B(n_645),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_742),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_764),
.A2(n_567),
.B(n_562),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_752),
.A2(n_567),
.B(n_562),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_701),
.B(n_541),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_693),
.A2(n_624),
.B(n_651),
.C(n_628),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_674),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_752),
.A2(n_567),
.B(n_562),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_733),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_742),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_659),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_713),
.B(n_670),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_782),
.A2(n_664),
.B(n_662),
.Y(n_845)
);

BUFx12f_ASAP7_75t_L g846 ( 
.A(n_671),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_786),
.A2(n_541),
.B(n_602),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_806),
.A2(n_308),
.B(n_319),
.C(n_650),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_703),
.B(n_538),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_695),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_677),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_658),
.B(n_640),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_758),
.A2(n_611),
.B(n_651),
.C(n_649),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_658),
.A2(n_637),
.B(n_598),
.Y(n_854)
);

BUFx4f_ASAP7_75t_L g855 ( 
.A(n_737),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_742),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_665),
.B(n_412),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_673),
.B(n_541),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_668),
.B(n_641),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_687),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_698),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_658),
.A2(n_637),
.B(n_598),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_786),
.A2(n_780),
.B(n_777),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_658),
.B(n_732),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_733),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_732),
.B(n_288),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_732),
.B(n_293),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_703),
.B(n_641),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_767),
.A2(n_611),
.B(n_649),
.C(n_648),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_704),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_704),
.B(n_229),
.Y(n_871)
);

AOI21x1_ASAP7_75t_L g872 ( 
.A1(n_777),
.A2(n_628),
.B(n_624),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_735),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_732),
.Y(n_874)
);

INVx11_ASAP7_75t_L g875 ( 
.A(n_657),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_755),
.B(n_641),
.Y(n_876)
);

O2A1O1Ixp5_ASAP7_75t_L g877 ( 
.A1(n_754),
.A2(n_646),
.B(n_648),
.C(n_603),
.Y(n_877)
);

OAI21xp33_ASAP7_75t_L g878 ( 
.A1(n_821),
.A2(n_237),
.B(n_230),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_715),
.A2(n_646),
.B(n_501),
.C(n_530),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_745),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_709),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_735),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_782),
.A2(n_637),
.B(n_609),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_681),
.A2(n_501),
.B(n_542),
.C(n_590),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_762),
.A2(n_542),
.B(n_555),
.C(n_530),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_756),
.B(n_641),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_766),
.B(n_776),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_742),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_734),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_780),
.A2(n_564),
.B(n_555),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_661),
.A2(n_654),
.B1(n_643),
.B2(n_642),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_779),
.B(n_642),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_666),
.A2(n_609),
.B(n_568),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_738),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_787),
.B(n_642),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_744),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_675),
.A2(n_718),
.B(n_680),
.Y(n_897)
);

OAI21x1_ASAP7_75t_L g898 ( 
.A1(n_694),
.A2(n_556),
.B(n_554),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_792),
.B(n_643),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_802),
.B(n_643),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_819),
.B(n_654),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_667),
.A2(n_691),
.B(n_680),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_738),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_SL g904 ( 
.A1(n_710),
.A2(n_712),
.B(n_726),
.C(n_722),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_L g905 ( 
.A(n_705),
.B(n_307),
.C(n_332),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_820),
.B(n_554),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_753),
.B(n_554),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_721),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_798),
.A2(n_571),
.B(n_564),
.C(n_580),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_721),
.Y(n_910)
);

BUFx12f_ASAP7_75t_L g911 ( 
.A(n_671),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_682),
.A2(n_580),
.B1(n_590),
.B2(n_571),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_667),
.A2(n_697),
.B(n_691),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_697),
.A2(n_568),
.B(n_607),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_724),
.B(n_415),
.Y(n_915)
);

BUFx4f_ASAP7_75t_L g916 ( 
.A(n_774),
.Y(n_916)
);

BUFx4f_ASAP7_75t_L g917 ( 
.A(n_759),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_683),
.A2(n_743),
.B(n_727),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_741),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_784),
.A2(n_607),
.B(n_556),
.C(n_619),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_753),
.B(n_556),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_753),
.B(n_603),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_814),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_683),
.A2(n_603),
.B(n_607),
.Y(n_924)
);

AO21x1_ASAP7_75t_L g925 ( 
.A1(n_686),
.A2(n_597),
.B(n_436),
.Y(n_925)
);

BUFx4f_ASAP7_75t_L g926 ( 
.A(n_757),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_729),
.B(n_317),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_800),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_716),
.B(n_610),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_716),
.B(n_700),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_799),
.B(n_243),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_727),
.B(n_743),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_696),
.B(n_663),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_679),
.A2(n_616),
.B(n_610),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_771),
.B(n_750),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_692),
.A2(n_616),
.B(n_610),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_740),
.A2(n_597),
.B(n_619),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_775),
.B(n_616),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_817),
.B(n_318),
.Y(n_939)
);

AO21x1_ASAP7_75t_L g940 ( 
.A1(n_686),
.A2(n_707),
.B(n_688),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_775),
.B(n_619),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_750),
.B(n_261),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_740),
.A2(n_594),
.B(n_632),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_669),
.A2(n_594),
.B(n_632),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_669),
.A2(n_594),
.B(n_632),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_685),
.B(n_320),
.Y(n_946)
);

AO21x1_ASAP7_75t_L g947 ( 
.A1(n_688),
.A2(n_448),
.B(n_443),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_748),
.B(n_626),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_768),
.Y(n_949)
);

BUFx12f_ASAP7_75t_L g950 ( 
.A(n_760),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_L g951 ( 
.A(n_660),
.B(n_275),
.C(n_266),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_682),
.A2(n_457),
.B(n_458),
.C(n_460),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_699),
.B(n_417),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_768),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_730),
.B(n_626),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_682),
.A2(n_457),
.B(n_458),
.C(n_460),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_788),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_751),
.B(n_812),
.C(n_789),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_730),
.B(n_626),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_L g960 ( 
.A(n_719),
.B(n_626),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_728),
.A2(n_632),
.B1(n_594),
.B2(n_272),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_790),
.A2(n_455),
.B(n_458),
.C(n_460),
.Y(n_962)
);

NAND2x2_ASAP7_75t_L g963 ( 
.A(n_678),
.B(n_270),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_788),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_731),
.A2(n_594),
.B(n_632),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_731),
.A2(n_582),
.B(n_430),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_801),
.A2(n_462),
.B(n_453),
.C(n_455),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_720),
.A2(n_325),
.B1(n_279),
.B2(n_327),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_791),
.B(n_492),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_791),
.B(n_492),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_746),
.A2(n_582),
.B(n_432),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_793),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_707),
.A2(n_448),
.B(n_443),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_794),
.B(n_280),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_746),
.A2(n_582),
.B(n_432),
.Y(n_975)
);

O2A1O1Ixp5_ASAP7_75t_L g976 ( 
.A1(n_711),
.A2(n_448),
.B(n_443),
.C(n_502),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_747),
.A2(n_462),
.B(n_455),
.C(n_453),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_814),
.Y(n_978)
);

AOI21xp33_ASAP7_75t_L g979 ( 
.A1(n_794),
.A2(n_296),
.B(n_291),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_818),
.B(n_298),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_778),
.A2(n_333),
.B1(n_301),
.B2(n_305),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_749),
.A2(n_582),
.B(n_438),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_676),
.A2(n_582),
.B(n_493),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_747),
.A2(n_462),
.B(n_453),
.C(n_502),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_795),
.B(n_493),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_676),
.A2(n_502),
.B(n_498),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_818),
.B(n_304),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_747),
.A2(n_265),
.B1(n_324),
.B2(n_495),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_796),
.B(n_493),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_810),
.A2(n_498),
.B(n_493),
.C(n_495),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_814),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_749),
.A2(n_432),
.B(n_426),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_810),
.B(n_421),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_810),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_719),
.B(n_265),
.Y(n_995)
);

CKINVDCx10_ASAP7_75t_R g996 ( 
.A(n_769),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_796),
.Y(n_997)
);

AND2x6_ASAP7_75t_L g998 ( 
.A(n_778),
.B(n_423),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_711),
.A2(n_437),
.B(n_432),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_813),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_761),
.A2(n_438),
.B(n_437),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_763),
.B(n_311),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_725),
.A2(n_438),
.B(n_430),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_736),
.A2(n_438),
.B(n_437),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_813),
.B(n_495),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_845),
.A2(n_739),
.B(n_785),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_933),
.A2(n_765),
.B(n_822),
.C(n_809),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_845),
.A2(n_804),
.B(n_783),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_915),
.B(n_953),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_844),
.B(n_823),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_962),
.A2(n_816),
.B(n_815),
.C(n_811),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_960),
.A2(n_807),
.B(n_805),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_828),
.A2(n_722),
.B1(n_726),
.B2(n_717),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_930),
.B(n_719),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_887),
.B(n_719),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_857),
.B(n_719),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_923),
.Y(n_1017)
);

O2A1O1Ixp5_ASAP7_75t_SL g1018 ( 
.A1(n_995),
.A2(n_717),
.B(n_803),
.C(n_797),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_926),
.B(n_719),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_841),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_850),
.B(n_770),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_967),
.A2(n_808),
.B(n_773),
.C(n_772),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_857),
.B(n_719),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_848),
.A2(n_808),
.B(n_498),
.C(n_495),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_926),
.B(n_814),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_872),
.A2(n_781),
.B(n_498),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_994),
.B(n_324),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1002),
.A2(n_324),
.B1(n_461),
.B2(n_459),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_865),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_843),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_955),
.A2(n_312),
.B1(n_316),
.B2(n_329),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_974),
.A2(n_330),
.B(n_331),
.C(n_461),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_980),
.B(n_461),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_832),
.A2(n_426),
.B(n_430),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_949),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_832),
.A2(n_863),
.B(n_858),
.Y(n_1036)
);

OAI21xp33_ASAP7_75t_SL g1037 ( 
.A1(n_852),
.A2(n_461),
.B(n_459),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_977),
.A2(n_459),
.B(n_452),
.C(n_430),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_954),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_870),
.B(n_324),
.Y(n_1040)
);

AND2x2_ASAP7_75t_SL g1041 ( 
.A(n_935),
.B(n_452),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_830),
.A2(n_426),
.B(n_437),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_830),
.A2(n_897),
.B(n_904),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_897),
.A2(n_426),
.B(n_444),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_L g1045 ( 
.A(n_942),
.B(n_452),
.C(n_459),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_916),
.B(n_452),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_928),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_959),
.A2(n_644),
.B1(n_456),
.B2(n_444),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_874),
.B(n_440),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_987),
.B(n_456),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_873),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_846),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_880),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_882),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_825),
.A2(n_440),
.B(n_441),
.C(n_444),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_902),
.A2(n_444),
.B(n_441),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_894),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_958),
.A2(n_440),
.B(n_441),
.C(n_444),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_979),
.A2(n_878),
.B(n_871),
.C(n_931),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_829),
.B(n_456),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_993),
.B(n_456),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_903),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_923),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_919),
.Y(n_1064)
);

NOR2x1_ASAP7_75t_L g1065 ( 
.A(n_910),
.B(n_441),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_831),
.A2(n_833),
.B1(n_908),
.B2(n_837),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_993),
.B(n_456),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_L g1068 ( 
.A(n_998),
.B(n_856),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_905),
.B(n_19),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_918),
.A2(n_441),
.B(n_444),
.C(n_456),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_911),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_946),
.A2(n_441),
.B(n_24),
.C(n_25),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_916),
.B(n_456),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_927),
.B(n_24),
.Y(n_1074)
);

OAI21xp33_ASAP7_75t_SL g1075 ( 
.A1(n_847),
.A2(n_864),
.B(n_839),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_981),
.B(n_26),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_856),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_951),
.A2(n_456),
.B1(n_644),
.B2(n_68),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_856),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_849),
.B(n_27),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_855),
.A2(n_456),
.B1(n_644),
.B2(n_76),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_826),
.B(n_456),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_851),
.B(n_28),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_SL g1084 ( 
.A1(n_920),
.A2(n_66),
.B(n_168),
.C(n_161),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_923),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_957),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_860),
.B(n_861),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_917),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_881),
.B(n_29),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_875),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_824),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_952),
.A2(n_30),
.B(n_35),
.C(n_37),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_964),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_855),
.B(n_644),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_902),
.A2(n_79),
.B(n_158),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_889),
.B(n_30),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_910),
.B(n_65),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_950),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_996),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_913),
.A2(n_102),
.B(n_156),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_932),
.A2(n_160),
.B1(n_154),
.B2(n_151),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_896),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_917),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_963),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_888),
.B(n_150),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_991),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_913),
.A2(n_133),
.B(n_141),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_888),
.B(n_147),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_972),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_908),
.A2(n_138),
.B1(n_135),
.B2(n_127),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_888),
.B(n_125),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_827),
.A2(n_42),
.B(n_43),
.C(n_45),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_898),
.A2(n_120),
.B(n_46),
.Y(n_1113)
);

INVx3_ASAP7_75t_SL g1114 ( 
.A(n_866),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_968),
.B(n_43),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1000),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_924),
.A2(n_48),
.B(n_49),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_956),
.A2(n_50),
.B(n_55),
.C(n_56),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_834),
.Y(n_1119)
);

BUFx8_ASAP7_75t_L g1120 ( 
.A(n_998),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_876),
.A2(n_886),
.B(n_907),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_997),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_SL g1123 ( 
.A(n_988),
.B(n_55),
.C(n_56),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_834),
.B(n_57),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_969),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_970),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_991),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_984),
.A2(n_60),
.B(n_853),
.C(n_869),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_L g1129 ( 
.A(n_842),
.B(n_978),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_842),
.B(n_901),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_892),
.B(n_899),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_921),
.A2(n_922),
.B(n_859),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_874),
.B(n_991),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_877),
.A2(n_838),
.B(n_936),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_978),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_868),
.A2(n_990),
.B(n_900),
.C(n_895),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_940),
.A2(n_929),
.B(n_989),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_939),
.B(n_867),
.Y(n_1138)
);

BUFx12f_ASAP7_75t_L g1139 ( 
.A(n_998),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_985),
.A2(n_1005),
.B(n_941),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_891),
.A2(n_938),
.B1(n_906),
.B2(n_912),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_R g1142 ( 
.A(n_998),
.B(n_948),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_884),
.A2(n_879),
.B(n_961),
.C(n_909),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_885),
.A2(n_976),
.B(n_937),
.C(n_890),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_925),
.B(n_973),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_893),
.A2(n_936),
.B(n_934),
.Y(n_1146)
);

INVx4_ASAP7_75t_L g1147 ( 
.A(n_998),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1001),
.Y(n_1148)
);

OAI21xp33_ASAP7_75t_L g1149 ( 
.A1(n_986),
.A2(n_934),
.B(n_1001),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_947),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_965),
.B(n_943),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_SL g1152 ( 
.A(n_965),
.B(n_943),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_914),
.A2(n_883),
.B1(n_893),
.B2(n_944),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_914),
.A2(n_945),
.B(n_983),
.C(n_975),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_883),
.A2(n_835),
.B1(n_854),
.B2(n_862),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_971),
.B(n_982),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_835),
.A2(n_836),
.B1(n_840),
.B2(n_966),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_966),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_992),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_836),
.B(n_840),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_971),
.A2(n_975),
.B(n_982),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1087),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1009),
.B(n_1004),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1044),
.A2(n_1004),
.B(n_992),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1047),
.B(n_999),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1044),
.A2(n_1003),
.B(n_999),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1007),
.A2(n_1041),
.B1(n_1013),
.B2(n_1010),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1021),
.B(n_1126),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1115),
.A2(n_1069),
.B1(n_1076),
.B2(n_1074),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1030),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1035),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1135),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1125),
.B(n_1131),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1042),
.A2(n_1146),
.B(n_1034),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1043),
.A2(n_1157),
.A3(n_1145),
.B(n_1036),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1039),
.B(n_1093),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_1016),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1043),
.A2(n_1036),
.A3(n_1146),
.B(n_1153),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1017),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1042),
.A2(n_1034),
.B(n_1161),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_1134),
.A2(n_1137),
.B(n_1149),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1122),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1132),
.A2(n_1121),
.B(n_1026),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1132),
.A2(n_1121),
.B(n_1006),
.Y(n_1184)
);

OAI21xp33_ASAP7_75t_L g1185 ( 
.A1(n_1080),
.A2(n_1040),
.B(n_1123),
.Y(n_1185)
);

INVx5_ASAP7_75t_L g1186 ( 
.A(n_1017),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1160),
.A2(n_1050),
.B(n_1033),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1031),
.A2(n_1092),
.B1(n_1102),
.B2(n_1118),
.C(n_1112),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_1139),
.B(n_1088),
.Y(n_1189)
);

AOI222xp33_ASAP7_75t_L g1190 ( 
.A1(n_1027),
.A2(n_1089),
.B1(n_1096),
.B2(n_1083),
.C1(n_1114),
.C2(n_1053),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1128),
.A2(n_1032),
.B(n_1072),
.C(n_1143),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1128),
.A2(n_1138),
.B(n_1075),
.C(n_1028),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1020),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1092),
.A2(n_1117),
.B(n_1124),
.C(n_1084),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1155),
.A2(n_1008),
.B(n_1015),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1008),
.A2(n_1006),
.B(n_1014),
.Y(n_1196)
);

INVx5_ASAP7_75t_L g1197 ( 
.A(n_1017),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1140),
.A2(n_1137),
.B(n_1056),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_SL g1199 ( 
.A1(n_1101),
.A2(n_1078),
.B(n_1117),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1091),
.Y(n_1200)
);

INVxp67_ASAP7_75t_SL g1201 ( 
.A(n_1023),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1029),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1025),
.A2(n_1066),
.B(n_1104),
.C(n_1097),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1140),
.A2(n_1056),
.B(n_1151),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1158),
.A2(n_1012),
.B(n_1113),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1063),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1012),
.A2(n_1152),
.B(n_1144),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1136),
.A2(n_1156),
.B(n_1011),
.Y(n_1208)
);

INVx4_ASAP7_75t_L g1209 ( 
.A(n_1063),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1051),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1158),
.A2(n_1148),
.B(n_1018),
.Y(n_1211)
);

BUFx10_ASAP7_75t_L g1212 ( 
.A(n_1090),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1103),
.B(n_1067),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1063),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1085),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1055),
.A2(n_1038),
.B(n_1022),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1054),
.B(n_1109),
.Y(n_1217)
);

O2A1O1Ixp5_ASAP7_75t_L g1218 ( 
.A1(n_1154),
.A2(n_1141),
.B(n_1073),
.C(n_1019),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1057),
.B(n_1086),
.Y(n_1219)
);

OA22x2_ASAP7_75t_L g1220 ( 
.A1(n_1099),
.A2(n_1119),
.B1(n_1081),
.B2(n_1105),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1062),
.A2(n_1116),
.B1(n_1064),
.B2(n_1045),
.Y(n_1221)
);

NAND2x1p5_ASAP7_75t_L g1222 ( 
.A(n_1079),
.B(n_1147),
.Y(n_1222)
);

AOI21xp33_ASAP7_75t_L g1223 ( 
.A1(n_1011),
.A2(n_1022),
.B(n_1037),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1130),
.B(n_1150),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1079),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1055),
.A2(n_1038),
.B(n_1082),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_SL g1227 ( 
.A1(n_1108),
.A2(n_1111),
.B(n_1094),
.C(n_1133),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1095),
.A2(n_1100),
.B(n_1107),
.C(n_1061),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1052),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1147),
.A2(n_1060),
.B1(n_1046),
.B2(n_1159),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1095),
.A2(n_1100),
.B(n_1107),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_1085),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1068),
.A2(n_1159),
.B(n_1070),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1077),
.B(n_1071),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1098),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1085),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1058),
.Y(n_1237)
);

AO21x2_ASAP7_75t_L g1238 ( 
.A1(n_1142),
.A2(n_1024),
.B(n_1048),
.Y(n_1238)
);

BUFx4_ASAP7_75t_SL g1239 ( 
.A(n_1120),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1049),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1110),
.A2(n_1024),
.A3(n_1159),
.B(n_1065),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1106),
.B(n_1127),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1129),
.A2(n_1049),
.B(n_1120),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1106),
.A2(n_525),
.B(n_511),
.C(n_714),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1106),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1127),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1127),
.B(n_880),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1036),
.A2(n_1137),
.B(n_845),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1134),
.A2(n_1043),
.B(n_1146),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1043),
.A2(n_533),
.B(n_960),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1043),
.A2(n_1157),
.A3(n_1145),
.B(n_1036),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1059),
.A2(n_511),
.B(n_933),
.C(n_714),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1044),
.A2(n_898),
.B(n_1042),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1036),
.A2(n_1137),
.B(n_845),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1043),
.A2(n_533),
.B(n_960),
.Y(n_1255)
);

OA21x2_ASAP7_75t_L g1256 ( 
.A1(n_1134),
.A2(n_1043),
.B(n_1146),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1030),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1087),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1043),
.A2(n_1157),
.A3(n_1145),
.B(n_1036),
.Y(n_1259)
);

INVx4_ASAP7_75t_L g1260 ( 
.A(n_1017),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1044),
.A2(n_898),
.B(n_1042),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1044),
.A2(n_898),
.B(n_1042),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1059),
.A2(n_525),
.B(n_511),
.C(n_714),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1059),
.A2(n_511),
.B(n_933),
.C(n_714),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1059),
.A2(n_511),
.B(n_933),
.C(n_714),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1043),
.A2(n_1157),
.A3(n_1145),
.B(n_1036),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1044),
.A2(n_898),
.B(n_1042),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1009),
.B(n_695),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1009),
.B(n_706),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1043),
.A2(n_533),
.B(n_960),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1009),
.A2(n_689),
.B1(n_535),
.B2(n_525),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1087),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1087),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1044),
.A2(n_898),
.B(n_1042),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1009),
.B(n_828),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1103),
.Y(n_1276)
);

AND3x2_ASAP7_75t_L g1277 ( 
.A(n_1115),
.B(n_685),
.C(n_771),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1009),
.B(n_706),
.Y(n_1278)
);

BUFx12f_ASAP7_75t_L g1279 ( 
.A(n_1090),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1122),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_SL g1281 ( 
.A1(n_1128),
.A2(n_1117),
.B(n_1118),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1009),
.B(n_708),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1052),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1091),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1087),
.Y(n_1285)
);

AO21x2_ASAP7_75t_L g1286 ( 
.A1(n_1043),
.A2(n_1134),
.B(n_1036),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1009),
.B(n_584),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1087),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1017),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1009),
.B(n_706),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1043),
.A2(n_533),
.B(n_960),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1044),
.A2(n_898),
.B(n_1042),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1059),
.A2(n_511),
.B(n_933),
.C(n_714),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1009),
.B(n_933),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1043),
.A2(n_533),
.B(n_960),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1009),
.B(n_708),
.Y(n_1296)
);

OAI22x1_ASAP7_75t_L g1297 ( 
.A1(n_1080),
.A2(n_702),
.B1(n_933),
.B2(n_663),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1059),
.B(n_511),
.C(n_714),
.Y(n_1298)
);

AOI221x1_ASAP7_75t_L g1299 ( 
.A1(n_1112),
.A2(n_1043),
.B1(n_1146),
.B2(n_660),
.C(n_1117),
.Y(n_1299)
);

O2A1O1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1059),
.A2(n_525),
.B(n_511),
.C(n_714),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1009),
.A2(n_689),
.B1(n_535),
.B2(n_525),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1043),
.A2(n_533),
.B(n_960),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1122),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1044),
.A2(n_898),
.B(n_1042),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1043),
.A2(n_1157),
.A3(n_1145),
.B(n_1036),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1009),
.B(n_708),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1135),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1009),
.B(n_584),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1044),
.A2(n_898),
.B(n_1042),
.Y(n_1309)
);

AO21x1_ASAP7_75t_L g1310 ( 
.A1(n_1059),
.A2(n_1128),
.B(n_1117),
.Y(n_1310)
);

NOR2x1_ASAP7_75t_SL g1311 ( 
.A(n_1139),
.B(n_1147),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1043),
.A2(n_533),
.B(n_960),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1043),
.A2(n_533),
.B(n_960),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1169),
.A2(n_1297),
.B1(n_1185),
.B2(n_1298),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1294),
.A2(n_1298),
.B1(n_1167),
.B2(n_1271),
.Y(n_1315)
);

INVx4_ASAP7_75t_L g1316 ( 
.A(n_1186),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1257),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1283),
.Y(n_1318)
);

BUFx8_ASAP7_75t_L g1319 ( 
.A(n_1279),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1169),
.A2(n_1287),
.B1(n_1308),
.B2(n_1168),
.Y(n_1320)
);

BUFx12f_ASAP7_75t_L g1321 ( 
.A(n_1235),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_1200),
.Y(n_1322)
);

CKINVDCx6p67_ASAP7_75t_R g1323 ( 
.A(n_1229),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1268),
.B(n_1162),
.Y(n_1324)
);

CKINVDCx8_ASAP7_75t_R g1325 ( 
.A(n_1284),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1247),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1185),
.A2(n_1188),
.B1(n_1190),
.B2(n_1301),
.Y(n_1327)
);

CKINVDCx11_ASAP7_75t_R g1328 ( 
.A(n_1212),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1190),
.A2(n_1301),
.B1(n_1271),
.B2(n_1310),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1167),
.A2(n_1208),
.B1(n_1281),
.B2(n_1220),
.Y(n_1330)
);

BUFx4f_ASAP7_75t_L g1331 ( 
.A(n_1189),
.Y(n_1331)
);

CKINVDCx11_ASAP7_75t_R g1332 ( 
.A(n_1212),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1186),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1170),
.Y(n_1334)
);

BUFx2_ASAP7_75t_SL g1335 ( 
.A(n_1197),
.Y(n_1335)
);

INVx4_ASAP7_75t_SL g1336 ( 
.A(n_1179),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1171),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1275),
.A2(n_1277),
.B1(n_1165),
.B2(n_1208),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1252),
.A2(n_1265),
.B(n_1264),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1269),
.A2(n_1278),
.B1(n_1290),
.B2(n_1273),
.Y(n_1340)
);

BUFx2_ASAP7_75t_SL g1341 ( 
.A(n_1197),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1182),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1269),
.A2(n_1290),
.B1(n_1278),
.B2(n_1272),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1276),
.Y(n_1344)
);

CKINVDCx6p67_ASAP7_75t_R g1345 ( 
.A(n_1197),
.Y(n_1345)
);

CKINVDCx11_ASAP7_75t_R g1346 ( 
.A(n_1189),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1258),
.A2(n_1285),
.B1(n_1288),
.B2(n_1168),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1280),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1237),
.A2(n_1163),
.B1(n_1223),
.B2(n_1173),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1249),
.A2(n_1256),
.B1(n_1181),
.B2(n_1286),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1250),
.A2(n_1313),
.B(n_1312),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1249),
.A2(n_1256),
.B1(n_1181),
.B2(n_1286),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1234),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1263),
.A2(n_1300),
.B1(n_1306),
.B2(n_1282),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1296),
.B(n_1173),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1163),
.A2(n_1223),
.B1(n_1224),
.B2(n_1303),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1224),
.A2(n_1210),
.B1(n_1202),
.B2(n_1193),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1207),
.A2(n_1254),
.B1(n_1248),
.B2(n_1177),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1248),
.A2(n_1254),
.B1(n_1201),
.B2(n_1219),
.Y(n_1359)
);

CKINVDCx6p67_ASAP7_75t_R g1360 ( 
.A(n_1189),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1217),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1199),
.A2(n_1192),
.B1(n_1244),
.B2(n_1191),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1172),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1247),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1213),
.B(n_1221),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1213),
.A2(n_1216),
.B1(n_1238),
.B2(n_1231),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1199),
.A2(n_1221),
.B1(n_1230),
.B2(n_1233),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1232),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1239),
.Y(n_1369)
);

BUFx8_ASAP7_75t_L g1370 ( 
.A(n_1206),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1206),
.Y(n_1371)
);

CKINVDCx16_ASAP7_75t_R g1372 ( 
.A(n_1209),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1245),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1203),
.B(n_1307),
.Y(n_1374)
);

INVx8_ASAP7_75t_L g1375 ( 
.A(n_1215),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1243),
.A2(n_1242),
.B1(n_1214),
.B2(n_1209),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1215),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1215),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1299),
.B(n_1246),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1246),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1236),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1230),
.A2(n_1194),
.B1(n_1228),
.B2(n_1222),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1236),
.Y(n_1383)
);

CKINVDCx6p67_ASAP7_75t_R g1384 ( 
.A(n_1236),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1238),
.A2(n_1195),
.B1(n_1196),
.B2(n_1180),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1187),
.A2(n_1243),
.B1(n_1240),
.B2(n_1226),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1289),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1222),
.A2(n_1295),
.B1(n_1255),
.B2(n_1302),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1311),
.A2(n_1270),
.B1(n_1291),
.B2(n_1184),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1289),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1175),
.B(n_1266),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1225),
.A2(n_1227),
.B(n_1218),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1175),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1225),
.A2(n_1260),
.B1(n_1214),
.B2(n_1204),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1260),
.Y(n_1395)
);

CKINVDCx11_ASAP7_75t_R g1396 ( 
.A(n_1241),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1198),
.A2(n_1174),
.B1(n_1183),
.B2(n_1211),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1205),
.A2(n_1164),
.B1(n_1166),
.B2(n_1309),
.Y(n_1398)
);

INVx8_ASAP7_75t_L g1399 ( 
.A(n_1241),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1251),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1253),
.A2(n_1267),
.B1(n_1304),
.B2(n_1292),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1259),
.B(n_1305),
.Y(n_1402)
);

BUFx8_ASAP7_75t_L g1403 ( 
.A(n_1266),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_SL g1404 ( 
.A1(n_1305),
.A2(n_1178),
.B1(n_1261),
.B2(n_1262),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1178),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1274),
.A2(n_1169),
.B1(n_1297),
.B2(n_771),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1250),
.A2(n_1270),
.B(n_1255),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1294),
.B(n_1287),
.Y(n_1408)
);

INVx6_ASAP7_75t_L g1409 ( 
.A(n_1186),
.Y(n_1409)
);

OAI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1169),
.A2(n_1297),
.B1(n_771),
.B2(n_1298),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1294),
.A2(n_771),
.B1(n_504),
.B2(n_600),
.Y(n_1411)
);

BUFx2_ASAP7_75t_SL g1412 ( 
.A(n_1257),
.Y(n_1412)
);

CKINVDCx6p67_ASAP7_75t_R g1413 ( 
.A(n_1283),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1294),
.A2(n_771),
.B1(n_504),
.B2(n_600),
.Y(n_1414)
);

INVx6_ASAP7_75t_L g1415 ( 
.A(n_1186),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1257),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1175),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1169),
.A2(n_933),
.B1(n_696),
.B2(n_1297),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1294),
.B(n_1287),
.Y(n_1419)
);

CKINVDCx11_ASAP7_75t_R g1420 ( 
.A(n_1235),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1294),
.A2(n_771),
.B1(n_504),
.B2(n_600),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1294),
.A2(n_771),
.B1(n_504),
.B2(n_600),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1169),
.A2(n_1293),
.B1(n_1252),
.B2(n_1265),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1176),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1169),
.A2(n_1297),
.B1(n_1185),
.B2(n_1298),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1169),
.A2(n_1293),
.B1(n_1252),
.B2(n_1265),
.Y(n_1426)
);

BUFx2_ASAP7_75t_SL g1427 ( 
.A(n_1257),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1212),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1169),
.A2(n_1293),
.B1(n_1252),
.B2(n_1265),
.Y(n_1429)
);

INVx11_ASAP7_75t_L g1430 ( 
.A(n_1279),
.Y(n_1430)
);

BUFx8_ASAP7_75t_SL g1431 ( 
.A(n_1279),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1176),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1351),
.A2(n_1407),
.B(n_1397),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1393),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1315),
.B(n_1400),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1408),
.B(n_1419),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1417),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1351),
.A2(n_1407),
.B(n_1339),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1397),
.A2(n_1401),
.B(n_1385),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1315),
.B(n_1329),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1417),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1405),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1385),
.A2(n_1391),
.B(n_1329),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1402),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1314),
.B(n_1425),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1403),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1320),
.B(n_1340),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1403),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1379),
.B(n_1314),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1320),
.B(n_1340),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1399),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1365),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1358),
.A2(n_1401),
.B(n_1356),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1388),
.A2(n_1398),
.B(n_1382),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1404),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1396),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1366),
.A2(n_1386),
.B(n_1358),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1337),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1330),
.B(n_1356),
.Y(n_1459)
);

INVxp33_ASAP7_75t_L g1460 ( 
.A(n_1416),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1342),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1359),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1359),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1374),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1424),
.Y(n_1465)
);

OR2x6_ASAP7_75t_L g1466 ( 
.A(n_1362),
.B(n_1367),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1432),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1361),
.Y(n_1468)
);

INVx1_ASAP7_75t_SL g1469 ( 
.A(n_1373),
.Y(n_1469)
);

AO21x1_ASAP7_75t_L g1470 ( 
.A1(n_1423),
.A2(n_1429),
.B(n_1426),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1350),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1350),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1412),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1330),
.B(n_1327),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1348),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1343),
.B(n_1347),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1406),
.A2(n_1410),
.B(n_1392),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1352),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1331),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1352),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1349),
.A2(n_1366),
.B(n_1386),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1349),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1324),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1389),
.A2(n_1410),
.B(n_1406),
.Y(n_1484)
);

AO21x2_ASAP7_75t_L g1485 ( 
.A1(n_1418),
.A2(n_1389),
.B(n_1355),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1363),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1331),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1368),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1357),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1394),
.A2(n_1357),
.B(n_1343),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1347),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1327),
.A2(n_1380),
.B(n_1383),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1338),
.A2(n_1381),
.B(n_1354),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1354),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1411),
.B(n_1414),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1322),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1409),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1334),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1427),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1376),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1378),
.A2(n_1387),
.B(n_1395),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1353),
.B(n_1325),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1360),
.A2(n_1336),
.B(n_1335),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1364),
.A2(n_1428),
.B(n_1414),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1341),
.A2(n_1346),
.B(n_1345),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1318),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1415),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1415),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1316),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1411),
.B(n_1422),
.Y(n_1510)
);

AO21x2_ASAP7_75t_L g1511 ( 
.A1(n_1421),
.A2(n_1422),
.B(n_1384),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1421),
.B(n_1326),
.Y(n_1512)
);

CKINVDCx6p67_ASAP7_75t_R g1513 ( 
.A(n_1420),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1333),
.Y(n_1514)
);

AOI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1495),
.A2(n_1317),
.B1(n_1372),
.B2(n_1369),
.C(n_1371),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1470),
.B(n_1326),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1436),
.B(n_1460),
.Y(n_1517)
);

NOR2x1_ASAP7_75t_SL g1518 ( 
.A(n_1466),
.B(n_1321),
.Y(n_1518)
);

NAND2x1p5_ASAP7_75t_L g1519 ( 
.A(n_1501),
.B(n_1377),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1452),
.B(n_1413),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1464),
.B(n_1323),
.Y(n_1521)
);

OR2x6_ASAP7_75t_L g1522 ( 
.A(n_1484),
.B(n_1466),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1484),
.A2(n_1370),
.B(n_1375),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1501),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1439),
.A2(n_1370),
.B(n_1375),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1439),
.A2(n_1390),
.B(n_1328),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1451),
.B(n_1332),
.Y(n_1527)
);

OAI211xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1495),
.A2(n_1344),
.B(n_1319),
.C(n_1431),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_SL g1529 ( 
.A1(n_1470),
.A2(n_1319),
.B(n_1430),
.Y(n_1529)
);

OR2x6_ASAP7_75t_L g1530 ( 
.A(n_1466),
.B(n_1454),
.Y(n_1530)
);

O2A1O1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1510),
.A2(n_1494),
.B(n_1466),
.C(n_1447),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1466),
.A2(n_1440),
.B1(n_1474),
.B2(n_1510),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1491),
.B(n_1482),
.Y(n_1533)
);

A2O1A1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1440),
.A2(n_1474),
.B(n_1459),
.C(n_1445),
.Y(n_1534)
);

AO32x2_ASAP7_75t_L g1535 ( 
.A1(n_1449),
.A2(n_1444),
.A3(n_1480),
.B1(n_1471),
.B2(n_1472),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1512),
.B(n_1435),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1512),
.B(n_1435),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1483),
.B(n_1504),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1459),
.A2(n_1494),
.B1(n_1447),
.B2(n_1450),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1504),
.B(n_1456),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1498),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1450),
.A2(n_1445),
.B(n_1490),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1504),
.B(n_1456),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1504),
.B(n_1456),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1511),
.B(n_1449),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1491),
.B(n_1482),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1456),
.B(n_1446),
.Y(n_1547)
);

AOI221xp5_ASAP7_75t_L g1548 ( 
.A1(n_1476),
.A2(n_1463),
.B1(n_1462),
.B2(n_1489),
.C(n_1511),
.Y(n_1548)
);

NAND2xp33_ASAP7_75t_R g1549 ( 
.A(n_1448),
.B(n_1496),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1458),
.B(n_1462),
.Y(n_1550)
);

AO32x2_ASAP7_75t_L g1551 ( 
.A1(n_1478),
.A2(n_1443),
.A3(n_1501),
.B1(n_1485),
.B2(n_1477),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1463),
.B(n_1461),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1475),
.B(n_1489),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1434),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1448),
.B(n_1485),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1498),
.Y(n_1556)
);

NAND2x1_ASAP7_75t_L g1557 ( 
.A(n_1501),
.B(n_1509),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1485),
.B(n_1488),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1511),
.B(n_1476),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1490),
.A2(n_1457),
.B(n_1454),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1493),
.B(n_1469),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1465),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1511),
.A2(n_1500),
.B(n_1469),
.C(n_1477),
.Y(n_1563)
);

O2A1O1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1500),
.A2(n_1477),
.B(n_1473),
.C(n_1499),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1465),
.A2(n_1467),
.B1(n_1468),
.B2(n_1479),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1493),
.A2(n_1438),
.B(n_1433),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1437),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1493),
.B(n_1486),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1467),
.B(n_1468),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1479),
.A2(n_1487),
.B1(n_1481),
.B2(n_1455),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1477),
.A2(n_1492),
.B(n_1507),
.C(n_1508),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1524),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1560),
.B(n_1438),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1522),
.A2(n_1539),
.B1(n_1559),
.B2(n_1545),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1560),
.B(n_1438),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1554),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1567),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1567),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1516),
.B(n_1497),
.Y(n_1579)
);

INVx3_ASAP7_75t_SL g1580 ( 
.A(n_1523),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1568),
.B(n_1540),
.Y(n_1581)
);

BUFx12f_ASAP7_75t_L g1582 ( 
.A(n_1520),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1543),
.B(n_1481),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1557),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1544),
.B(n_1481),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1524),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1538),
.B(n_1441),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1558),
.B(n_1442),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1569),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1566),
.B(n_1551),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1559),
.B(n_1443),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1553),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1545),
.B(n_1443),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1548),
.B(n_1443),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1551),
.B(n_1453),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1550),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1552),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1541),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1530),
.B(n_1453),
.Y(n_1599)
);

AND2x4_ASAP7_75t_SL g1600 ( 
.A(n_1530),
.B(n_1487),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1519),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1555),
.B(n_1453),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1581),
.B(n_1526),
.Y(n_1603)
);

OAI211xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1574),
.A2(n_1563),
.B(n_1548),
.C(n_1564),
.Y(n_1604)
);

NOR3xp33_ASAP7_75t_L g1605 ( 
.A(n_1594),
.B(n_1563),
.C(n_1528),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1582),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1591),
.B(n_1561),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1581),
.B(n_1526),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1577),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1577),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1578),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1591),
.B(n_1542),
.Y(n_1612)
);

OAI33xp33_ASAP7_75t_L g1613 ( 
.A1(n_1594),
.A2(n_1539),
.A3(n_1564),
.B1(n_1531),
.B2(n_1533),
.B3(n_1546),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1588),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1581),
.B(n_1535),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1572),
.Y(n_1616)
);

INVx4_ASAP7_75t_L g1617 ( 
.A(n_1582),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1587),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1593),
.B(n_1570),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1602),
.B(n_1535),
.Y(n_1620)
);

OAI31xp33_ASAP7_75t_L g1621 ( 
.A1(n_1574),
.A2(n_1534),
.A3(n_1531),
.B(n_1528),
.Y(n_1621)
);

OAI33xp33_ASAP7_75t_L g1622 ( 
.A1(n_1593),
.A2(n_1533),
.A3(n_1546),
.B1(n_1570),
.B2(n_1565),
.B3(n_1562),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1602),
.B(n_1535),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1578),
.B(n_1596),
.Y(n_1624)
);

INVx4_ASAP7_75t_L g1625 ( 
.A(n_1582),
.Y(n_1625)
);

AO22x1_ASAP7_75t_L g1626 ( 
.A1(n_1579),
.A2(n_1527),
.B1(n_1542),
.B2(n_1536),
.Y(n_1626)
);

AOI221xp5_ASAP7_75t_L g1627 ( 
.A1(n_1590),
.A2(n_1532),
.B1(n_1537),
.B2(n_1515),
.C(n_1571),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1576),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1572),
.Y(n_1629)
);

INVx4_ASAP7_75t_L g1630 ( 
.A(n_1600),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1587),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1586),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1580),
.A2(n_1515),
.B1(n_1522),
.B2(n_1517),
.C(n_1521),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1602),
.B(n_1547),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1599),
.B(n_1525),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1590),
.A2(n_1571),
.B(n_1505),
.C(n_1573),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1598),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1601),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1599),
.B(n_1583),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1586),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1639),
.B(n_1590),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1639),
.B(n_1583),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1609),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1612),
.B(n_1589),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1603),
.B(n_1608),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1628),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1609),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1619),
.B(n_1588),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1619),
.B(n_1592),
.Y(n_1649)
);

INVx6_ASAP7_75t_L g1650 ( 
.A(n_1617),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1630),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1610),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1628),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1614),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1630),
.B(n_1584),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_SL g1656 ( 
.A(n_1621),
.B(n_1513),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1630),
.B(n_1584),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1612),
.B(n_1589),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1616),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1605),
.A2(n_1522),
.B1(n_1579),
.B2(n_1599),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1617),
.B(n_1513),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1610),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1617),
.B(n_1527),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1616),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1607),
.B(n_1597),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1607),
.B(n_1597),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1608),
.B(n_1585),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1638),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1620),
.B(n_1595),
.Y(n_1669)
);

NAND2xp33_ASAP7_75t_R g1670 ( 
.A(n_1638),
.B(n_1523),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1611),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1629),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1620),
.B(n_1597),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1611),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1618),
.B(n_1592),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1623),
.B(n_1595),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1646),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1661),
.B(n_1637),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1643),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1648),
.B(n_1624),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1646),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1646),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1643),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1651),
.B(n_1623),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1644),
.B(n_1605),
.Y(n_1685)
);

NOR4xp25_ASAP7_75t_L g1686 ( 
.A(n_1656),
.B(n_1604),
.C(n_1636),
.D(n_1627),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1653),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1647),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1653),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1651),
.B(n_1615),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1663),
.B(n_1617),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1641),
.B(n_1615),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1647),
.Y(n_1693)
);

AOI32xp33_ASAP7_75t_L g1694 ( 
.A1(n_1656),
.A2(n_1604),
.A3(n_1627),
.B1(n_1633),
.B2(n_1625),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1641),
.B(n_1635),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1650),
.B(n_1625),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1653),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1652),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1648),
.B(n_1624),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1644),
.B(n_1621),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1652),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1650),
.B(n_1625),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1658),
.B(n_1626),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1641),
.B(n_1635),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1654),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1658),
.B(n_1626),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1671),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1649),
.B(n_1634),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1671),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1674),
.Y(n_1710)
);

OR2x6_ASAP7_75t_L g1711 ( 
.A(n_1650),
.B(n_1625),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1655),
.B(n_1634),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1674),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1662),
.Y(n_1714)
);

NAND2x1_ASAP7_75t_L g1715 ( 
.A(n_1655),
.B(n_1657),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1650),
.B(n_1606),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1649),
.B(n_1618),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1662),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1660),
.B(n_1631),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1679),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1684),
.B(n_1655),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1708),
.B(n_1673),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1684),
.B(n_1655),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1685),
.B(n_1673),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1700),
.B(n_1665),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1690),
.B(n_1655),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1715),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1679),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1690),
.B(n_1657),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1683),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1712),
.B(n_1657),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1677),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1683),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1686),
.B(n_1665),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1688),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1712),
.B(n_1657),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1688),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1678),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1693),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1694),
.B(n_1633),
.C(n_1670),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1677),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1680),
.B(n_1659),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1681),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1692),
.B(n_1657),
.Y(n_1744)
);

AOI211x1_ASAP7_75t_L g1745 ( 
.A1(n_1703),
.A2(n_1676),
.B(n_1669),
.C(n_1645),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1693),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1694),
.B(n_1666),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1692),
.B(n_1711),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1706),
.B(n_1666),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1680),
.B(n_1659),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1716),
.B(n_1668),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1699),
.B(n_1664),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1699),
.B(n_1664),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1698),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1681),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1724),
.B(n_1717),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1740),
.A2(n_1696),
.B(n_1702),
.C(n_1719),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1734),
.A2(n_1613),
.B(n_1691),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1727),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1720),
.Y(n_1760)
);

OAI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1738),
.A2(n_1650),
.B1(n_1711),
.B2(n_1714),
.C(n_1718),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1720),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1724),
.B(n_1711),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1747),
.A2(n_1613),
.B1(n_1622),
.B2(n_1714),
.C(n_1718),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1738),
.A2(n_1711),
.B1(n_1622),
.B2(n_1715),
.Y(n_1765)
);

A2O1A1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1725),
.A2(n_1606),
.B(n_1573),
.C(n_1575),
.Y(n_1766)
);

OAI31xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1748),
.A2(n_1668),
.A3(n_1502),
.B(n_1704),
.Y(n_1767)
);

O2A1O1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1751),
.A2(n_1672),
.B(n_1606),
.C(n_1529),
.Y(n_1768)
);

AOI32xp33_ASAP7_75t_L g1769 ( 
.A1(n_1748),
.A2(n_1704),
.A3(n_1695),
.B1(n_1645),
.B2(n_1575),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1728),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1728),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1749),
.B(n_1695),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1722),
.B(n_1645),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1730),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1745),
.B(n_1698),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1730),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1745),
.B(n_1701),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1731),
.B(n_1642),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1731),
.B(n_1642),
.Y(n_1779)
);

OAI21xp33_ASAP7_75t_L g1780 ( 
.A1(n_1721),
.A2(n_1575),
.B(n_1573),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1733),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1760),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1758),
.B(n_1721),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1762),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1770),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1771),
.Y(n_1786)
);

OAI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1765),
.A2(n_1727),
.B1(n_1750),
.B2(n_1753),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1757),
.A2(n_1723),
.B1(n_1729),
.B2(n_1726),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1774),
.Y(n_1789)
);

NAND5xp2_ASAP7_75t_SL g1790 ( 
.A(n_1761),
.B(n_1723),
.C(n_1726),
.D(n_1729),
.E(n_1736),
.Y(n_1790)
);

AOI32xp33_ASAP7_75t_L g1791 ( 
.A1(n_1764),
.A2(n_1744),
.A3(n_1736),
.B1(n_1739),
.B2(n_1737),
.Y(n_1791)
);

INVxp67_ASAP7_75t_SL g1792 ( 
.A(n_1767),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1767),
.B(n_1744),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1759),
.B(n_1742),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1776),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1761),
.A2(n_1739),
.B1(n_1754),
.B2(n_1733),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1775),
.A2(n_1753),
.B1(n_1752),
.B2(n_1750),
.Y(n_1797)
);

INVxp67_ASAP7_75t_SL g1798 ( 
.A(n_1768),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1763),
.B(n_1742),
.Y(n_1799)
);

NAND2x1p5_ASAP7_75t_L g1800 ( 
.A(n_1781),
.B(n_1637),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1778),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1792),
.A2(n_1777),
.B1(n_1775),
.B2(n_1756),
.Y(n_1802)
);

AOI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1787),
.A2(n_1777),
.B1(n_1772),
.B2(n_1766),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1800),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1794),
.Y(n_1805)
);

AOI322xp5_ASAP7_75t_L g1806 ( 
.A1(n_1783),
.A2(n_1780),
.A3(n_1779),
.B1(n_1669),
.B2(n_1676),
.C1(n_1754),
.C2(n_1735),
.Y(n_1806)
);

O2A1O1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1790),
.A2(n_1798),
.B(n_1800),
.C(n_1797),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1791),
.B(n_1769),
.Y(n_1808)
);

AOI211x1_ASAP7_75t_L g1809 ( 
.A1(n_1793),
.A2(n_1735),
.B(n_1737),
.C(n_1746),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1801),
.B(n_1773),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1788),
.A2(n_1796),
.B1(n_1799),
.B2(n_1797),
.Y(n_1811)
);

OA22x2_ASAP7_75t_L g1812 ( 
.A1(n_1782),
.A2(n_1746),
.B1(n_1707),
.B2(n_1701),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1784),
.Y(n_1813)
);

XOR2x2_ASAP7_75t_L g1814 ( 
.A(n_1785),
.B(n_1637),
.Y(n_1814)
);

AOI21xp33_ASAP7_75t_L g1815 ( 
.A1(n_1807),
.A2(n_1789),
.B(n_1786),
.Y(n_1815)
);

NAND4xp25_ASAP7_75t_SL g1816 ( 
.A(n_1811),
.B(n_1795),
.C(n_1752),
.D(n_1722),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1804),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1812),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1803),
.A2(n_1741),
.B(n_1732),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1810),
.Y(n_1820)
);

NOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1813),
.B(n_1506),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1808),
.A2(n_1741),
.B(n_1732),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1814),
.Y(n_1823)
);

OAI22xp33_ASAP7_75t_SL g1824 ( 
.A1(n_1802),
.A2(n_1755),
.B1(n_1743),
.B2(n_1741),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_SL g1825 ( 
.A1(n_1815),
.A2(n_1805),
.B(n_1549),
.Y(n_1825)
);

AOI211x1_ASAP7_75t_SL g1826 ( 
.A1(n_1819),
.A2(n_1809),
.B(n_1755),
.C(n_1743),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1816),
.A2(n_1755),
.B1(n_1743),
.B2(n_1732),
.C(n_1806),
.Y(n_1827)
);

AOI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1824),
.A2(n_1556),
.B(n_1580),
.C(n_1479),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1822),
.A2(n_1709),
.B(n_1707),
.Y(n_1829)
);

AOI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1827),
.A2(n_1821),
.B1(n_1823),
.B2(n_1817),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1828),
.A2(n_1820),
.B1(n_1818),
.B2(n_1713),
.Y(n_1831)
);

AOI21xp33_ASAP7_75t_L g1832 ( 
.A1(n_1825),
.A2(n_1705),
.B(n_1709),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1829),
.Y(n_1833)
);

OAI321xp33_ASAP7_75t_L g1834 ( 
.A1(n_1826),
.A2(n_1713),
.A3(n_1710),
.B1(n_1705),
.B2(n_1479),
.C(n_1487),
.Y(n_1834)
);

NOR3xp33_ASAP7_75t_SL g1835 ( 
.A(n_1827),
.B(n_1710),
.C(n_1514),
.Y(n_1835)
);

NOR2x1_ASAP7_75t_L g1836 ( 
.A(n_1833),
.B(n_1682),
.Y(n_1836)
);

NOR2x1_ASAP7_75t_L g1837 ( 
.A(n_1834),
.B(n_1682),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1830),
.B(n_1672),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1831),
.A2(n_1697),
.B1(n_1687),
.B2(n_1689),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1832),
.B(n_1687),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_SL g1841 ( 
.A1(n_1838),
.A2(n_1835),
.B(n_1487),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1836),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1840),
.B(n_1837),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1842),
.Y(n_1844)
);

OAI22x1_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1843),
.B1(n_1841),
.B2(n_1697),
.Y(n_1845)
);

INVxp67_ASAP7_75t_SL g1846 ( 
.A(n_1845),
.Y(n_1846)
);

AOI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1845),
.A2(n_1839),
.B(n_1689),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1846),
.A2(n_1847),
.B1(n_1654),
.B2(n_1675),
.Y(n_1848)
);

CKINVDCx20_ASAP7_75t_R g1849 ( 
.A(n_1846),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1849),
.A2(n_1487),
.B1(n_1640),
.B2(n_1676),
.Y(n_1850)
);

INVxp67_ASAP7_75t_SL g1851 ( 
.A(n_1848),
.Y(n_1851)
);

OAI21xp33_ASAP7_75t_L g1852 ( 
.A1(n_1851),
.A2(n_1669),
.B(n_1667),
.Y(n_1852)
);

OAI21x1_ASAP7_75t_SL g1853 ( 
.A1(n_1852),
.A2(n_1850),
.B(n_1518),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1853),
.Y(n_1854)
);

OAI221xp5_ASAP7_75t_R g1855 ( 
.A1(n_1854),
.A2(n_1640),
.B1(n_1654),
.B2(n_1580),
.C(n_1632),
.Y(n_1855)
);

AOI211xp5_ASAP7_75t_L g1856 ( 
.A1(n_1855),
.A2(n_1487),
.B(n_1503),
.C(n_1580),
.Y(n_1856)
);


endmodule