module fake_jpeg_28121_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_7),
.B(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_27),
.B1(n_24),
.B2(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_21),
.B1(n_33),
.B2(n_27),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_39),
.B1(n_38),
.B2(n_36),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_33),
.B1(n_21),
.B2(n_20),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_42),
.B1(n_39),
.B2(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_41),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_33),
.B1(n_27),
.B2(n_24),
.Y(n_51)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_20),
.B1(n_24),
.B2(n_29),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_30),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_40),
.B(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_28),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_63),
.C(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_88),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_40),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_64),
.B(n_68),
.Y(n_114)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_66),
.A2(n_56),
.B(n_58),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_30),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_80),
.B1(n_57),
.B2(n_58),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_30),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_32),
.B1(n_25),
.B2(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_25),
.B1(n_32),
.B2(n_37),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_37),
.B1(n_17),
.B2(n_18),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_23),
.B1(n_29),
.B2(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_43),
.B(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_83),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_55),
.B(n_17),
.CI(n_26),
.CON(n_83),
.SN(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_29),
.B1(n_23),
.B2(n_18),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_78),
.B1(n_64),
.B2(n_87),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_49),
.B(n_18),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_22),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_56),
.Y(n_97)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_93),
.A2(n_97),
.B(n_63),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_62),
.B1(n_76),
.B2(n_65),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_118),
.B1(n_44),
.B2(n_48),
.Y(n_135)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_113),
.Y(n_125)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_111),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_22),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_119),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_86),
.B1(n_68),
.B2(n_73),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_94),
.B1(n_93),
.B2(n_114),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_90),
.B1(n_89),
.B2(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_52),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_63),
.B1(n_66),
.B2(n_83),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_124),
.A2(n_130),
.B1(n_134),
.B2(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_138),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_63),
.C(n_67),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_140),
.C(n_101),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_60),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_111),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_119),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_142),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_71),
.B(n_67),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_146),
.B(n_112),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_71),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_141),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_80),
.B1(n_70),
.B2(n_69),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_136),
.B1(n_145),
.B2(n_98),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_69),
.B1(n_52),
.B2(n_48),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_17),
.B(n_26),
.C(n_70),
.D(n_16),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_146),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_52),
.C(n_48),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_62),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_85),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_117),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_85),
.B1(n_29),
.B2(n_23),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_94),
.A2(n_17),
.B(n_30),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_104),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_149),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_155),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_154),
.Y(n_191)
);

NAND2x1_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_92),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_152),
.A2(n_161),
.B(n_165),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_92),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_102),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_139),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_159),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_166),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_108),
.B(n_102),
.C(n_107),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_122),
.B(n_137),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_170),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_98),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_180),
.C(n_140),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_178),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_174),
.A2(n_0),
.B(n_1),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_142),
.A2(n_98),
.B1(n_112),
.B2(n_26),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_126),
.B1(n_121),
.B2(n_167),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_16),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_147),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_23),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_26),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_184),
.A2(n_189),
.B1(n_192),
.B2(n_198),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_180),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_10),
.B(n_13),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_133),
.C(n_135),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_203),
.C(n_208),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_145),
.B1(n_133),
.B2(n_121),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_193),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_26),
.B1(n_16),
.B2(n_9),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_0),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_192),
.B1(n_186),
.B2(n_193),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_1),
.Y(n_201)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_7),
.C(n_14),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_170),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_207),
.Y(n_217)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_182),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_6),
.C(n_13),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_156),
.A2(n_162),
.B1(n_169),
.B2(n_168),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_209),
.A2(n_176),
.B1(n_152),
.B2(n_161),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_227),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_214),
.B(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_160),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_219),
.B(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_194),
.B(n_153),
.Y(n_220)
);

AOI22x1_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_157),
.B1(n_171),
.B2(n_150),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_187),
.B1(n_208),
.B2(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_226),
.Y(n_238)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_191),
.C(n_185),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_225),
.C(n_233),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_155),
.C(n_9),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_6),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_6),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_231),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_229)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_197),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_232),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_5),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_212),
.C(n_225),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_218),
.C(n_233),
.Y(n_254)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_242),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_206),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_183),
.B(n_199),
.Y(n_258)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_203),
.Y(n_259)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_251),
.Y(n_257)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_213),
.B(n_195),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_252),
.B(n_10),
.Y(n_267)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_238),
.B(n_221),
.CI(n_201),
.CON(n_253),
.SN(n_253)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_250),
.Y(n_278)
);

AOI32xp33_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_247),
.A3(n_249),
.B1(n_241),
.B2(n_218),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_248),
.B(n_251),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_258),
.B(n_247),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_234),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_189),
.C(n_228),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_264),
.C(n_237),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_200),
.B(n_227),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_262),
.A2(n_236),
.B(n_235),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_265),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_205),
.C(n_5),
.Y(n_264)
);

BUFx12_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_10),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_12),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_267),
.A2(n_244),
.B1(n_236),
.B2(n_243),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_272),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_271),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_235),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_275),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_237),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_280),
.C(n_254),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_240),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_278),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_263),
.B1(n_260),
.B2(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_274),
.B(n_256),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_284),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_287),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_272),
.B(n_253),
.CI(n_264),
.CON(n_288),
.SN(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_273),
.C(n_258),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_296),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_277),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_292),
.A2(n_283),
.B(n_285),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_295),
.A2(n_286),
.B1(n_290),
.B2(n_287),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_288),
.A2(n_265),
.B1(n_12),
.B2(n_15),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_12),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_300),
.Y(n_305)
);

OAI211xp5_ASAP7_75t_L g304 ( 
.A1(n_301),
.A2(n_302),
.B(n_303),
.C(n_298),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_265),
.B(n_3),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_299),
.B(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_295),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_293),
.Y(n_310)
);


endmodule