module fake_jpeg_1492_n_89 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_89);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_89;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_37),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_30),
.B1(n_31),
.B2(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_2),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_47),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_34),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_29),
.B(n_27),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_49),
.A2(n_29),
.B(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

AO21x2_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_26),
.B(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_56),
.C(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_3),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_6),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_52),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_7),
.B(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_74),
.C(n_59),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_17),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_65),
.B(n_59),
.Y(n_78)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_7),
.CI(n_8),
.CON(n_76),
.SN(n_76)
);

AOI322xp5_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_16),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_81),
.B(n_72),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_80),
.C(n_82),
.Y(n_83)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_74),
.C(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_83),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_76),
.B(n_81),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_77),
.B(n_66),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_88),
.Y(n_89)
);


endmodule