module fake_jpeg_7418_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_26),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_17),
.B1(n_22),
.B2(n_24),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_22),
.B1(n_17),
.B2(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_17),
.B1(n_22),
.B2(n_28),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_53),
.B1(n_39),
.B2(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_41),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_66),
.B(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_57),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_72),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_10),
.C(n_9),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_73),
.C(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_48),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_40),
.C(n_13),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_45),
.B1(n_56),
.B2(n_53),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_68),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_49),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.C(n_85),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_51),
.C(n_39),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_62),
.B1(n_65),
.B2(n_50),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_26),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_48),
.C(n_43),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_96),
.C(n_98),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_81),
.B1(n_12),
.B2(n_50),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_70),
.A3(n_69),
.B1(n_68),
.B2(n_63),
.C1(n_72),
.C2(n_9),
.Y(n_95)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_43),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_87),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_43),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_86),
.C(n_78),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_105),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_82),
.B(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_50),
.B1(n_89),
.B2(n_21),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_104),
.A2(n_14),
.B1(n_19),
.B2(n_96),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_36),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_12),
.B(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_0),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_104),
.Y(n_117)
);

AOI321xp33_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_19),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_114),
.B(n_116),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_0),
.Y(n_115)
);

AOI31xp67_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_19),
.A3(n_46),
.B(n_36),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_106),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_114),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_112),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_107),
.B(n_121),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_126),
.A3(n_108),
.B1(n_14),
.B2(n_46),
.C1(n_6),
.C2(n_7),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_108),
.A3(n_101),
.B1(n_100),
.B2(n_105),
.C1(n_1),
.C2(n_7),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

AOI221xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_123),
.B1(n_6),
.B2(n_7),
.C(n_3),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_131),
.B(n_3),
.Y(n_134)
);


endmodule