module fake_jpeg_5008_n_137 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_24),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

NOR3xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_29),
.C(n_12),
.Y(n_34)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_15),
.Y(n_36)
);

BUFx2_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_13),
.Y(n_40)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_16),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_16),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_14),
.Y(n_50)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_50),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_31),
.B1(n_24),
.B2(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_38),
.Y(n_58)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_29),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_29),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_45),
.B1(n_32),
.B2(n_50),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_67),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_37),
.C(n_33),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_45),
.B(n_53),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_64),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_78),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_57),
.B1(n_31),
.B2(n_51),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_31),
.B1(n_43),
.B2(n_30),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_59),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_12),
.B(n_17),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_79),
.A2(n_18),
.B(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_76),
.B(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_89),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_88),
.B1(n_91),
.B2(n_77),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_56),
.B1(n_30),
.B2(n_46),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_26),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_18),
.B1(n_11),
.B2(n_13),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_72),
.B1(n_22),
.B2(n_26),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_20),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_98),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_101),
.B1(n_93),
.B2(n_99),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_68),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_68),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_102),
.B(n_92),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_20),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_107),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_84),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_106),
.Y(n_116)
);

OA21x2_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_84),
.B(n_20),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_111),
.B(n_20),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_22),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_23),
.C(n_20),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_13),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_20),
.B(n_13),
.C(n_11),
.D(n_19),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_118),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_10),
.Y(n_118)
);

AOI21x1_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_108),
.B(n_104),
.Y(n_120)
);

OAI21x1_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_116),
.B(n_112),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_111),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_19),
.C(n_21),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_130),
.A3(n_124),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_10),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_21),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

OAI21x1_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_9),
.B(n_19),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_131),
.A2(n_2),
.B(n_5),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_125),
.C(n_5),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_132),
.B1(n_133),
.B2(n_6),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_136),
.B1(n_7),
.B2(n_19),
.C(n_38),
.Y(n_137)
);


endmodule