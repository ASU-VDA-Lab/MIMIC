module fake_jpeg_7587_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_5),
.B(n_1),
.Y(n_7)
);

AOI21xp33_ASAP7_75t_SL g8 ( 
.A1(n_4),
.A2(n_1),
.B(n_0),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx2_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

HB1xp67_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_3),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_14),
.B(n_20),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_9),
.A2(n_10),
.B1(n_8),
.B2(n_6),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_16),
.B1(n_17),
.B2(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_9),
.A2(n_10),
.B1(n_8),
.B2(n_6),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_6),
.A2(n_3),
.B1(n_5),
.B2(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_1),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_26),
.B(n_27),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_32),
.B1(n_25),
.B2(n_14),
.Y(n_35)
);

AO22x1_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_29),
.B(n_32),
.Y(n_37)
);

OA21x2_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_18),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_32),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_20),
.B(n_18),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_40),
.B(n_36),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_40),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.C(n_37),
.Y(n_43)
);


endmodule