module fake_jpeg_19587_n_99 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_51),
.B1(n_37),
.B2(n_43),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_54),
.B(n_4),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_46),
.B1(n_45),
.B2(n_39),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_1),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_40),
.B1(n_36),
.B2(n_20),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_36),
.B1(n_1),
.B2(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_64),
.Y(n_66)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_75),
.B1(n_3),
.B2(n_34),
.Y(n_83)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_74),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_3),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_64),
.B(n_5),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_66),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_86),
.A3(n_87),
.B1(n_88),
.B2(n_77),
.C1(n_21),
.C2(n_22),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_70),
.B1(n_11),
.B2(n_13),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_8),
.B1(n_14),
.B2(n_15),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_79),
.A3(n_23),
.B1(n_25),
.B2(n_26),
.C1(n_28),
.C2(n_30),
.Y(n_90)
);

OA21x2_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_85),
.B(n_90),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_18),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_31),
.Y(n_95)
);

INVxp33_ASAP7_75t_SL g96 ( 
.A(n_95),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_96),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_33),
.B(n_81),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_81),
.Y(n_99)
);


endmodule