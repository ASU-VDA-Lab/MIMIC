module fake_aes_4262_n_51 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_51);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_51;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_48;
wire n_46;
wire n_25;
wire n_30;
wire n_26;
wire n_16;
wire n_33;
wire n_50;
wire n_49;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_8), .A2(n_15), .B1(n_6), .B2(n_10), .Y(n_16) );
BUFx3_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_2), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_5), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_5), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_0), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_1), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_3), .Y(n_23) );
AOI22xp5_ASAP7_75t_L g24 ( .A1(n_17), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_24) );
AND2x4_ASAP7_75t_L g25 ( .A(n_17), .B(n_3), .Y(n_25) );
NAND2xp5_ASAP7_75t_SL g26 ( .A(n_18), .B(n_4), .Y(n_26) );
BUFx3_ASAP7_75t_L g27 ( .A(n_18), .Y(n_27) );
AO22x1_ASAP7_75t_L g28 ( .A1(n_19), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_28) );
AOI221xp5_ASAP7_75t_SL g29 ( .A1(n_26), .A2(n_23), .B1(n_21), .B2(n_19), .C(n_20), .Y(n_29) );
AOI21xp5_ASAP7_75t_L g30 ( .A1(n_25), .A2(n_22), .B(n_20), .Y(n_30) );
AOI21xp5_ASAP7_75t_L g31 ( .A1(n_25), .A2(n_22), .B(n_23), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_33), .B(n_25), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
AND2x2_ASAP7_75t_L g38 ( .A(n_35), .B(n_34), .Y(n_38) );
AOI211x1_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_28), .B(n_35), .C(n_21), .Y(n_39) );
OAI221xp5_ASAP7_75t_L g40 ( .A1(n_38), .A2(n_24), .B1(n_29), .B2(n_16), .C(n_32), .Y(n_40) );
OAI22xp33_ASAP7_75t_L g41 ( .A1(n_36), .A2(n_16), .B1(n_35), .B2(n_28), .Y(n_41) );
NAND3xp33_ASAP7_75t_L g42 ( .A(n_39), .B(n_18), .C(n_36), .Y(n_42) );
OAI221xp5_ASAP7_75t_L g43 ( .A1(n_40), .A2(n_37), .B1(n_32), .B2(n_18), .C(n_27), .Y(n_43) );
NOR2xp33_ASAP7_75t_SL g44 ( .A(n_41), .B(n_37), .Y(n_44) );
NOR2x1_ASAP7_75t_L g45 ( .A(n_42), .B(n_18), .Y(n_45) );
NOR2x1_ASAP7_75t_L g46 ( .A(n_43), .B(n_27), .Y(n_46) );
OR3x2_ASAP7_75t_L g47 ( .A(n_44), .B(n_7), .C(n_8), .Y(n_47) );
OAI22xp5_ASAP7_75t_SL g48 ( .A1(n_47), .A2(n_9), .B1(n_11), .B2(n_12), .Y(n_48) );
AO22x2_ASAP7_75t_L g49 ( .A1(n_45), .A2(n_9), .B1(n_11), .B2(n_12), .Y(n_49) );
OAI22xp5_ASAP7_75t_L g50 ( .A1(n_48), .A2(n_46), .B1(n_13), .B2(n_14), .Y(n_50) );
OR2x6_ASAP7_75t_L g51 ( .A(n_50), .B(n_49), .Y(n_51) );
endmodule