module real_jpeg_548_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_1),
.A2(n_28),
.B1(n_32),
.B2(n_38),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_28),
.B1(n_49),
.B2(n_50),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_1),
.A2(n_28),
.B1(n_62),
.B2(n_66),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_62),
.B1(n_66),
.B2(n_71),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_2),
.A2(n_32),
.B1(n_38),
.B2(n_71),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_3),
.A2(n_32),
.B1(n_38),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_54),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_3),
.A2(n_54),
.B1(n_62),
.B2(n_66),
.Y(n_157)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_32),
.B1(n_38),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_57),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_5),
.A2(n_57),
.B1(n_62),
.B2(n_66),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_6),
.B(n_25),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_6),
.B(n_165),
.Y(n_202)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_6),
.A2(n_7),
.B(n_38),
.C(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_6),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_6),
.B(n_48),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_6),
.A2(n_32),
.B1(n_38),
.B2(n_215),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_6),
.B(n_62),
.C(n_65),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_215),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_6),
.B(n_87),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_6),
.B(n_60),
.Y(n_276)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_7),
.A2(n_38),
.B(n_47),
.C(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_7),
.B(n_38),
.Y(n_47)
);

AO22x2_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_8),
.A2(n_32),
.B1(n_38),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_8),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_8),
.A2(n_41),
.B1(n_62),
.B2(n_66),
.Y(n_190)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_12),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_12),
.A2(n_32),
.B1(n_38),
.B2(n_97),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_97),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_12),
.A2(n_62),
.B1(n_66),
.B2(n_97),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_13),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_13),
.A2(n_32),
.B1(n_38),
.B2(n_136),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_136),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_13),
.A2(n_62),
.B1(n_66),
.B2(n_136),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_15),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_15),
.A2(n_32),
.B1(n_38),
.B2(n_164),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_164),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_15),
.A2(n_62),
.B1(n_66),
.B2(n_164),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_111),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_109),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_20),
.B(n_98),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.C(n_79),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_21),
.B(n_73),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_42),
.B2(n_72),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_22),
.A2(n_23),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_23),
.B(n_43),
.C(n_59),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_31),
.B2(n_40),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_24),
.A2(n_31),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI32xp33_ASAP7_75t_L g185 ( 
.A1(n_26),
.A2(n_35),
.A3(n_38),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_26),
.A2(n_29),
.B(n_215),
.C(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_29),
.A2(n_31),
.B1(n_40),
.B2(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_29),
.A2(n_134),
.B(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_30),
.B(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_30),
.A2(n_135),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_31),
.B(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_31),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_31),
.A2(n_94),
.B(n_179),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_31)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_32),
.B(n_36),
.Y(n_187)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_53),
.B1(n_55),
.B2(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_45),
.A2(n_55),
.B1(n_56),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_45),
.A2(n_55),
.B1(n_75),
.B2(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_45),
.A2(n_181),
.B(n_183),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_45),
.A2(n_183),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_46),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_46),
.A2(n_48),
.B1(n_182),
.B2(n_199),
.Y(n_227)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_48),
.B(n_161),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_49),
.A2(n_52),
.B(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_50),
.B(n_260),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_55),
.A2(n_132),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_55),
.A2(n_160),
.B(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_59),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_67),
.B(n_69),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_60),
.A2(n_67),
.B1(n_92),
.B2(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_60),
.A2(n_67),
.B1(n_130),
.B2(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_60),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_70),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_77),
.B1(n_78),
.B2(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_61),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_61),
.A2(n_231),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_61),
.A2(n_77),
.B1(n_208),
.B2(n_242),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_62),
.B(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_67),
.A2(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_67),
.B(n_211),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_74),
.B(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_77),
.A2(n_210),
.B(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_93),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_80),
.A2(n_81),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_83),
.B1(n_93),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_82),
.A2(n_83),
.B1(n_90),
.B2(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_87),
.B(n_88),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_84),
.A2(n_87),
.B1(n_127),
.B2(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_84),
.A2(n_215),
.B(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_85),
.A2(n_86),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_85),
.A2(n_86),
.B1(n_190),
.B2(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_85),
.B(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_85),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_85),
.A2(n_86),
.B1(n_246),
.B2(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_86),
.A2(n_205),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_86),
.B(n_219),
.Y(n_248)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_87),
.A2(n_218),
.B(n_275),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_90),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_108),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_139),
.B(n_312),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_113),
.B(n_115),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_131),
.C(n_133),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_124),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_176),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_125),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_133),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_138),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_166),
.B(n_311),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_142),
.B(n_145),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_158),
.C(n_162),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_153),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_154),
.B(n_156),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_155),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_157),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_192),
.B(n_310),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_168),
.B(n_170),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.C(n_177),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_171),
.B(n_175),
.Y(n_295)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_177),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_184),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_178),
.B(n_180),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_184),
.B(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_188),
.B1(n_189),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI31xp33_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_292),
.A3(n_302),
.B(n_307),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_236),
.B(n_291),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_220),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_195),
.B(n_220),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.C(n_212),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_196),
.B(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_201),
.C(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_206),
.B(n_212),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_216),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_232),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_221),
.B(n_233),
.C(n_235),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_222),
.B(n_227),
.C(n_228),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_286),
.B(n_290),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_255),
.B(n_285),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_249),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_249),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_245),
.B1(n_264),
.B2(n_266),
.Y(n_263)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_253),
.C(n_254),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_267),
.B(n_284),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_263),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_263),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_278),
.B(n_283),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_273),
.B(n_277),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_276),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_281),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_289),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_296),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.C(n_300),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_306),
.Y(n_308)
);


endmodule