module fake_jpeg_3487_n_711 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_711);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_711;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_544;
wire n_455;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_62),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_111),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_64),
.Y(n_201)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_65),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_68),
.Y(n_224)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g207 ( 
.A(n_71),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_72),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_74),
.Y(n_184)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_75),
.Y(n_200)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_77),
.B(n_112),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_80),
.Y(n_183)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_82),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_83),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_90),
.Y(n_220)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_92),
.Y(n_229)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_93),
.Y(n_196)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_96),
.Y(n_215)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_29),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_99),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_105),
.Y(n_214)
);

BUFx16f_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_108),
.Y(n_225)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_26),
.B(n_19),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_26),
.B(n_18),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_119),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_115),
.Y(n_231)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_116),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_117),
.Y(n_181)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_44),
.B(n_18),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_53),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_33),
.Y(n_123)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

BUFx8_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_126),
.B(n_130),
.Y(n_191)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_47),
.Y(n_129)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

BUFx12f_ASAP7_75t_SL g130 ( 
.A(n_47),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_132),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_47),
.Y(n_133)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_139),
.B(n_186),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_77),
.B(n_50),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_141),
.B(n_157),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_71),
.A2(n_21),
.B1(n_22),
.B2(n_31),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_149),
.B(n_166),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_44),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_21),
.B1(n_22),
.B2(n_38),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g263 ( 
.A1(n_165),
.A2(n_172),
.B1(n_198),
.B2(n_37),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_80),
.B(n_50),
.Y(n_166)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_116),
.A2(n_22),
.B1(n_38),
.B2(n_31),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_82),
.B(n_59),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_173),
.B(n_132),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_92),
.A2(n_59),
.B1(n_40),
.B2(n_30),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_180),
.A2(n_197),
.B1(n_219),
.B2(n_221),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_66),
.B(n_38),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_72),
.B(n_21),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_187),
.B(n_192),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_84),
.B(n_31),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_133),
.B(n_20),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_195),
.B(n_210),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_96),
.A2(n_59),
.B1(n_20),
.B2(n_30),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_85),
.A2(n_20),
.B1(n_40),
.B2(n_30),
.Y(n_198)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_128),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_85),
.B(n_57),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_216),
.Y(n_234)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_61),
.Y(n_217)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_62),
.Y(n_218)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_60),
.A2(n_40),
.B1(n_55),
.B2(n_52),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_64),
.A2(n_41),
.B1(n_55),
.B2(n_52),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_88),
.Y(n_222)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_90),
.B(n_41),
.Y(n_223)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_223),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_78),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_197),
.B1(n_113),
.B2(n_115),
.Y(n_253)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_100),
.Y(n_228)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_97),
.B(n_41),
.Y(n_230)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_233),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_191),
.A2(n_32),
.B1(n_24),
.B2(n_28),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_237),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_239),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_191),
.A2(n_195),
.B1(n_207),
.B2(n_28),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_SL g377 ( 
.A(n_241),
.B(n_153),
.C(n_151),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_152),
.B(n_32),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_242),
.B(n_254),
.Y(n_354)
);

O2A1O1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_93),
.B(n_32),
.C(n_57),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_243),
.A2(n_273),
.B(n_136),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_180),
.A2(n_104),
.B1(n_120),
.B2(n_117),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_246),
.A2(n_253),
.B1(n_309),
.B2(n_224),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_207),
.A2(n_49),
.B1(n_24),
.B2(n_35),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_247),
.A2(n_251),
.B1(n_283),
.B2(n_292),
.Y(n_337)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_140),
.Y(n_248)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_248),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_162),
.A2(n_52),
.B1(n_35),
.B2(n_37),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_154),
.A2(n_49),
.B1(n_35),
.B2(n_37),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_252),
.B(n_3),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_135),
.B(n_28),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_177),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_258),
.B(n_267),
.Y(n_338)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_134),
.Y(n_260)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_260),
.Y(n_321)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_213),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_261),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_159),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_262),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_263),
.B(n_282),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_150),
.B(n_45),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_265),
.B(n_274),
.Y(n_369)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_137),
.Y(n_266)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_177),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_143),
.Y(n_268)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_268),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_138),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_269),
.Y(n_319)
);

INVx4_ASAP7_75t_SL g270 ( 
.A(n_232),
.Y(n_270)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_270),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_169),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_271),
.B(n_288),
.Y(n_370)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_145),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_272),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_172),
.A2(n_57),
.B(n_55),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_158),
.B(n_45),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_147),
.B(n_107),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_275),
.B(n_277),
.Y(n_330)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_140),
.Y(n_276)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_276),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_148),
.B(n_0),
.Y(n_277)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_164),
.Y(n_279)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_279),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_165),
.A2(n_129),
.B1(n_49),
.B2(n_45),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_280),
.A2(n_295),
.B1(n_297),
.B2(n_299),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_194),
.A2(n_47),
.B1(n_15),
.B2(n_14),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_281),
.A2(n_310),
.B1(n_315),
.B2(n_208),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_200),
.B(n_0),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_200),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_176),
.Y(n_284)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_284),
.Y(n_376)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_220),
.Y(n_285)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_285),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_190),
.B(n_0),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_296),
.C(n_178),
.Y(n_336)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_174),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_287),
.B(n_304),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_205),
.B(n_1),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_289),
.Y(n_349)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_160),
.Y(n_290)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_203),
.Y(n_291)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

INVx11_ASAP7_75t_L g292 ( 
.A(n_142),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_193),
.Y(n_293)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_293),
.Y(n_360)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_189),
.Y(n_294)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_185),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_161),
.B(n_15),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_215),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_185),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_168),
.Y(n_300)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_145),
.Y(n_301)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_301),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_188),
.B(n_1),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_302),
.B(n_312),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_201),
.Y(n_303)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_303),
.Y(n_371)
);

BUFx12f_ASAP7_75t_L g304 ( 
.A(n_171),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_194),
.Y(n_305)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_144),
.Y(n_308)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_183),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_156),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_144),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_311),
.B(n_316),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_181),
.B(n_2),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_182),
.A2(n_206),
.B1(n_146),
.B2(n_199),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_313),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_201),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_314),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_175),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_169),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_184),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_317),
.B(n_9),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_250),
.A2(n_231),
.B1(n_227),
.B2(n_184),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_320),
.Y(n_397)
);

OR2x4_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_214),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_322),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_265),
.A2(n_231),
.B1(n_227),
.B2(n_224),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_324),
.A2(n_374),
.B1(n_233),
.B2(n_303),
.Y(n_416)
);

NAND2xp67_ASAP7_75t_L g325 ( 
.A(n_263),
.B(n_243),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_325),
.A2(n_344),
.B(n_372),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_326),
.A2(n_347),
.B1(n_313),
.B2(n_289),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_329),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_254),
.B(n_212),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_331),
.B(n_334),
.C(n_348),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_245),
.B(n_202),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_336),
.B(n_270),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_264),
.B(n_179),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_339),
.B(n_341),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_259),
.B(n_225),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_278),
.A2(n_208),
.B(n_178),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_241),
.A2(n_146),
.B1(n_199),
.B2(n_229),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_211),
.C(n_142),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_274),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_350),
.B(n_353),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_239),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_307),
.B(n_211),
.C(n_142),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_275),
.C(n_282),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_362),
.A2(n_5),
.B(n_6),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_366),
.Y(n_392)
);

AOI32xp33_ASAP7_75t_L g367 ( 
.A1(n_298),
.A2(n_229),
.A3(n_209),
.B1(n_183),
.B2(n_155),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_367),
.B(n_380),
.Y(n_424)
);

AO22x1_ASAP7_75t_L g372 ( 
.A1(n_246),
.A2(n_151),
.B1(n_209),
.B2(n_136),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_234),
.A2(n_155),
.B1(n_153),
.B2(n_151),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_273),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_5),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_385),
.A2(n_396),
.B1(n_399),
.B2(n_407),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_386),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_322),
.A2(n_263),
.B1(n_236),
.B2(n_242),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_388),
.A2(n_406),
.B(n_411),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_318),
.B(n_288),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_404),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_390),
.B(n_395),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_391),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_331),
.B(n_296),
.C(n_260),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_413),
.C(n_422),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_350),
.A2(n_263),
.B1(n_312),
.B2(n_302),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_326),
.A2(n_286),
.B1(n_277),
.B2(n_275),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_398),
.A2(n_400),
.B1(n_405),
.B2(n_414),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_369),
.A2(n_252),
.B1(n_286),
.B2(n_277),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_357),
.A2(n_282),
.B1(n_244),
.B2(n_255),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_321),
.Y(n_401)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_401),
.Y(n_442)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_402),
.Y(n_449)
);

INVx11_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_403),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_293),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_357),
.A2(n_305),
.B1(n_284),
.B2(n_279),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_357),
.A2(n_256),
.B(n_235),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_357),
.A2(n_272),
.B1(n_249),
.B2(n_238),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_318),
.B(n_249),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_408),
.B(n_410),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_238),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_335),
.A2(n_292),
.B1(n_311),
.B2(n_308),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_334),
.B(n_354),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_412),
.B(n_417),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_354),
.B(n_268),
.C(n_266),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_357),
.A2(n_257),
.B1(n_294),
.B2(n_276),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_349),
.Y(n_415)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_415),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_416),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_336),
.B(n_257),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_347),
.A2(n_314),
.B1(n_301),
.B2(n_248),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_418),
.A2(n_425),
.B1(n_397),
.B2(n_372),
.Y(n_437)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_419),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_332),
.A2(n_300),
.B(n_285),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_420),
.A2(n_427),
.B(n_337),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_330),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_348),
.B(n_261),
.C(n_291),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_341),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_428),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_362),
.A2(n_262),
.B1(n_290),
.B2(n_304),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_351),
.Y(n_426)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_426),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_335),
.A2(n_304),
.B1(n_287),
.B2(n_8),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_373),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_429),
.B(n_430),
.Y(n_440)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_360),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_356),
.B(n_287),
.C(n_6),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_330),
.C(n_332),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_432),
.A2(n_366),
.B(n_344),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_409),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_435),
.B(n_447),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_437),
.A2(n_453),
.B1(n_383),
.B2(n_458),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_443),
.A2(n_426),
.B1(n_411),
.B2(n_375),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_409),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_448),
.B(n_384),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_452),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_404),
.B(n_330),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_394),
.A2(n_325),
.B1(n_363),
.B2(n_329),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_454),
.B(n_467),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_421),
.B(n_360),
.C(n_338),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_466),
.C(n_468),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_396),
.A2(n_372),
.B1(n_381),
.B2(n_327),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_458),
.A2(n_434),
.B1(n_453),
.B2(n_435),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_389),
.B(n_378),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_460),
.B(n_462),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_432),
.A2(n_353),
.B(n_319),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_394),
.A2(n_319),
.B(n_342),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_463),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_426),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_469),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_408),
.B(n_339),
.Y(n_465)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_465),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_384),
.B(n_361),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_410),
.B(n_361),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_417),
.B(n_359),
.C(n_364),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_388),
.A2(n_359),
.B(n_364),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_387),
.A2(n_323),
.B(n_328),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_471),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_399),
.B(n_340),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_472),
.B(n_431),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_387),
.A2(n_327),
.B1(n_351),
.B2(n_371),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_474),
.A2(n_407),
.B1(n_390),
.B2(n_400),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_406),
.A2(n_358),
.B(n_375),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_475),
.B(n_469),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_476),
.A2(n_504),
.B1(n_512),
.B2(n_472),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_479),
.A2(n_477),
.B1(n_490),
.B2(n_481),
.Y(n_535)
);

FAx1_ASAP7_75t_L g481 ( 
.A(n_436),
.B(n_424),
.CI(n_405),
.CON(n_481),
.SN(n_481)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_481),
.A2(n_503),
.B(n_513),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_485),
.B(n_493),
.C(n_499),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_412),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_459),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_473),
.A2(n_434),
.B1(n_458),
.B2(n_453),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_488),
.A2(n_494),
.B1(n_495),
.B2(n_502),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_489),
.A2(n_436),
.B1(n_474),
.B2(n_457),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_440),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_497),
.Y(n_517)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_491),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_439),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_492),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_446),
.B(n_413),
.C(n_393),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_434),
.A2(n_424),
.B1(n_385),
.B2(n_397),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_447),
.A2(n_382),
.B1(n_398),
.B2(n_425),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_445),
.Y(n_496)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_496),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_445),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_470),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_498),
.B(n_464),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_466),
.B(n_386),
.C(n_422),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_467),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_500),
.B(n_511),
.Y(n_539)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_442),
.Y(n_501)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_501),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_460),
.A2(n_382),
.B1(n_392),
.B2(n_414),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_441),
.A2(n_395),
.B1(n_418),
.B2(n_420),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_436),
.A2(n_395),
.B1(n_401),
.B2(n_402),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_506),
.A2(n_451),
.B1(n_437),
.B2(n_470),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_508),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_444),
.B(n_454),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_509),
.B(n_510),
.C(n_514),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_444),
.B(n_419),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_442),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_441),
.A2(n_395),
.B1(n_416),
.B2(n_415),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_444),
.B(n_429),
.C(n_428),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_454),
.B(n_430),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_515),
.B(n_448),
.C(n_463),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_456),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_516),
.B(n_518),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_456),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_520),
.B(n_545),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_459),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_521),
.B(n_540),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_526),
.A2(n_537),
.B1(n_505),
.B2(n_480),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_496),
.B(n_465),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_527),
.B(n_549),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_529),
.A2(n_531),
.B1(n_533),
.B2(n_555),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_484),
.B(n_438),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_530),
.B(n_501),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_489),
.A2(n_474),
.B1(n_462),
.B2(n_436),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_494),
.A2(n_462),
.B1(n_471),
.B2(n_457),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_482),
.A2(n_471),
.B(n_450),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_534),
.Y(n_587)
);

OAI22x1_ASAP7_75t_L g565 ( 
.A1(n_535),
.A2(n_533),
.B1(n_555),
.B2(n_504),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_482),
.A2(n_478),
.B(n_433),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_536),
.A2(n_443),
.B(n_476),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_481),
.A2(n_450),
.B1(n_438),
.B2(n_437),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_538),
.B(n_498),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_486),
.B(n_468),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_505),
.B(n_468),
.Y(n_541)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_541),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_483),
.B(n_448),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_SL g558 ( 
.A(n_542),
.B(n_516),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_500),
.B(n_452),
.Y(n_543)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_543),
.Y(n_582)
);

CKINVDCx14_ASAP7_75t_R g544 ( 
.A(n_505),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_544),
.A2(n_507),
.B1(n_480),
.B2(n_498),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_486),
.B(n_499),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_546),
.B(n_553),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_514),
.B(n_463),
.C(n_475),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_548),
.B(n_550),
.C(n_493),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_484),
.B(n_455),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_487),
.B(n_433),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_491),
.B(n_449),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_552),
.B(n_355),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_515),
.B(n_449),
.Y(n_553)
);

AND2x4_ASAP7_75t_SL g554 ( 
.A(n_507),
.B(n_455),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_554),
.B(n_508),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_556),
.A2(n_568),
.B(n_524),
.Y(n_605)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_557),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_SL g598 ( 
.A(n_558),
.B(n_560),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_559),
.A2(n_579),
.B1(n_581),
.B2(n_588),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_554),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_561),
.B(n_562),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_554),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_506),
.Y(n_563)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_563),
.Y(n_606)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_565),
.Y(n_608)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_522),
.Y(n_566)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_566),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_521),
.B(n_358),
.Y(n_569)
);

NOR2xp67_ASAP7_75t_L g616 ( 
.A(n_569),
.B(n_574),
.Y(n_616)
);

CKINVDCx14_ASAP7_75t_R g609 ( 
.A(n_570),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_539),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_572),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_517),
.B(n_511),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_573),
.B(n_580),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_532),
.B(n_439),
.Y(n_574)
);

XNOR2x1_ASAP7_75t_L g578 ( 
.A(n_550),
.B(n_483),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_578),
.B(n_518),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_528),
.A2(n_512),
.B1(n_513),
.B2(n_451),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_526),
.A2(n_492),
.B1(n_461),
.B2(n_368),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_583),
.B(n_355),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_525),
.B(n_379),
.C(n_343),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_584),
.B(n_585),
.C(n_586),
.Y(n_592)
);

BUFx24_ASAP7_75t_SL g585 ( 
.A(n_546),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_525),
.B(n_379),
.C(n_343),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_538),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_588),
.A2(n_590),
.B1(n_551),
.B2(n_522),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_529),
.A2(n_368),
.B1(n_371),
.B2(n_351),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_591),
.B(n_601),
.Y(n_631)
);

INVx13_ASAP7_75t_L g593 ( 
.A(n_566),
.Y(n_593)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_593),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g594 ( 
.A1(n_579),
.A2(n_531),
.B1(n_519),
.B2(n_537),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_594),
.A2(n_603),
.B1(n_610),
.B2(n_580),
.Y(n_634)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_596),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_523),
.C(n_540),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_599),
.B(n_613),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_600),
.A2(n_391),
.B1(n_345),
.B2(n_340),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_577),
.B(n_575),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_SL g602 ( 
.A(n_578),
.B(n_547),
.Y(n_602)
);

OAI21xp33_ASAP7_75t_L g639 ( 
.A1(n_602),
.A2(n_391),
.B(n_333),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_559),
.A2(n_536),
.B1(n_534),
.B2(n_524),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_605),
.A2(n_617),
.B(n_365),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_582),
.A2(n_548),
.B1(n_553),
.B2(n_545),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_577),
.B(n_523),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g640 ( 
.A(n_611),
.B(n_352),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_612),
.B(n_590),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_589),
.B(n_564),
.C(n_575),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_564),
.B(n_520),
.C(n_542),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_614),
.B(n_618),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_587),
.A2(n_403),
.B(n_323),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_584),
.B(n_355),
.C(n_345),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_SL g619 ( 
.A1(n_608),
.A2(n_587),
.B(n_571),
.C(n_557),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_619),
.A2(n_637),
.B(n_639),
.Y(n_654)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_620),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_601),
.B(n_611),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_621),
.B(n_624),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_616),
.Y(n_622)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_622),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_608),
.A2(n_568),
.B1(n_563),
.B2(n_576),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_SL g643 ( 
.A1(n_623),
.A2(n_600),
.B1(n_597),
.B2(n_604),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_610),
.B(n_565),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_599),
.B(n_560),
.C(n_586),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_625),
.B(n_626),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_609),
.B(n_567),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_605),
.A2(n_571),
.B(n_573),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_627),
.A2(n_595),
.B(n_596),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_613),
.B(n_558),
.C(n_580),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_632),
.B(n_633),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_607),
.A2(n_581),
.B1(n_580),
.B2(n_403),
.Y(n_633)
);

XOR2xp5_ASAP7_75t_L g649 ( 
.A(n_634),
.B(n_638),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_592),
.B(n_614),
.C(n_598),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_635),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_592),
.B(n_598),
.C(n_618),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_636),
.B(n_640),
.C(n_642),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_603),
.B(n_591),
.C(n_615),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_643),
.B(n_648),
.Y(n_668)
);

OAI21xp33_ASAP7_75t_L g672 ( 
.A1(n_647),
.A2(n_650),
.B(n_619),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_625),
.B(n_615),
.C(n_594),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_SL g650 ( 
.A1(n_627),
.A2(n_604),
.B(n_597),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_628),
.B(n_606),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_651),
.B(n_652),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_642),
.B(n_602),
.C(n_606),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_621),
.B(n_617),
.C(n_612),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_655),
.B(n_658),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_629),
.B(n_593),
.C(n_333),
.Y(n_658)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_630),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_660),
.A2(n_662),
.B1(n_376),
.B2(n_352),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_623),
.B(n_346),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g665 ( 
.A(n_661),
.B(n_624),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_641),
.B(n_346),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_657),
.B(n_620),
.Y(n_663)
);

AOI21xp33_ASAP7_75t_L g685 ( 
.A1(n_663),
.A2(n_674),
.B(n_654),
.Y(n_685)
);

XNOR2xp5_ASAP7_75t_L g664 ( 
.A(n_646),
.B(n_636),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_664),
.B(n_669),
.Y(n_690)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_665),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_659),
.B(n_634),
.Y(n_666)
);

NAND2x1_ASAP7_75t_L g689 ( 
.A(n_666),
.B(n_667),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_SL g667 ( 
.A1(n_656),
.A2(n_632),
.B(n_637),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_653),
.B(n_635),
.C(n_631),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g670 ( 
.A(n_646),
.B(n_648),
.C(n_652),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_670),
.B(n_671),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g671 ( 
.A(n_658),
.B(n_640),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g684 ( 
.A(n_672),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_644),
.B(n_631),
.C(n_619),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_673),
.B(n_655),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_645),
.B(n_619),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_676),
.B(n_678),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_644),
.B(n_376),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_680),
.B(n_681),
.Y(n_692)
);

MAJIxp5_ASAP7_75t_L g681 ( 
.A(n_666),
.B(n_649),
.C(n_647),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_677),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_682),
.B(n_668),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_663),
.B(n_650),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_683),
.A2(n_688),
.B(n_352),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_685),
.A2(n_672),
.B(n_674),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_675),
.B(n_662),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_SL g700 ( 
.A1(n_691),
.A2(n_694),
.B(n_684),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_693),
.B(n_695),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_SL g694 ( 
.A1(n_690),
.A2(n_643),
.B(n_654),
.Y(n_694)
);

MAJIxp5_ASAP7_75t_L g695 ( 
.A(n_687),
.B(n_678),
.C(n_649),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_696),
.A2(n_698),
.B(n_689),
.Y(n_702)
);

XOR2xp5_ASAP7_75t_L g697 ( 
.A(n_681),
.B(n_5),
.Y(n_697)
);

XOR2xp5_ASAP7_75t_L g699 ( 
.A(n_697),
.B(n_689),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_SL g698 ( 
.A1(n_684),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_698)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_699),
.A2(n_700),
.B(n_701),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g701 ( 
.A(n_692),
.B(n_679),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_SL g704 ( 
.A1(n_702),
.A2(n_692),
.B(n_686),
.Y(n_704)
);

XNOR2xp5_ASAP7_75t_L g707 ( 
.A(n_704),
.B(n_706),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_SL g706 ( 
.A1(n_703),
.A2(n_682),
.B(n_686),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_705),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_708),
.B(n_698),
.Y(n_709)
);

XOR2xp5_ASAP7_75t_L g710 ( 
.A(n_709),
.B(n_707),
.Y(n_710)
);

XOR2xp5_ASAP7_75t_L g711 ( 
.A(n_710),
.B(n_8),
.Y(n_711)
);


endmodule