module fake_jpeg_16344_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g84 ( 
.A(n_46),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_20),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_17),
.B1(n_29),
.B2(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_57),
.B1(n_19),
.B2(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_62),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_SL g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_19),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_32),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_63),
.B1(n_16),
.B2(n_18),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_29),
.B1(n_24),
.B2(n_30),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_77),
.B1(n_94),
.B2(n_61),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_74),
.B(n_88),
.Y(n_117)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_29),
.B1(n_45),
.B2(n_27),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_83),
.Y(n_122)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_28),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_33),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_95),
.Y(n_123)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_16),
.B1(n_18),
.B2(n_27),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_33),
.B1(n_23),
.B2(n_34),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_24),
.B1(n_30),
.B2(n_16),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_33),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_99),
.Y(n_110)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_18),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_46),
.B(n_27),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_61),
.B(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_54),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_113),
.B1(n_125),
.B2(n_78),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_108),
.B1(n_71),
.B2(n_91),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_87),
.B1(n_78),
.B2(n_89),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_64),
.B1(n_66),
.B2(n_46),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_119),
.Y(n_131)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_68),
.B(n_31),
.CI(n_33),
.CON(n_120),
.SN(n_120)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_127),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_76),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_31),
.B(n_1),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_126),
.B(n_73),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_68),
.A2(n_66),
.B1(n_14),
.B2(n_15),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_34),
.B1(n_30),
.B2(n_21),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_135),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_67),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_134),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_88),
.A3(n_74),
.B1(n_67),
.B2(n_87),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_136),
.B(n_147),
.Y(n_165)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_98),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_146),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_87),
.B1(n_101),
.B2(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_145),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_117),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_100),
.B1(n_75),
.B2(n_84),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_150),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_99),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_154),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_157),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_115),
.B1(n_112),
.B2(n_123),
.Y(n_172)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_155),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_77),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_127),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_159),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_77),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_59),
.C(n_92),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_125),
.C(n_102),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_77),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_117),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_110),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_164),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_124),
.B1(n_113),
.B2(n_118),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_171),
.B1(n_172),
.B2(n_188),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_123),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_183),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_115),
.B1(n_126),
.B2(n_121),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_186),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_119),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_138),
.B1(n_154),
.B2(n_78),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_129),
.B(n_102),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_143),
.B(n_158),
.Y(n_204)
);

AOI221xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_150),
.B1(n_139),
.B2(n_34),
.C(n_32),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_180),
.B(n_132),
.CI(n_12),
.CON(n_215),
.SN(n_215)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_114),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_31),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_66),
.Y(n_185)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_21),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_82),
.B1(n_83),
.B2(n_97),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_148),
.B1(n_153),
.B2(n_160),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_82),
.B1(n_92),
.B2(n_70),
.Y(n_218)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_59),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_59),
.C(n_70),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_132),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_134),
.B(n_86),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_199),
.B(n_200),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_174),
.B(n_131),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_218),
.B1(n_196),
.B2(n_184),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_211),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_183),
.C(n_186),
.Y(n_233)
);

OA21x2_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_177),
.B(n_215),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_132),
.B(n_1),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_172),
.B(n_191),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_215),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_169),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_21),
.Y(n_217)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_163),
.B(n_33),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_220),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_223),
.A2(n_224),
.B1(n_211),
.B2(n_219),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_225),
.C(n_192),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_169),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_227),
.A2(n_235),
.B1(n_247),
.B2(n_248),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_170),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_209),
.A2(n_196),
.B1(n_168),
.B2(n_167),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_232),
.A2(n_197),
.B1(n_217),
.B2(n_206),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_234),
.C(n_243),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_165),
.C(n_176),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_241),
.Y(n_264)
);

AO22x1_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_175),
.B1(n_168),
.B2(n_164),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_165),
.C(n_189),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_201),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_173),
.C(n_180),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_207),
.C(n_212),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_179),
.B1(n_188),
.B2(n_185),
.Y(n_247)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_213),
.B1(n_202),
.B2(n_197),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_261),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_237),
.B1(n_202),
.B2(n_249),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_260),
.C(n_267),
.Y(n_271)
);

AOI22x1_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_215),
.B1(n_210),
.B2(n_212),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_258),
.B(n_262),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_247),
.A2(n_237),
.B1(n_227),
.B2(n_249),
.Y(n_259)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_219),
.C(n_214),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_179),
.B1(n_214),
.B2(n_220),
.Y(n_261)
);

NAND2x1_ASAP7_75t_SL g262 ( 
.A(n_226),
.B(n_171),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_266),
.Y(n_276)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_166),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_243),
.C(n_232),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_223),
.B1(n_184),
.B2(n_192),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_240),
.B1(n_190),
.B2(n_193),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_282),
.C(n_254),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_229),
.C(n_230),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_284),
.C(n_285),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_258),
.B(n_242),
.CI(n_228),
.CON(n_278),
.SN(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_226),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_259),
.B(n_240),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_242),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_25),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_248),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_269),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_190),
.C(n_23),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_267),
.C(n_252),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_286),
.A2(n_262),
.B1(n_2),
.B2(n_3),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

OAI221xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_253),
.B1(n_256),
.B2(n_261),
.C(n_263),
.Y(n_288)
);

NOR2x1p5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_300),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_292),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_296),
.C(n_271),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_274),
.B1(n_284),
.B2(n_273),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_23),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_32),
.C(n_25),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_299),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_25),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_301),
.A2(n_312),
.A3(n_10),
.B1(n_9),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_307),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_290),
.A2(n_281),
.B1(n_282),
.B2(n_278),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_308),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_285),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_15),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_311),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_58),
.B(n_12),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_297),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_316),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_300),
.B1(n_11),
.B2(n_10),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_318),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_58),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_23),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_1),
.C2(n_6),
.Y(n_319)
);

AOI31xp67_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_321),
.A3(n_5),
.B(n_7),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_304),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_309),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_316),
.A2(n_304),
.B1(n_6),
.B2(n_7),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_323),
.B(n_326),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_5),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_317),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_325),
.A2(n_320),
.B(n_314),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_320),
.C(n_328),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_329),
.C(n_8),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_8),
.Y(n_333)
);


endmodule