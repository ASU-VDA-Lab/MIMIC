module fake_jpeg_216_n_694 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_694);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_694;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_553;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_SL g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_61),
.B(n_68),
.Y(n_210)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_64),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_65),
.Y(n_223)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_67),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_19),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_71),
.B(n_84),
.Y(n_148)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_73),
.Y(n_220)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_76),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_78),
.Y(n_183)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_79),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_81),
.Y(n_194)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_82),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_86),
.Y(n_207)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_88),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_30),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_89),
.B(n_92),
.Y(n_164)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_30),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_93),
.Y(n_233)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_31),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_100),
.B(n_101),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_31),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_102),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_37),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_105),
.B(n_106),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_22),
.B(n_19),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_32),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_120),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_27),
.B(n_1),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_112),
.B(n_43),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_37),
.B(n_19),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_29),
.Y(n_143)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_115),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_35),
.Y(n_116)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_40),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_124),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_127),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx6_ASAP7_75t_SL g129 ( 
.A(n_39),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g180 ( 
.A(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_27),
.Y(n_130)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_132),
.Y(n_201)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_28),
.Y(n_133)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_143),
.B(n_177),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_76),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_150),
.B(n_175),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_56),
.B1(n_54),
.B2(n_43),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_153),
.A2(n_169),
.B1(n_9),
.B2(n_10),
.Y(n_292)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_62),
.B(n_54),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_154),
.B(n_228),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_69),
.A2(n_48),
.B1(n_56),
.B2(n_58),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g313 ( 
.A1(n_160),
.A2(n_218),
.B1(n_14),
.B2(n_15),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_161),
.B(n_219),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_77),
.A2(n_56),
.B1(n_29),
.B2(n_50),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_70),
.B(n_44),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_80),
.B(n_44),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_73),
.Y(n_179)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_179),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_83),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_186),
.B(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_187),
.Y(n_271)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_60),
.Y(n_191)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_74),
.Y(n_196)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_196),
.Y(n_286)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_63),
.B(n_1),
.Y(n_198)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_198),
.A2(n_42),
.A3(n_55),
.B1(n_49),
.B2(n_24),
.Y(n_254)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_81),
.Y(n_199)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_199),
.Y(n_288)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_93),
.Y(n_202)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_202),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_80),
.B(n_28),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_211),
.Y(n_246)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_95),
.Y(n_208)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_88),
.B(n_33),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_127),
.B(n_33),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_213),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_88),
.B(n_50),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_104),
.B(n_34),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_224),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_65),
.A2(n_48),
.B1(n_56),
.B2(n_55),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_86),
.B(n_53),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_96),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_104),
.B(n_53),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_116),
.B(n_34),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_226),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_65),
.B(n_58),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_108),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_230),
.B(n_234),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_116),
.B(n_58),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_110),
.Y(n_234)
);

HAxp5_ASAP7_75t_SL g235 ( 
.A(n_180),
.B(n_48),
.CON(n_235),
.SN(n_235)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_235),
.B(n_238),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_118),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_239),
.Y(n_336)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_135),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_241),
.Y(n_359)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_149),
.Y(n_242)
);

BUFx4f_ASAP7_75t_SL g373 ( 
.A(n_242),
.Y(n_373)
);

OR2x2_ASAP7_75t_SL g243 ( 
.A(n_156),
.B(n_36),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g333 ( 
.A(n_243),
.B(n_254),
.C(n_296),
.Y(n_333)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_183),
.Y(n_244)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_244),
.Y(n_343)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_245),
.Y(n_348)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_135),
.Y(n_247)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_247),
.Y(n_370)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_248),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_145),
.A2(n_94),
.B1(n_90),
.B2(n_36),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_250),
.A2(n_251),
.B1(n_283),
.B2(n_297),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_145),
.A2(n_24),
.B1(n_55),
.B2(n_49),
.Y(n_251)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_184),
.Y(n_255)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_255),
.Y(n_367)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_197),
.Y(n_257)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_257),
.Y(n_382)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_134),
.Y(n_258)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_258),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_175),
.A2(n_24),
.B1(n_49),
.B2(n_36),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_158),
.A2(n_131),
.B1(n_128),
.B2(n_126),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_210),
.A2(n_124),
.B1(n_123),
.B2(n_122),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_261),
.A2(n_317),
.B1(n_318),
.B2(n_174),
.Y(n_380)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_262),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_198),
.A2(n_1),
.B(n_2),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_263),
.A2(n_283),
.B(n_276),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_154),
.A2(n_121),
.B1(n_119),
.B2(n_117),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_264),
.A2(n_276),
.B1(n_292),
.B2(n_300),
.Y(n_369)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_136),
.Y(n_265)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_265),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_165),
.B(n_118),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_267),
.B(n_273),
.Y(n_330)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_188),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_268),
.Y(n_332)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_167),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_270),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_148),
.B(n_111),
.Y(n_273)
);

AO22x2_ASAP7_75t_L g274 ( 
.A1(n_142),
.A2(n_45),
.B1(n_42),
.B2(n_4),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_274),
.B(n_289),
.Y(n_357)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_134),
.Y(n_275)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_275),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_L g276 ( 
.A1(n_160),
.A2(n_45),
.B1(n_42),
.B2(n_4),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_152),
.Y(n_277)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_277),
.Y(n_365)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_136),
.Y(n_278)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_278),
.Y(n_362)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_152),
.Y(n_279)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_279),
.Y(n_371)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_178),
.Y(n_280)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_280),
.Y(n_378)
);

A2O1A1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_166),
.A2(n_42),
.B(n_2),
.C(n_5),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_282),
.B(n_287),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_159),
.A2(n_42),
.B1(n_2),
.B2(n_5),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_164),
.B(n_1),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_284),
.B(n_290),
.Y(n_344)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_178),
.Y(n_285)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_285),
.Y(n_385)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_228),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_287)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_138),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_176),
.B(n_7),
.Y(n_290)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_163),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_291),
.Y(n_324)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_190),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_294),
.Y(n_331)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_163),
.Y(n_294)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_181),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_295),
.B(n_302),
.Y(n_335)
);

CKINVDCx9p33_ASAP7_75t_R g296 ( 
.A(n_173),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_151),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_137),
.B(n_10),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_298),
.B(n_304),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_218),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_300)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_206),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_201),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_306),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_141),
.B(n_11),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_157),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_305),
.B(n_308),
.Y(n_384)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_214),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_141),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_151),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_309),
.A2(n_162),
.B1(n_159),
.B2(n_209),
.Y(n_345)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_144),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_312),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_215),
.B(n_13),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_313),
.A2(n_319),
.B1(n_320),
.B2(n_140),
.Y(n_355)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_181),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_315),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_221),
.B(n_15),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_221),
.B(n_16),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_316),
.B(n_321),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_168),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_139),
.A2(n_16),
.B1(n_18),
.B2(n_232),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_168),
.Y(n_319)
);

INVx13_ASAP7_75t_L g320 ( 
.A(n_223),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_146),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_220),
.B(n_18),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_322),
.B(n_18),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_238),
.B(n_229),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_326),
.B(n_327),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_249),
.B(n_182),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_266),
.B(n_182),
.C(n_207),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_328),
.B(n_334),
.C(n_305),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_237),
.B(n_195),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_263),
.B(n_195),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_337),
.B(n_349),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_189),
.B1(n_204),
.B2(n_200),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_338),
.A2(n_345),
.B1(n_278),
.B2(n_265),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_282),
.B(n_207),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_287),
.A2(n_162),
.B(n_157),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_351),
.A2(n_358),
.B(n_291),
.Y(n_418)
);

OAI22xp33_ASAP7_75t_L g352 ( 
.A1(n_313),
.A2(n_232),
.B1(n_139),
.B2(n_209),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_352),
.A2(n_360),
.B1(n_375),
.B2(n_380),
.Y(n_406)
);

AOI32xp33_ASAP7_75t_L g354 ( 
.A1(n_246),
.A2(n_206),
.A3(n_147),
.B1(n_205),
.B2(n_170),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_354),
.B(n_235),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_355),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_272),
.B(n_140),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_356),
.B(n_366),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_272),
.A2(n_253),
.B1(n_252),
.B2(n_307),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_317),
.A2(n_189),
.B1(n_204),
.B2(n_200),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_313),
.A2(n_227),
.B1(n_170),
.B2(n_140),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_174),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_374),
.B(n_155),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_273),
.A2(n_227),
.B1(n_193),
.B2(n_172),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_269),
.B(n_271),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_377),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_274),
.B(n_172),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_274),
.B(n_193),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_381),
.B(n_386),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_SL g387 ( 
.A(n_383),
.B(n_257),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_251),
.A2(n_192),
.B1(n_155),
.B2(n_147),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_387),
.A2(n_390),
.B(n_418),
.Y(n_442)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_323),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_388),
.B(n_408),
.Y(n_444)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_370),
.Y(n_391)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_391),
.Y(n_439)
);

O2A1O1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_326),
.A2(n_250),
.B(n_281),
.C(n_288),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_392),
.A2(n_402),
.B(n_432),
.Y(n_457)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_384),
.Y(n_393)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_393),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g394 ( 
.A(n_323),
.B(n_320),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_394),
.B(n_401),
.Y(n_449)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

INVx8_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_397),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_346),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g401 ( 
.A(n_333),
.B(n_314),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_351),
.A2(n_280),
.B(n_285),
.Y(n_402)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_379),
.Y(n_404)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_404),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_407),
.Y(n_462)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_409),
.A2(n_433),
.B1(n_329),
.B2(n_380),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_240),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_410),
.B(n_421),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_377),
.A2(n_192),
.B1(n_241),
.B2(n_247),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_412),
.A2(n_416),
.B1(n_372),
.B2(n_348),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_349),
.B(n_236),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_414),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_334),
.B(n_286),
.Y(n_414)
);

INVx13_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_415),
.Y(n_443)
);

OAI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_381),
.A2(n_302),
.B1(n_299),
.B2(n_319),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_347),
.B(n_301),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_420),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_419),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_350),
.B(n_256),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_327),
.B(n_321),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_429),
.Y(n_456)
);

OA22x2_ASAP7_75t_L g423 ( 
.A1(n_369),
.A2(n_239),
.B1(n_294),
.B2(n_295),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_423),
.B(n_425),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_325),
.A2(n_223),
.B(n_242),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_424),
.A2(n_389),
.B(n_411),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_368),
.B(n_297),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_358),
.B(n_242),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_427),
.C(n_434),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_328),
.B(n_223),
.C(n_155),
.Y(n_427)
);

INVx13_ASAP7_75t_L g428 ( 
.A(n_373),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_428),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_366),
.B(n_363),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_385),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_325),
.B(n_330),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_431),
.B(n_344),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_357),
.A2(n_354),
.B(n_340),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_369),
.A2(n_330),
.B1(n_337),
.B2(n_383),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_356),
.B(n_341),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_335),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_436),
.Y(n_463)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_342),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_331),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_437),
.B(n_448),
.C(n_451),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_440),
.B(n_452),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_432),
.A2(n_357),
.B1(n_329),
.B2(n_345),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_441),
.A2(n_454),
.B1(n_478),
.B2(n_412),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_402),
.A2(n_357),
.B(n_324),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_447),
.A2(n_450),
.B(n_459),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_418),
.A2(n_324),
.B(n_386),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_365),
.C(n_371),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_406),
.A2(n_352),
.B1(n_360),
.B2(n_344),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_424),
.A2(n_382),
.B(n_372),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_461),
.A2(n_465),
.B(n_475),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_393),
.B(n_371),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_469),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_392),
.A2(n_389),
.B(n_411),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_407),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_472),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_403),
.B(n_396),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_476),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_426),
.B(n_365),
.C(n_378),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_474),
.B(n_408),
.C(n_332),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_398),
.A2(n_348),
.B(n_378),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_420),
.B(n_385),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_405),
.A2(n_403),
.B1(n_413),
.B2(n_396),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_477),
.A2(n_479),
.B1(n_425),
.B2(n_400),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_405),
.A2(n_353),
.B1(n_359),
.B2(n_362),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_406),
.A2(n_359),
.B1(n_353),
.B2(n_362),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_459),
.Y(n_480)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_480),
.Y(n_523)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_481),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_482),
.A2(n_440),
.B1(n_450),
.B2(n_479),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_468),
.A2(n_398),
.B1(n_430),
.B2(n_434),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_483),
.A2(n_496),
.B1(n_444),
.B2(n_438),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_452),
.B(n_417),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_487),
.B(n_499),
.Y(n_528)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_488),
.Y(n_526)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_466),
.Y(n_489)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_489),
.Y(n_535)
);

BUFx5_ASAP7_75t_L g490 ( 
.A(n_439),
.Y(n_490)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_490),
.Y(n_545)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_439),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_494),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_457),
.A2(n_431),
.B(n_400),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_495),
.A2(n_515),
.B(n_516),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_468),
.A2(n_450),
.B1(n_454),
.B2(n_441),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_436),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_497),
.B(n_502),
.Y(n_548)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_463),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_498),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_445),
.B(n_429),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_463),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_500),
.B(n_508),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_449),
.B(n_401),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_445),
.B(n_332),
.Y(n_503)
);

CKINVDCx14_ASAP7_75t_R g549 ( 
.A(n_503),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_448),
.B(n_427),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_504),
.B(n_438),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_449),
.B(n_394),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_505),
.B(n_509),
.Y(n_551)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_469),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_506),
.A2(n_512),
.B1(n_514),
.B2(n_519),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_438),
.C(n_448),
.Y(n_530)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_476),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_464),
.B(n_423),
.Y(n_509)
);

CKINVDCx10_ASAP7_75t_R g510 ( 
.A(n_443),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_510),
.Y(n_525)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_446),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_511),
.B(n_518),
.Y(n_540)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_446),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_467),
.B(n_422),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_513),
.B(n_517),
.Y(n_547)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_453),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_457),
.A2(n_442),
.B(n_447),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_442),
.A2(n_397),
.B(n_423),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_455),
.B(n_339),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_455),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_478),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_423),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_520),
.B(n_475),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_521),
.A2(n_531),
.B1(n_537),
.B2(n_550),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_492),
.A2(n_480),
.B(n_501),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_524),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_510),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_527),
.B(n_534),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_530),
.B(n_542),
.C(n_556),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_496),
.A2(n_485),
.B1(n_482),
.B2(n_506),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_491),
.B(n_437),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_532),
.B(n_539),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_492),
.B(n_483),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_485),
.A2(n_479),
.B1(n_447),
.B2(n_458),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_498),
.B(n_458),
.Y(n_538)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_538),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_491),
.B(n_437),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_541),
.B(n_553),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_504),
.B(n_474),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_544),
.B(n_484),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_486),
.B(n_467),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_546),
.B(n_554),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_509),
.A2(n_465),
.B1(n_461),
.B2(n_474),
.Y(n_550)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_552),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_497),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_486),
.B(n_507),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_520),
.A2(n_472),
.B1(n_444),
.B2(n_456),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_555),
.A2(n_557),
.B1(n_481),
.B2(n_493),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_495),
.B(n_451),
.C(n_456),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_519),
.A2(n_451),
.B1(n_471),
.B2(n_460),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_515),
.B(n_453),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_558),
.B(n_364),
.C(n_367),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_543),
.A2(n_501),
.B(n_516),
.Y(n_560)
);

OAI21xp33_ASAP7_75t_L g604 ( 
.A1(n_560),
.A2(n_523),
.B(n_551),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_563),
.A2(n_567),
.B1(n_589),
.B2(n_553),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_564),
.B(n_591),
.Y(n_592)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_526),
.Y(n_565)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_565),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_521),
.A2(n_493),
.B1(n_484),
.B2(n_505),
.Y(n_567)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_536),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_568),
.B(n_569),
.Y(n_606)
);

OAI21xp33_ASAP7_75t_L g569 ( 
.A1(n_556),
.A2(n_493),
.B(n_502),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_522),
.A2(n_514),
.B1(n_488),
.B2(n_489),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_570),
.A2(n_587),
.B1(n_533),
.B2(n_527),
.Y(n_593)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_526),
.Y(n_574)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_574),
.Y(n_609)
);

OAI21xp33_ASAP7_75t_L g576 ( 
.A1(n_543),
.A2(n_470),
.B(n_443),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_576),
.B(n_577),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_528),
.B(n_470),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_542),
.B(n_512),
.C(n_404),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_578),
.B(n_580),
.C(n_585),
.Y(n_596)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_535),
.Y(n_579)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_579),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_532),
.B(n_395),
.C(n_391),
.Y(n_580)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_535),
.Y(n_582)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_582),
.Y(n_617)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_559),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_583),
.B(n_584),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_528),
.B(n_460),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_539),
.B(n_530),
.C(n_544),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_522),
.A2(n_494),
.B1(n_462),
.B2(n_419),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_550),
.B(n_382),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_588),
.B(n_590),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_531),
.A2(n_537),
.B1(n_555),
.B2(n_552),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_540),
.Y(n_590)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_593),
.Y(n_628)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_595),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_573),
.B(n_541),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_597),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_573),
.B(n_534),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_598),
.B(n_575),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_578),
.B(n_558),
.C(n_524),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_601),
.C(n_605),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_SL g600 ( 
.A(n_586),
.B(n_564),
.Y(n_600)
);

XNOR2x1_ASAP7_75t_L g618 ( 
.A(n_600),
.B(n_612),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_580),
.B(n_557),
.C(n_523),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_581),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_602),
.B(n_611),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_571),
.A2(n_562),
.B1(n_589),
.B2(n_563),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_603),
.A2(n_615),
.B1(n_583),
.B2(n_561),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_604),
.A2(n_588),
.B(n_570),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_585),
.B(n_586),
.C(n_591),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_572),
.B(n_548),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g635 ( 
.A(n_607),
.B(n_545),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_566),
.A2(n_548),
.B(n_551),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_608),
.B(n_587),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_567),
.A2(n_559),
.B1(n_529),
.B2(n_538),
.Y(n_611)
);

XOR2x2_ASAP7_75t_L g612 ( 
.A(n_588),
.B(n_547),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_562),
.A2(n_549),
.B1(n_533),
.B2(n_525),
.Y(n_615)
);

XNOR2x1_ASAP7_75t_L g644 ( 
.A(n_619),
.B(n_624),
.Y(n_644)
);

AOI21x1_ASAP7_75t_SL g621 ( 
.A1(n_610),
.A2(n_560),
.B(n_566),
.Y(n_621)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_621),
.Y(n_649)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_623),
.B(n_629),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_614),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_625),
.B(n_627),
.Y(n_642)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_626),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_615),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_596),
.B(n_525),
.C(n_579),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_611),
.B(n_582),
.Y(n_630)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_630),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_596),
.B(n_574),
.C(n_565),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_631),
.B(n_639),
.C(n_594),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_606),
.B(n_545),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_633),
.B(n_609),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_604),
.B(n_601),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_634),
.A2(n_598),
.B(n_612),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g640 ( 
.A(n_635),
.B(n_636),
.Y(n_640)
);

INVx13_ASAP7_75t_L g636 ( 
.A(n_593),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_616),
.B(n_490),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_637),
.A2(n_617),
.B(n_613),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_597),
.B(n_359),
.C(n_364),
.Y(n_639)
);

XOR2xp5_ASAP7_75t_L g641 ( 
.A(n_621),
.B(n_599),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_641),
.B(n_646),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_645),
.A2(n_648),
.B1(n_637),
.B2(n_619),
.Y(n_663)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_635),
.B(n_592),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_639),
.B(n_592),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_647),
.B(n_631),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_652),
.B(n_654),
.Y(n_660)
);

BUFx24_ASAP7_75t_SL g653 ( 
.A(n_625),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_653),
.B(n_629),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_633),
.B(n_607),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_655),
.A2(n_618),
.B(n_620),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_638),
.B(n_605),
.C(n_603),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_656),
.B(n_657),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_622),
.B(n_595),
.C(n_600),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_658),
.B(n_662),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_659),
.B(n_661),
.Y(n_672)
);

XOR2xp5_ASAP7_75t_L g661 ( 
.A(n_641),
.B(n_626),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_656),
.B(n_622),
.C(n_628),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_663),
.B(n_665),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_643),
.B(n_632),
.C(n_620),
.Y(n_665)
);

XOR2xp5_ASAP7_75t_L g666 ( 
.A(n_640),
.B(n_618),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_666),
.B(n_668),
.C(n_669),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_667),
.A2(n_644),
.B(n_646),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_657),
.B(n_632),
.C(n_628),
.Y(n_668)
);

XOR2xp5_ASAP7_75t_L g669 ( 
.A(n_640),
.B(n_624),
.Y(n_669)
);

MAJx2_ASAP7_75t_L g671 ( 
.A(n_670),
.B(n_649),
.C(n_642),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g681 ( 
.A(n_671),
.B(n_677),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_662),
.B(n_650),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_673),
.B(n_676),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_660),
.B(n_652),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_659),
.B(n_644),
.C(n_647),
.Y(n_679)
);

MAJIxp5_ASAP7_75t_L g682 ( 
.A(n_679),
.B(n_664),
.C(n_666),
.Y(n_682)
);

AOI322xp5_ASAP7_75t_L g680 ( 
.A1(n_678),
.A2(n_636),
.A3(n_651),
.B1(n_627),
.B2(n_664),
.C1(n_630),
.C2(n_661),
.Y(n_680)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_680),
.Y(n_686)
);

AOI21x1_ASAP7_75t_L g685 ( 
.A1(n_682),
.A2(n_684),
.B(n_672),
.Y(n_685)
);

NOR2x1_ASAP7_75t_L g684 ( 
.A(n_674),
.B(n_669),
.Y(n_684)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_685),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_SL g687 ( 
.A1(n_683),
.A2(n_672),
.B(n_675),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_687),
.B(n_682),
.C(n_684),
.Y(n_689)
);

MAJIxp5_ASAP7_75t_L g690 ( 
.A(n_689),
.B(n_686),
.C(n_681),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_690),
.A2(n_688),
.B1(n_636),
.B2(n_415),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_691),
.A2(n_428),
.B(n_339),
.Y(n_692)
);

AO21x2_ASAP7_75t_L g693 ( 
.A1(n_692),
.A2(n_343),
.B(n_367),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_693),
.B(n_343),
.Y(n_694)
);


endmodule