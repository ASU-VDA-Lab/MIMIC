module fake_jpeg_4483_n_319 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_37),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_11),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_40),
.B(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_35),
.B(n_16),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_33),
.C(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_50),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_19),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_49),
.B(n_35),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_20),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_17),
.B1(n_26),
.B2(n_22),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_64),
.B1(n_90),
.B2(n_97),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_25),
.B1(n_17),
.B2(n_26),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_25),
.B1(n_17),
.B2(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_58),
.B(n_65),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_25),
.B1(n_14),
.B2(n_34),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_87),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_14),
.B1(n_18),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_18),
.B1(n_22),
.B2(n_32),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_62),
.A2(n_68),
.B1(n_73),
.B2(n_78),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_63),
.A2(n_85),
.B(n_4),
.C(n_5),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_31),
.B1(n_29),
.B2(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_67),
.B(n_101),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_37),
.A2(n_28),
.B1(n_23),
.B2(n_30),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_76),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_37),
.A2(n_28),
.B1(n_23),
.B2(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_30),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_89),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_30),
.B1(n_35),
.B2(n_16),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_81),
.A2(n_86),
.B1(n_92),
.B2(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_38),
.B(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_39),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_0),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_43),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_102),
.Y(n_118)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_42),
.A2(n_8),
.B1(n_10),
.B2(n_3),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_8),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_42),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_64),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_112),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_72),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_110),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_77),
.Y(n_112)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_117),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_130),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_65),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_4),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_56),
.B(n_5),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_74),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_63),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_139),
.B(n_157),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_75),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_138),
.Y(n_171)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_143),
.Y(n_190)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_141),
.B(n_149),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_90),
.C(n_58),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_142),
.B(n_164),
.C(n_95),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_67),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_101),
.B(n_94),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_167),
.C(n_124),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_91),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_147),
.C(n_153),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_105),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_154),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_103),
.A2(n_69),
.B1(n_84),
.B2(n_66),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_156),
.B1(n_128),
.B2(n_93),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_60),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_166),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_103),
.A2(n_129),
.B1(n_104),
.B2(n_115),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_5),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_87),
.Y(n_161)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_56),
.C(n_83),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_165),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_104),
.B(n_71),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_122),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_169),
.B(n_175),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_SL g227 ( 
.A1(n_173),
.A2(n_177),
.B(n_186),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_107),
.B1(n_66),
.B2(n_69),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_200),
.B1(n_156),
.B2(n_154),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_107),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_112),
.B(n_117),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_162),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_179),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_84),
.B1(n_119),
.B2(n_131),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_184),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_163),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_128),
.B1(n_117),
.B2(n_112),
.C(n_113),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_185),
.A2(n_192),
.B(n_148),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_127),
.B1(n_159),
.B2(n_5),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_121),
.B(n_117),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_136),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_193),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_113),
.Y(n_194)
);

NOR2x1_ASAP7_75t_R g203 ( 
.A(n_194),
.B(n_149),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_143),
.B(n_98),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_202),
.C(n_137),
.Y(n_211)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_146),
.A2(n_95),
.B1(n_127),
.B2(n_102),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_155),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_206),
.B(n_208),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_190),
.B(n_194),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_210),
.B1(n_198),
.B2(n_172),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_209),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_148),
.B1(n_137),
.B2(n_141),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_219),
.C(n_168),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_212),
.B(n_215),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_157),
.B(n_160),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_214),
.A2(n_221),
.B1(n_227),
.B2(n_181),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_216),
.B(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_157),
.C(n_138),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_224),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_226),
.Y(n_233)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_241),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_234),
.B(n_240),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_175),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_229),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_246),
.C(n_249),
.Y(n_256)
);

AO22x1_ASAP7_75t_L g238 ( 
.A1(n_206),
.A2(n_177),
.B1(n_169),
.B2(n_188),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_252),
.B1(n_210),
.B2(n_217),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_239),
.A2(n_213),
.B1(n_205),
.B2(n_221),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_204),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_225),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_208),
.A2(n_168),
.B(n_176),
.C(n_177),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_170),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_211),
.C(n_228),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_209),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_250),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_201),
.C(n_170),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_236),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_261),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_235),
.B1(n_230),
.B2(n_248),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_242),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_239),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_267),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_213),
.C(n_219),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_264),
.C(n_237),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_214),
.C(n_207),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_266),
.B(n_269),
.Y(n_283)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_227),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_256),
.C(n_263),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_254),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_266),
.B1(n_257),
.B2(n_243),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_267),
.B1(n_230),
.B2(n_240),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_258),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_279),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_268),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_277),
.B(n_282),
.Y(n_287)
);

AOI221xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_232),
.B1(n_233),
.B2(n_244),
.C(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_265),
.A2(n_232),
.B(n_247),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_281),
.Y(n_286)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_284),
.B(n_272),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_294),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_256),
.C(n_249),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_293),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_257),
.C(n_253),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_259),
.C(n_251),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_295),
.A2(n_280),
.B(n_281),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_302),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_298),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_279),
.B1(n_283),
.B2(n_270),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_299),
.A2(n_294),
.B1(n_289),
.B2(n_284),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_222),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_287),
.A2(n_231),
.B(n_245),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_286),
.B(n_293),
.Y(n_305)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_224),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_292),
.B(n_217),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_308),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_312),
.A2(n_309),
.B1(n_300),
.B2(n_306),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_314),
.A2(n_315),
.B(n_305),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_310),
.C(n_296),
.Y(n_315)
);

AOI21x1_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_311),
.B(n_304),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_318),
.Y(n_319)
);


endmodule