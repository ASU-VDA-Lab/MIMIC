module fake_jpeg_14564_n_355 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_355);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_10),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_10),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_54),
.B(n_31),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_59),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_22),
.B1(n_26),
.B2(n_29),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_73),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_68),
.A2(n_35),
.B1(n_33),
.B2(n_31),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_76),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_82),
.Y(n_120)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_85),
.Y(n_108)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_42),
.B(n_32),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_61),
.B(n_42),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_98),
.B(n_37),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_104),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_38),
.C(n_21),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_121),
.C(n_39),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_22),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_26),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_115),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_88),
.Y(n_146)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_62),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_124),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_65),
.A2(n_25),
.B1(n_35),
.B2(n_33),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_65),
.B1(n_85),
.B2(n_69),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_38),
.C(n_27),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_79),
.A2(n_59),
.B1(n_83),
.B2(n_69),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_67),
.B1(n_92),
.B2(n_71),
.Y(n_129)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx12_ASAP7_75t_R g124 ( 
.A(n_62),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_30),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_144),
.B1(n_149),
.B2(n_113),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_33),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_148),
.C(n_154),
.Y(n_162)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_35),
.B1(n_59),
.B2(n_30),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_151),
.B1(n_96),
.B2(n_108),
.Y(n_159)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_139),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_94),
.CI(n_86),
.CON(n_139),
.SN(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_37),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_146),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_34),
.B1(n_56),
.B2(n_3),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_57),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_1),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_107),
.B1(n_97),
.B2(n_32),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_112),
.A2(n_121),
.B1(n_102),
.B2(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_66),
.C(n_70),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_157),
.Y(n_178)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_111),
.B1(n_110),
.B2(n_103),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_66),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_159),
.A2(n_161),
.B1(n_163),
.B2(n_169),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_156),
.A2(n_108),
.B1(n_96),
.B2(n_103),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_164),
.B(n_155),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_122),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_166),
.A2(n_174),
.B(n_145),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_110),
.B1(n_113),
.B2(n_99),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_127),
.C(n_100),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_129),
.C(n_100),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_172),
.A2(n_146),
.B1(n_134),
.B2(n_154),
.Y(n_192)
);

AO22x1_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_93),
.B1(n_84),
.B2(n_72),
.Y(n_175)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_173),
.B1(n_170),
.B2(n_141),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_145),
.B1(n_149),
.B2(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_180),
.A2(n_185),
.B1(n_172),
.B2(n_164),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_183),
.B(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_177),
.B(n_137),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_197),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_137),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_191),
.C(n_196),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_139),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_196),
.B1(n_198),
.B2(n_181),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_159),
.B(n_150),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_198),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_150),
.B(n_140),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_195),
.B(n_178),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_166),
.A2(n_152),
.B(n_147),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

XNOR2x1_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_128),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_200),
.B(n_41),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_205),
.B1(n_207),
.B2(n_41),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_209),
.B(n_220),
.Y(n_227)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_174),
.B1(n_178),
.B2(n_165),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_177),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_143),
.C(n_27),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_168),
.B1(n_173),
.B2(n_167),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_138),
.B(n_176),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_195),
.B1(n_185),
.B2(n_192),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_135),
.B1(n_141),
.B2(n_170),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_40),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_131),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_217),
.B(n_153),
.Y(n_229)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_2),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_183),
.A2(n_167),
.B(n_160),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_160),
.B(n_34),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_220),
.B(n_210),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_133),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_2),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_170),
.B1(n_143),
.B2(n_133),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_237),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_214),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_228),
.B(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_234),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_84),
.C(n_95),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_235),
.C(n_201),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_210),
.B(n_41),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_38),
.C(n_27),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_206),
.B(n_41),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_245),
.B1(n_230),
.B2(n_216),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_242),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_224),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_246),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_246),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_252),
.C(n_253),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_219),
.C(n_222),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_199),
.B1(n_219),
.B2(n_215),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_231),
.B1(n_223),
.B2(n_228),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_209),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_260),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_214),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_200),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_260),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_225),
.B(n_204),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_221),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_264),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_211),
.C(n_212),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_253),
.C(n_252),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_268),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_238),
.B(n_231),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_277),
.B(n_249),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_254),
.B(n_226),
.CI(n_236),
.CON(n_273),
.SN(n_273)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_286),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_287),
.C(n_258),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_276),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_251),
.B(n_258),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_285),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_241),
.B1(n_8),
.B2(n_9),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_247),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_241),
.C(n_8),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_289),
.B(n_283),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_250),
.C(n_263),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_297),
.Y(n_305)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_302),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_265),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_271),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_255),
.C(n_256),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_7),
.C(n_10),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_287),
.B(n_278),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_7),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_7),
.Y(n_310)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_270),
.B(n_273),
.Y(n_302)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_283),
.Y(n_313)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_306)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_307),
.B(n_311),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_285),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_288),
.C(n_293),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_313),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_303),
.A2(n_273),
.B1(n_269),
.B2(n_279),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_314),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_291),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_12),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_295),
.B(n_14),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_301),
.B(n_299),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_319),
.A2(n_302),
.B(n_294),
.C(n_314),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_20),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_308),
.C(n_292),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_301),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_325),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_309),
.A2(n_302),
.B(n_300),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_312),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_331),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_330),
.B(n_334),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_332),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_14),
.C(n_15),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_323),
.C(n_17),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_16),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_335),
.A2(n_337),
.B(n_16),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_325),
.B(n_318),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_336),
.B(n_328),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_339),
.B(n_340),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_320),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_344),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_338),
.A2(n_16),
.B(n_17),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_347),
.Y(n_349)
);

BUFx4f_ASAP7_75t_SL g348 ( 
.A(n_341),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_348),
.B(n_339),
.C(n_343),
.Y(n_350)
);

AO21x1_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_346),
.B(n_345),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_349),
.Y(n_352)
);

AOI221xp5_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.C(n_343),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_18),
.C(n_19),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_SL g355 ( 
.A(n_354),
.B(n_18),
.Y(n_355)
);


endmodule