module fake_netlist_6_2784_n_2052 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2052);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2052;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_175),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_46),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

HB1xp67_ASAP7_75t_SL g205 ( 
.A(n_33),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_53),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_16),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_1),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_94),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_59),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_66),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_19),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_108),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_112),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_33),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_185),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_6),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_106),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_173),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_147),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_116),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_148),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_77),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_165),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_43),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_122),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_63),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_74),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_59),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_60),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_111),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_29),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_92),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_85),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_5),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_57),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_145),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_109),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_52),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_155),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_36),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_21),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_34),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_102),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_150),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_129),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_53),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_16),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_131),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_35),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_3),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_24),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_75),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_49),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_68),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_158),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_104),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_115),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_154),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_56),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_13),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_132),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_188),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_127),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_113),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_64),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_0),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_26),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_17),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_164),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_3),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_177),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_72),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_64),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_67),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_72),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_199),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_50),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_176),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_62),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_76),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_128),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_74),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_121),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_13),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_96),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_80),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_58),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_82),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_5),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_69),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_123),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_191),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_73),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_45),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_57),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_126),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_7),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_180),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_2),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_160),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_49),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_90),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_100),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_118),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_71),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_35),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_83),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_10),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_182),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_6),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_44),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_149),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_66),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_14),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_20),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_55),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_91),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_163),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_36),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_186),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_124),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_139),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_23),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_17),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_60),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_76),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_58),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_69),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_51),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_138),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_107),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_79),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_29),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_63),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_87),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_197),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_189),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_28),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_26),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_50),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_37),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_88),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_39),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_179),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_168),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_93),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_153),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_125),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_62),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_192),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_11),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_170),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_130),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_161),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_171),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_166),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_114),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_143),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_75),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_4),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_4),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_14),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_174),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_151),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_120),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_21),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_37),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_146),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_156),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_39),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_48),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_81),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_97),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_7),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_32),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_200),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_51),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_41),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_190),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_71),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_9),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_136),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_43),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_45),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_99),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_20),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_46),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_194),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_119),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_198),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_98),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_32),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_61),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_324),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_231),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_254),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_256),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_237),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_258),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_259),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_260),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_284),
.B(n_0),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_284),
.B(n_1),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_261),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_316),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_238),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_267),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_238),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_266),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_243),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_278),
.B(n_2),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_263),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_363),
.B(n_8),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_264),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_221),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_272),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_306),
.B(n_8),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_238),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_273),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_238),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_238),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_253),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_253),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_253),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_296),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_282),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_205),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_310),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_253),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_R g439 ( 
.A(n_201),
.B(n_9),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_327),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_274),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_253),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_307),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_283),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_283),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_275),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_281),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_283),
.Y(n_448)
);

INVxp33_ASAP7_75t_SL g449 ( 
.A(n_206),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_221),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_287),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_218),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_283),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_288),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_297),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_283),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_203),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_242),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_248),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_298),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_285),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_301),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_311),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_292),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_295),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_302),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_320),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_325),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_255),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_305),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_303),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_309),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_322),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_206),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_262),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_334),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_367),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_313),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_369),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_245),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_268),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_314),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_270),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_375),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_382),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_383),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_319),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_389),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_277),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_269),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_269),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_304),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_331),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_332),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_304),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_333),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_336),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_337),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_279),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_286),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_245),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_361),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_361),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_204),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_245),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_289),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_306),
.B(n_10),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_342),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_207),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_346),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_347),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_210),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_209),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_349),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_226),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_401),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_232),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_209),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_469),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_475),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_442),
.Y(n_524)
);

AO22x1_ASAP7_75t_L g525 ( 
.A1(n_426),
.A2(n_378),
.B1(n_318),
.B2(n_335),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_403),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_442),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_436),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_481),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_492),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_415),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_402),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_417),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_424),
.B(n_290),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_421),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_483),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_R g537 ( 
.A(n_490),
.B(n_291),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_427),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_407),
.B(n_362),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_402),
.B(n_452),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_421),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_502),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_429),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_503),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_405),
.B(n_213),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_421),
.Y(n_547)
);

AND2x2_ASAP7_75t_R g548 ( 
.A(n_439),
.B(n_239),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_431),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_421),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_508),
.B(n_344),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_432),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_509),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_433),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_492),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_438),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_444),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_406),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_448),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_507),
.B(n_362),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_406),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_408),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_408),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_409),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_409),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_450),
.B(n_494),
.Y(n_567)
);

NOR2xp67_ASAP7_75t_L g568 ( 
.A(n_495),
.B(n_240),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_453),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_498),
.B(n_212),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_456),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_521),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_512),
.B(n_201),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_419),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_457),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_515),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_458),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_518),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_410),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_SL g580 ( 
.A(n_420),
.B(n_290),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_413),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_459),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_461),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_464),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_413),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_465),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_418),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_418),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_R g589 ( 
.A(n_425),
.B(n_294),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_425),
.B(n_344),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_520),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_435),
.A2(n_388),
.B1(n_359),
.B2(n_348),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_471),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_472),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_473),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_423),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_476),
.Y(n_597)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_505),
.B(n_252),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_506),
.B(n_404),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_477),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_414),
.B(n_212),
.Y(n_601)
);

OA21x2_ASAP7_75t_L g602 ( 
.A1(n_411),
.A2(n_250),
.B(n_216),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_428),
.B(n_344),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_428),
.B(n_350),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_479),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_484),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_412),
.A2(n_250),
.B(n_216),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_485),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_486),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_441),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_487),
.B(n_318),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_567),
.B(n_516),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_567),
.B(n_446),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_552),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_539),
.B(n_276),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_592),
.B(n_474),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_573),
.B(n_449),
.Y(n_617)
);

AND3x2_ASAP7_75t_L g618 ( 
.A(n_532),
.B(n_422),
.C(n_510),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_550),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_573),
.B(n_449),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_530),
.B(n_276),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_534),
.B(n_330),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_572),
.B(n_446),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_575),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_535),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_550),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_537),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_550),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_575),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_572),
.B(n_447),
.Y(n_630)
);

INVx6_ASAP7_75t_L g631 ( 
.A(n_530),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_577),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_555),
.B(n_330),
.Y(n_633)
);

BUFx4f_ASAP7_75t_L g634 ( 
.A(n_579),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_555),
.B(n_451),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_577),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_589),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_534),
.B(n_451),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_525),
.B(n_454),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_525),
.B(n_455),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_582),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_531),
.B(n_455),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_552),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_531),
.B(n_460),
.Y(n_644)
);

OAI21xp33_ASAP7_75t_SL g645 ( 
.A1(n_607),
.A2(n_374),
.B(n_335),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_608),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_582),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_599),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_592),
.B(n_443),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_528),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_533),
.B(n_460),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_583),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_533),
.B(n_462),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_590),
.B(n_462),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_611),
.B(n_343),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_550),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_608),
.B(n_355),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_557),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_608),
.B(n_355),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_608),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_583),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_597),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_557),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_603),
.B(n_470),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_597),
.B(n_371),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_584),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_547),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_522),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_532),
.B(n_480),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_597),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_584),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_586),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_586),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_535),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_547),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_611),
.B(n_489),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_609),
.B(n_371),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_535),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_538),
.B(n_470),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_593),
.Y(n_680)
);

BUFx4f_ASAP7_75t_L g681 ( 
.A(n_579),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_580),
.B(n_263),
.Y(n_682)
);

CKINVDCx16_ASAP7_75t_R g683 ( 
.A(n_526),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_541),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_557),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_593),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_541),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_594),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_560),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_546),
.B(n_482),
.C(n_478),
.Y(n_690)
);

AND2x2_ASAP7_75t_SL g691 ( 
.A(n_602),
.B(n_263),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_538),
.B(n_478),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_602),
.A2(n_257),
.B1(n_230),
.B2(n_341),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_L g694 ( 
.A(n_559),
.B(n_519),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_594),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_604),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_574),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_541),
.Y(n_698)
);

AND2x6_ASAP7_75t_L g699 ( 
.A(n_540),
.B(n_263),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_595),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_595),
.B(n_491),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_602),
.A2(n_341),
.B1(n_230),
.B2(n_208),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_543),
.B(n_545),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_551),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_605),
.B(n_263),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_543),
.B(n_482),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_605),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_606),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_560),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_562),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_606),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_576),
.B(n_271),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_547),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_563),
.B(n_488),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_545),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_561),
.B(n_488),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_602),
.A2(n_257),
.B1(n_208),
.B2(n_211),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_564),
.A2(n_497),
.B1(n_517),
.B2(n_514),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_549),
.B(n_496),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_607),
.A2(n_211),
.B1(n_374),
.B2(n_440),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_576),
.B(n_271),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_561),
.A2(n_466),
.B1(n_213),
.B2(n_351),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_549),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_570),
.B(n_497),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_554),
.B(n_499),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_554),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_556),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_565),
.B(n_499),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_556),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_558),
.B(n_500),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_578),
.B(n_271),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_547),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_560),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_601),
.A2(n_416),
.B1(n_493),
.B2(n_293),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_578),
.B(n_271),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_558),
.Y(n_736)
);

AO22x2_ASAP7_75t_L g737 ( 
.A1(n_548),
.A2(n_373),
.B1(n_397),
.B2(n_265),
.Y(n_737)
);

INVx5_ASAP7_75t_L g738 ( 
.A(n_547),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_569),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_596),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_569),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_566),
.A2(n_214),
.B1(n_215),
.B2(n_219),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_571),
.B(n_500),
.Y(n_743)
);

AND2x2_ASAP7_75t_SL g744 ( 
.A(n_548),
.B(n_271),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_591),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_591),
.B(n_501),
.Y(n_746)
);

OR2x6_ASAP7_75t_L g747 ( 
.A(n_600),
.B(n_504),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_571),
.B(n_501),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_568),
.B(n_511),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_617),
.B(n_581),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_617),
.B(n_620),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_661),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_620),
.B(n_585),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_638),
.B(n_587),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_661),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_638),
.A2(n_568),
.B(n_598),
.C(n_317),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_680),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_680),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_700),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_691),
.A2(n_547),
.B(n_591),
.Y(n_760)
);

NOR2x1p5_ASAP7_75t_L g761 ( 
.A(n_627),
.B(n_588),
.Y(n_761)
);

INVxp33_ASAP7_75t_SL g762 ( 
.A(n_668),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_716),
.B(n_610),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_724),
.B(n_670),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_700),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_624),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_693),
.A2(n_323),
.B1(n_228),
.B2(n_321),
.Y(n_767)
);

OAI21xp33_ASAP7_75t_L g768 ( 
.A1(n_654),
.A2(n_513),
.B(n_215),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_629),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_744),
.B(n_293),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_724),
.B(n_744),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_632),
.Y(n_772)
);

INVx8_ASAP7_75t_L g773 ( 
.A(n_747),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_696),
.B(n_293),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_636),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_639),
.B(n_244),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_640),
.B(n_746),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_622),
.B(n_312),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_641),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_622),
.B(n_315),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_622),
.B(n_326),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_623),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_647),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_613),
.B(n_308),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_642),
.B(n_366),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_644),
.B(n_202),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_652),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_674),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_622),
.B(n_345),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_654),
.A2(n_434),
.B1(n_468),
.B2(n_467),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_631),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_612),
.B(n_523),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_614),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_666),
.Y(n_794)
);

BUFx5_ASAP7_75t_L g795 ( 
.A(n_691),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_614),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_697),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_622),
.B(n_662),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_699),
.B(n_299),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_664),
.B(n_536),
.C(n_529),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_671),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_651),
.B(n_202),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_672),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_747),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_662),
.B(n_364),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_664),
.B(n_542),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_693),
.A2(n_280),
.B1(n_293),
.B2(n_339),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_737),
.A2(n_437),
.B1(n_463),
.B2(n_300),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_653),
.B(n_217),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_740),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_630),
.Y(n_811)
);

NOR2xp67_ASAP7_75t_L g812 ( 
.A(n_690),
.B(n_718),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_637),
.B(n_544),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_676),
.Y(n_814)
);

NOR3xp33_ASAP7_75t_L g815 ( 
.A(n_704),
.B(n_553),
.C(n_219),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_702),
.A2(n_293),
.B1(n_339),
.B2(n_396),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_616),
.B(n_214),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_673),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_650),
.B(n_600),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_648),
.B(n_600),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_674),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_643),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_686),
.B(n_393),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_725),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_676),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_679),
.B(n_217),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_688),
.B(n_524),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_695),
.B(n_524),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_655),
.A2(n_328),
.B1(n_329),
.B2(n_338),
.Y(n_829)
);

NAND3xp33_ASAP7_75t_L g830 ( 
.A(n_725),
.B(n_353),
.C(n_223),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_702),
.B(n_717),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_631),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_707),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_708),
.B(n_527),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_711),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_655),
.A2(n_340),
.B1(n_399),
.B2(n_398),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_692),
.B(n_220),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_648),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_SL g839 ( 
.A1(n_634),
.A2(n_350),
.B1(n_222),
.B2(n_233),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_SL g840 ( 
.A(n_634),
.B(n_350),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_715),
.B(n_339),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_SL g842 ( 
.A(n_714),
.B(n_222),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_706),
.B(n_223),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_723),
.B(n_339),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_726),
.B(n_339),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_645),
.A2(n_356),
.B(n_399),
.C(n_398),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_719),
.B(n_224),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_727),
.B(n_224),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_L g849 ( 
.A(n_694),
.B(n_400),
.C(n_392),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_730),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_729),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_743),
.B(n_225),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_736),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_739),
.B(n_227),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_741),
.B(n_227),
.Y(n_855)
);

CKINVDCx11_ASAP7_75t_R g856 ( 
.A(n_710),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_748),
.B(n_229),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_SL g858 ( 
.A1(n_683),
.A2(n_400),
.B1(n_392),
.B2(n_391),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_655),
.A2(n_356),
.B1(n_390),
.B2(n_387),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_655),
.A2(n_354),
.B1(n_390),
.B2(n_387),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_L g861 ( 
.A(n_699),
.B(n_229),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_747),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_615),
.A2(n_391),
.B1(n_386),
.B2(n_234),
.Y(n_863)
);

OAI22x1_ASAP7_75t_SL g864 ( 
.A1(n_742),
.A2(n_386),
.B1(n_234),
.B2(n_235),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_681),
.Y(n_865)
);

OAI22xp33_ASAP7_75t_L g866 ( 
.A1(n_649),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_728),
.B(n_236),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_701),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_703),
.A2(n_633),
.B(n_621),
.Y(n_869)
);

OAI22x1_ASAP7_75t_SL g870 ( 
.A1(n_742),
.A2(n_241),
.B1(n_247),
.B2(n_249),
.Y(n_870)
);

OAI22xp33_ASAP7_75t_L g871 ( 
.A1(n_722),
.A2(n_241),
.B1(n_247),
.B2(n_249),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_720),
.A2(n_351),
.B1(n_357),
.B2(n_368),
.Y(n_872)
);

NOR2x1p5_ASAP7_75t_L g873 ( 
.A(n_749),
.B(n_357),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_658),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_663),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_701),
.Y(n_876)
);

NOR2xp67_ASAP7_75t_L g877 ( 
.A(n_635),
.B(n_246),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_745),
.B(n_251),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_674),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_720),
.A2(n_368),
.B1(n_370),
.B2(n_379),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_681),
.B(n_251),
.Y(n_881)
);

NAND2x1_ASAP7_75t_L g882 ( 
.A(n_619),
.B(n_78),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_745),
.B(n_352),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_635),
.A2(n_384),
.B1(n_381),
.B2(n_380),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_655),
.B(n_352),
.Y(n_885)
);

AND2x2_ASAP7_75t_SL g886 ( 
.A(n_734),
.B(n_84),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_674),
.B(n_353),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_621),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_633),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_SL g890 ( 
.A(n_682),
.B(n_370),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_699),
.B(n_354),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_663),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_831),
.A2(n_665),
.B(n_677),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_876),
.B(n_682),
.Y(n_894)
);

BUFx4f_ASAP7_75t_L g895 ( 
.A(n_773),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_811),
.B(n_710),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_831),
.B(n_618),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_771),
.A2(n_734),
.B1(n_669),
.B2(n_677),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_816),
.A2(n_646),
.B(n_660),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_777),
.B(n_722),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_816),
.A2(n_646),
.B(n_660),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_777),
.B(n_358),
.Y(n_902)
);

CKINVDCx10_ASAP7_75t_R g903 ( 
.A(n_856),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_795),
.B(n_618),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_824),
.B(n_358),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_820),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_850),
.B(n_360),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_SL g908 ( 
.A(n_762),
.B(n_669),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_793),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_782),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_764),
.A2(n_628),
.B(n_626),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_795),
.B(n_685),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_760),
.A2(n_628),
.B(n_626),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_869),
.A2(n_659),
.B(n_657),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_795),
.B(n_685),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_751),
.A2(n_699),
.B1(n_665),
.B2(n_657),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_795),
.B(n_689),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_753),
.B(n_360),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_797),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_838),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_795),
.B(n_689),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_795),
.B(n_709),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_886),
.B(n_709),
.Y(n_923)
);

AOI21x1_ASAP7_75t_L g924 ( 
.A1(n_805),
.A2(n_687),
.B(n_625),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_819),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_819),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_753),
.B(n_365),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_810),
.Y(n_928)
);

AND2x4_ASAP7_75t_SL g929 ( 
.A(n_819),
.B(n_678),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_791),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_886),
.B(n_733),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_766),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_867),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_785),
.B(n_365),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_770),
.A2(n_699),
.B(n_735),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_778),
.A2(n_656),
.B(n_675),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_796),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_780),
.A2(n_656),
.B(n_675),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_791),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_770),
.A2(n_731),
.B(n_721),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_781),
.A2(n_738),
.B(n_667),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_776),
.A2(n_731),
.B(n_721),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_791),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_784),
.B(n_379),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_785),
.B(n_733),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_789),
.A2(n_738),
.B(n_667),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_879),
.A2(n_738),
.B(n_667),
.Y(n_947)
);

OR2x6_ASAP7_75t_SL g948 ( 
.A(n_817),
.B(n_372),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_769),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_772),
.Y(n_950)
);

NOR2xp67_ASAP7_75t_L g951 ( 
.A(n_865),
.B(n_712),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_788),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_784),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_750),
.B(n_372),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_812),
.A2(n_684),
.B1(n_678),
.B2(n_698),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_807),
.A2(n_712),
.B1(n_377),
.B2(n_380),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_807),
.A2(n_376),
.B1(n_377),
.B2(n_381),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_822),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_888),
.B(n_684),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_827),
.A2(n_678),
.B(n_698),
.Y(n_960)
);

OAI321xp33_ASAP7_75t_L g961 ( 
.A1(n_871),
.A2(n_11),
.A3(n_12),
.B1(n_15),
.B2(n_18),
.C(n_19),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_889),
.A2(n_705),
.B(n_376),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_832),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_775),
.Y(n_964)
);

CKINVDCx10_ASAP7_75t_R g965 ( 
.A(n_864),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_786),
.B(n_678),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_786),
.B(n_698),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_879),
.A2(n_738),
.B(n_667),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_879),
.A2(n_675),
.B(n_713),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_788),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_873),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_879),
.A2(n_732),
.B(n_713),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_779),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_763),
.B(n_384),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_763),
.B(n_698),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_767),
.B(n_12),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_842),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_783),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_787),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_773),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_885),
.A2(n_732),
.B(n_713),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_882),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_821),
.B(n_732),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_821),
.A2(n_732),
.B(n_713),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_802),
.A2(n_705),
.B(n_22),
.C(n_23),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_767),
.A2(n_705),
.B1(n_103),
.B2(n_105),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_840),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_809),
.B(n_705),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_874),
.A2(n_101),
.B(n_195),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_875),
.A2(n_95),
.B(n_187),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_814),
.B(n_825),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_826),
.A2(n_89),
.B1(n_184),
.B2(n_183),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_773),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_892),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_799),
.A2(n_196),
.B(n_181),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_826),
.B(n_172),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_861),
.A2(n_169),
.B(n_162),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_877),
.B(n_157),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_837),
.B(n_843),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_843),
.A2(n_141),
.B1(n_140),
.B2(n_137),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_847),
.B(n_135),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_847),
.B(n_852),
.Y(n_1002)
);

NOR2x1_ASAP7_75t_L g1003 ( 
.A(n_813),
.B(n_134),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_852),
.B(n_133),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_794),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_857),
.B(n_110),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_857),
.B(n_117),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_801),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_803),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_792),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_818),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_754),
.B(n_25),
.Y(n_1012)
);

AND2x2_ASAP7_75t_SL g1013 ( 
.A(n_790),
.B(n_27),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_SL g1014 ( 
.A1(n_756),
.A2(n_27),
.B(n_28),
.C(n_30),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_752),
.B(n_30),
.Y(n_1015)
);

NOR2x1p5_ASAP7_75t_SL g1016 ( 
.A(n_833),
.B(n_31),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_878),
.A2(n_31),
.B(n_34),
.Y(n_1017)
);

CKINVDCx10_ASAP7_75t_R g1018 ( 
.A(n_870),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_768),
.A2(n_835),
.B(n_851),
.C(n_853),
.Y(n_1019)
);

NAND2x1p5_ASAP7_75t_L g1020 ( 
.A(n_755),
.B(n_38),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_828),
.A2(n_38),
.B(n_40),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_757),
.B(n_40),
.Y(n_1022)
);

AO21x1_ASAP7_75t_L g1023 ( 
.A1(n_887),
.A2(n_41),
.B(n_42),
.Y(n_1023)
);

INVx11_ASAP7_75t_L g1024 ( 
.A(n_890),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_834),
.A2(n_42),
.B(n_44),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_758),
.B(n_759),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_765),
.A2(n_47),
.B(n_48),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_868),
.B(n_47),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_830),
.A2(n_77),
.B(n_54),
.C(n_55),
.Y(n_1029)
);

INVx3_ASAP7_75t_SL g1030 ( 
.A(n_806),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_887),
.A2(n_52),
.B(n_54),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_804),
.Y(n_1032)
);

CKINVDCx10_ASAP7_75t_R g1033 ( 
.A(n_858),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_804),
.B(n_73),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_823),
.A2(n_61),
.B(n_65),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_891),
.A2(n_65),
.B(n_67),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_841),
.A2(n_70),
.B(n_845),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_844),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_839),
.B(n_70),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_848),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_859),
.A2(n_860),
.B1(n_836),
.B2(n_862),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_829),
.A2(n_855),
.B(n_854),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_774),
.A2(n_883),
.B(n_881),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_872),
.B(n_880),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_883),
.A2(n_881),
.B(n_884),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_862),
.B(n_866),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_866),
.B(n_808),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_849),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_815),
.A2(n_800),
.B(n_863),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_863),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_872),
.A2(n_880),
.B(n_871),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_771),
.A2(n_751),
.B1(n_777),
.B2(n_886),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_791),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_831),
.A2(n_816),
.B(n_798),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_820),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_831),
.A2(n_816),
.B(n_798),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_925),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_999),
.A2(n_1002),
.B(n_1051),
.C(n_1047),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_999),
.B(n_1002),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_919),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1054),
.A2(n_1056),
.B(n_967),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_897),
.A2(n_1052),
.B(n_893),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_944),
.B(n_953),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_897),
.A2(n_931),
.B(n_923),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1040),
.B(n_945),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_980),
.B(n_993),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_945),
.B(n_906),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_909),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_933),
.B(n_896),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_937),
.Y(n_1070)
);

NOR2xp67_ASAP7_75t_SL g1071 ( 
.A(n_961),
.B(n_976),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1055),
.B(n_1044),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_918),
.A2(n_927),
.B(n_1045),
.C(n_1044),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_932),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_949),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_924),
.A2(n_911),
.B(n_981),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_974),
.A2(n_900),
.B1(n_904),
.B2(n_1048),
.Y(n_1077)
);

AOI221x1_ASAP7_75t_L g1078 ( 
.A1(n_1049),
.A2(n_1001),
.B1(n_1007),
.B2(n_1006),
.C(n_1004),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_993),
.Y(n_1079)
);

NAND2x1_ASAP7_75t_L g1080 ( 
.A(n_952),
.B(n_970),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_926),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_966),
.A2(n_901),
.B(n_899),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1050),
.B(n_923),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1009),
.B(n_975),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_904),
.A2(n_954),
.B1(n_1012),
.B2(n_1041),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1009),
.B(n_912),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_913),
.A2(n_915),
.B(n_912),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_915),
.A2(n_922),
.B(n_921),
.Y(n_1088)
);

CKINVDCx11_ASAP7_75t_R g1089 ( 
.A(n_948),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_934),
.A2(n_1010),
.B1(n_894),
.B2(n_1004),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_910),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_930),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_980),
.B(n_993),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_917),
.A2(n_921),
.B(n_922),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_987),
.B(n_1030),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_984),
.A2(n_972),
.B(n_959),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_959),
.A2(n_983),
.B(n_940),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_903),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1001),
.A2(n_1007),
.B(n_1006),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1042),
.A2(n_935),
.B(n_988),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_936),
.A2(n_938),
.B(n_969),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1043),
.A2(n_916),
.B(n_942),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_941),
.A2(n_946),
.B(n_955),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_928),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_930),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_950),
.B(n_964),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_973),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_978),
.B(n_979),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1005),
.B(n_1019),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_939),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_898),
.A2(n_986),
.B(n_962),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_989),
.A2(n_990),
.B(n_995),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_1024),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_905),
.B(n_907),
.Y(n_1114)
);

NAND2x1p5_ASAP7_75t_L g1115 ( 
.A(n_1053),
.B(n_895),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_939),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1026),
.B(n_994),
.Y(n_1117)
);

AOI21x1_ASAP7_75t_L g1118 ( 
.A1(n_998),
.A2(n_951),
.B(n_958),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1028),
.A2(n_956),
.B(n_1046),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_997),
.A2(n_982),
.B(n_894),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_1034),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_977),
.B(n_902),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1028),
.A2(n_1031),
.B(n_1037),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_920),
.Y(n_1124)
);

OR2x6_ASAP7_75t_L g1125 ( 
.A(n_963),
.B(n_1032),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_943),
.B(n_1013),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_947),
.A2(n_968),
.B(n_1025),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_908),
.B(n_963),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_1023),
.A2(n_985),
.A3(n_1029),
.B(n_1036),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_963),
.B(n_991),
.Y(n_1130)
);

AO21x2_ASAP7_75t_L g1131 ( 
.A1(n_992),
.A2(n_1000),
.B(n_1017),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1003),
.A2(n_1027),
.B(n_1021),
.Y(n_1132)
);

AOI21xp33_ASAP7_75t_L g1133 ( 
.A1(n_957),
.A2(n_1039),
.B(n_1008),
.Y(n_1133)
);

INVx3_ASAP7_75t_SL g1134 ( 
.A(n_971),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_991),
.B(n_895),
.Y(n_1135)
);

AND3x4_ASAP7_75t_L g1136 ( 
.A(n_1033),
.B(n_965),
.C(n_1018),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_939),
.B(n_929),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1053),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_982),
.A2(n_1015),
.B(n_1022),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1020),
.A2(n_1035),
.B1(n_1014),
.B2(n_1016),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1020),
.A2(n_960),
.B(n_914),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_999),
.B(n_1002),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_944),
.B(n_811),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_944),
.B(n_811),
.Y(n_1144)
);

INVx4_ASAP7_75t_L g1145 ( 
.A(n_993),
.Y(n_1145)
);

AOI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_999),
.A2(n_1002),
.B(n_751),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1054),
.A2(n_1056),
.B(n_897),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_999),
.B(n_1002),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1011),
.Y(n_1149)
);

AOI22x1_ASAP7_75t_L g1150 ( 
.A1(n_1043),
.A2(n_942),
.B1(n_1042),
.B2(n_1038),
.Y(n_1150)
);

NOR2x1_ASAP7_75t_SL g1151 ( 
.A(n_998),
.B(n_831),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_944),
.B(n_811),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1054),
.A2(n_831),
.B(n_816),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_999),
.B(n_1002),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_944),
.B(n_811),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_999),
.B(n_1002),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_932),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_999),
.B(n_1002),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_999),
.A2(n_1002),
.B(n_1051),
.C(n_1047),
.Y(n_1159)
);

OAI22x1_ASAP7_75t_L g1160 ( 
.A1(n_1047),
.A2(n_751),
.B1(n_753),
.B2(n_976),
.Y(n_1160)
);

AND2x6_ASAP7_75t_L g1161 ( 
.A(n_976),
.B(n_923),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_910),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1054),
.A2(n_831),
.B(n_816),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_993),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1011),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_925),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_896),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_993),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_999),
.B(n_1002),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_993),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1054),
.A2(n_1056),
.B(n_897),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_999),
.B(n_1002),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_993),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_999),
.A2(n_1002),
.B1(n_918),
.B2(n_927),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_999),
.A2(n_751),
.B(n_1002),
.C(n_900),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_999),
.B(n_1002),
.Y(n_1176)
);

NOR2x1_ASAP7_75t_L g1177 ( 
.A(n_896),
.B(n_761),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1054),
.A2(n_1056),
.B(n_897),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_999),
.B(n_1002),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_932),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1051),
.A2(n_816),
.B1(n_807),
.B2(n_1044),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1054),
.A2(n_831),
.B(n_816),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1054),
.A2(n_831),
.B(n_816),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_999),
.B(n_1002),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1051),
.A2(n_816),
.B1(n_807),
.B2(n_1044),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_993),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1054),
.A2(n_831),
.B(n_1056),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_944),
.B(n_811),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_999),
.A2(n_1002),
.B1(n_1051),
.B2(n_886),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1054),
.A2(n_1056),
.A3(n_1023),
.B(n_846),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_999),
.A2(n_1002),
.B(n_1051),
.C(n_1047),
.Y(n_1191)
);

AO21x1_ASAP7_75t_L g1192 ( 
.A1(n_999),
.A2(n_1002),
.B(n_996),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1069),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1143),
.B(n_1144),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1104),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1059),
.B(n_1142),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1138),
.B(n_1093),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1112),
.A2(n_1099),
.B(n_1061),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1081),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1099),
.A2(n_1163),
.B(n_1153),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1074),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1182),
.A2(n_1183),
.B(n_1100),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1075),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1107),
.Y(n_1204)
);

OAI21xp33_ASAP7_75t_L g1205 ( 
.A1(n_1174),
.A2(n_1189),
.B(n_1073),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1142),
.B(n_1154),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1157),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1154),
.B(n_1156),
.Y(n_1208)
);

OR2x6_ASAP7_75t_L g1209 ( 
.A(n_1066),
.B(n_1079),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1152),
.B(n_1155),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1113),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1180),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_1164),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1106),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1156),
.B(n_1158),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1124),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1158),
.B(n_1169),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_1138),
.B(n_1093),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1169),
.B(n_1172),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1060),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1172),
.B(n_1176),
.Y(n_1221)
);

BUFx4_ASAP7_75t_SL g1222 ( 
.A(n_1098),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1176),
.A2(n_1179),
.B1(n_1184),
.B2(n_1058),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1091),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1164),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1188),
.B(n_1063),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1179),
.B(n_1184),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1121),
.B(n_1160),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1130),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1164),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1111),
.A2(n_1159),
.B(n_1191),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1168),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_L g1233 ( 
.A(n_1167),
.B(n_1095),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1148),
.B(n_1065),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1168),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1138),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1065),
.B(n_1146),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1130),
.B(n_1066),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1149),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1125),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1146),
.B(n_1175),
.Y(n_1241)
);

OAI21xp33_ASAP7_75t_L g1242 ( 
.A1(n_1085),
.A2(n_1133),
.B(n_1119),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1066),
.B(n_1135),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1126),
.B(n_1122),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1125),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1082),
.A2(n_1111),
.B(n_1102),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1168),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1072),
.B(n_1108),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1181),
.A2(n_1185),
.B1(n_1119),
.B2(n_1067),
.Y(n_1249)
);

AND2x2_ASAP7_75t_SL g1250 ( 
.A(n_1128),
.B(n_1114),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1170),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1165),
.Y(n_1252)
);

OR2x6_ASAP7_75t_L g1253 ( 
.A(n_1115),
.B(n_1125),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1108),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1170),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1090),
.B(n_1077),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1137),
.Y(n_1257)
);

NOR2x1_ASAP7_75t_SL g1258 ( 
.A(n_1084),
.B(n_1086),
.Y(n_1258)
);

BUFx10_ASAP7_75t_L g1259 ( 
.A(n_1170),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1145),
.B(n_1173),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1173),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1173),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_1084),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_1186),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1117),
.B(n_1083),
.Y(n_1265)
);

AO21x2_ASAP7_75t_L g1266 ( 
.A1(n_1147),
.A2(n_1171),
.B(n_1178),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_L g1267 ( 
.A(n_1145),
.B(n_1068),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1070),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_1089),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1137),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1181),
.A2(n_1185),
.B1(n_1109),
.B2(n_1083),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1187),
.A2(n_1078),
.B(n_1120),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1186),
.B(n_1177),
.Y(n_1273)
);

INVx3_ASAP7_75t_SL g1274 ( 
.A(n_1134),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1116),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1057),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1186),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1064),
.B(n_1133),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1166),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1064),
.B(n_1062),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1062),
.B(n_1071),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1192),
.B(n_1139),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1105),
.B(n_1092),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1086),
.A2(n_1178),
.B1(n_1150),
.B2(n_1140),
.Y(n_1284)
);

BUFx12f_ASAP7_75t_L g1285 ( 
.A(n_1116),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1115),
.Y(n_1286)
);

BUFx10_ASAP7_75t_L g1287 ( 
.A(n_1161),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1161),
.A2(n_1131),
.B1(n_1151),
.B2(n_1140),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1110),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1161),
.Y(n_1290)
);

OR2x2_ASAP7_75t_SL g1291 ( 
.A(n_1136),
.B(n_1161),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1080),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1118),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1088),
.B(n_1094),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1123),
.A2(n_1132),
.B(n_1141),
.C(n_1097),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1127),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1131),
.A2(n_1129),
.B1(n_1190),
.B2(n_1087),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1129),
.B(n_1096),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1129),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1190),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1103),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1076),
.A2(n_751),
.B(n_1002),
.C(n_999),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1101),
.B(n_1093),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1189),
.A2(n_1174),
.B1(n_816),
.B2(n_1142),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1074),
.Y(n_1305)
);

NAND2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1138),
.B(n_1093),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1069),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1074),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1138),
.Y(n_1309)
);

AOI222xp33_ASAP7_75t_L g1310 ( 
.A1(n_1071),
.A2(n_1013),
.B1(n_1047),
.B2(n_1044),
.C1(n_976),
.C2(n_751),
.Y(n_1310)
);

NAND2xp33_ASAP7_75t_SL g1311 ( 
.A(n_1164),
.B(n_1168),
.Y(n_1311)
);

OR2x4_ASAP7_75t_L g1312 ( 
.A(n_1095),
.B(n_753),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1189),
.A2(n_1174),
.B1(n_816),
.B2(n_1142),
.Y(n_1313)
);

INVxp67_ASAP7_75t_SL g1314 ( 
.A(n_1162),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1112),
.A2(n_1099),
.B(n_831),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1059),
.B(n_1142),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1059),
.B(n_1142),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1189),
.A2(n_1174),
.B1(n_816),
.B2(n_1142),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1112),
.A2(n_1099),
.B(n_831),
.Y(n_1319)
);

OAI21xp33_ASAP7_75t_L g1320 ( 
.A1(n_1174),
.A2(n_767),
.B(n_753),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1074),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1059),
.B(n_1142),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1069),
.Y(n_1323)
);

O2A1O1Ixp5_ASAP7_75t_SL g1324 ( 
.A1(n_1140),
.A2(n_900),
.B(n_751),
.C(n_1146),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1174),
.A2(n_753),
.B1(n_927),
.B2(n_918),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1112),
.A2(n_1099),
.B(n_831),
.Y(n_1326)
);

OR2x6_ASAP7_75t_L g1327 ( 
.A(n_1066),
.B(n_1079),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1174),
.A2(n_1002),
.B(n_999),
.Y(n_1328)
);

AND2x6_ASAP7_75t_L g1329 ( 
.A(n_1138),
.B(n_976),
.Y(n_1329)
);

CKINVDCx6p67_ASAP7_75t_R g1330 ( 
.A(n_1079),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1174),
.B(n_753),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1143),
.B(n_1144),
.Y(n_1332)
);

AOI221x1_ASAP7_75t_L g1333 ( 
.A1(n_1073),
.A2(n_1099),
.B1(n_1111),
.B2(n_1112),
.C(n_1191),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1112),
.A2(n_1099),
.B(n_831),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1104),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1143),
.B(n_1144),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1138),
.Y(n_1337)
);

NOR2x1_ASAP7_75t_SL g1338 ( 
.A(n_1066),
.B(n_1084),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1174),
.B(n_634),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1104),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1203),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1212),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1320),
.A2(n_1331),
.B1(n_1242),
.B2(n_1205),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1216),
.Y(n_1344)
);

BUFx2_ASAP7_75t_SL g1345 ( 
.A(n_1195),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1250),
.A2(n_1278),
.B1(n_1256),
.B2(n_1231),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1325),
.A2(n_1318),
.B1(n_1313),
.B2(n_1304),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1220),
.Y(n_1348)
);

OR2x6_ASAP7_75t_L g1349 ( 
.A(n_1253),
.B(n_1290),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1305),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1310),
.A2(n_1328),
.B1(n_1231),
.B2(n_1281),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1194),
.B(n_1210),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1225),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1310),
.A2(n_1328),
.B1(n_1313),
.B2(n_1304),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1321),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1318),
.A2(n_1339),
.B1(n_1249),
.B2(n_1280),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1243),
.B(n_1286),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1335),
.Y(n_1358)
);

AO21x1_ASAP7_75t_L g1359 ( 
.A1(n_1223),
.A2(n_1249),
.B(n_1282),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1299),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1201),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1204),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1207),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1269),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1283),
.Y(n_1365)
);

INVx6_ASAP7_75t_L g1366 ( 
.A(n_1259),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1225),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1244),
.A2(n_1329),
.B1(n_1228),
.B2(n_1208),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1227),
.A2(n_1312),
.B1(n_1316),
.B2(n_1196),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_SL g1370 ( 
.A(n_1209),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1223),
.A2(n_1266),
.B1(n_1246),
.B2(n_1241),
.Y(n_1371)
);

NAND2x1p5_ASAP7_75t_L g1372 ( 
.A(n_1286),
.B(n_1243),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1308),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1312),
.A2(n_1219),
.B1(n_1217),
.B2(n_1196),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1266),
.A2(n_1246),
.B1(n_1241),
.B2(n_1219),
.Y(n_1375)
);

CKINVDCx11_ASAP7_75t_R g1376 ( 
.A(n_1276),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1299),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1199),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1298),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1283),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1198),
.A2(n_1200),
.B(n_1272),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1229),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1239),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1215),
.B(n_1332),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1252),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1268),
.Y(n_1386)
);

AO21x2_ASAP7_75t_L g1387 ( 
.A1(n_1295),
.A2(n_1334),
.B(n_1315),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1336),
.B(n_1226),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1225),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1302),
.A2(n_1333),
.B(n_1324),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1329),
.A2(n_1193),
.B1(n_1323),
.B2(n_1307),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1298),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1329),
.A2(n_1307),
.B1(n_1323),
.B2(n_1338),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1259),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1206),
.A2(n_1221),
.B1(n_1317),
.B2(n_1322),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1214),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1222),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1211),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1254),
.A2(n_1248),
.B1(n_1265),
.B2(n_1233),
.Y(n_1399)
);

OR2x6_ASAP7_75t_L g1400 ( 
.A(n_1253),
.B(n_1209),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1302),
.A2(n_1319),
.B(n_1326),
.Y(n_1401)
);

AO21x2_ASAP7_75t_L g1402 ( 
.A1(n_1326),
.A2(n_1334),
.B(n_1202),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1253),
.B(n_1238),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1237),
.A2(n_1271),
.B1(n_1263),
.B2(n_1234),
.Y(n_1404)
);

NOR2x1_ASAP7_75t_R g1405 ( 
.A(n_1340),
.B(n_1285),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1329),
.A2(n_1245),
.B1(n_1240),
.B2(n_1270),
.Y(n_1406)
);

OR2x6_ASAP7_75t_L g1407 ( 
.A(n_1209),
.B(n_1327),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1257),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1197),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1293),
.Y(n_1410)
);

INVx6_ASAP7_75t_L g1411 ( 
.A(n_1264),
.Y(n_1411)
);

INVx5_ASAP7_75t_L g1412 ( 
.A(n_1327),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1293),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1293),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1258),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1294),
.A2(n_1297),
.B(n_1284),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1301),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1314),
.B(n_1291),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1287),
.A2(n_1284),
.B1(n_1238),
.B2(n_1273),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1300),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1273),
.B(n_1327),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1247),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1303),
.B(n_1337),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1292),
.A2(n_1288),
.B(n_1296),
.Y(n_1424)
);

BUFx4f_ASAP7_75t_SL g1425 ( 
.A(n_1274),
.Y(n_1425)
);

BUFx2_ASAP7_75t_SL g1426 ( 
.A(n_1224),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1296),
.A2(n_1287),
.B(n_1267),
.Y(n_1427)
);

INVx5_ASAP7_75t_L g1428 ( 
.A(n_1247),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1275),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1197),
.A2(n_1306),
.B(n_1218),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1306),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1236),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1279),
.A2(n_1289),
.B1(n_1261),
.B2(n_1255),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1236),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1309),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1230),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1232),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1337),
.A2(n_1330),
.B1(n_1260),
.B2(n_1251),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1247),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1262),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1262),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1262),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1277),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1277),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1260),
.B(n_1213),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1213),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1277),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1311),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1235),
.Y(n_1449)
);

INVx5_ASAP7_75t_L g1450 ( 
.A(n_1253),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1203),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1203),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_SL g1453 ( 
.A1(n_1331),
.A2(n_1013),
.B1(n_1047),
.B2(n_753),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1195),
.Y(n_1454)
);

INVx4_ASAP7_75t_SL g1455 ( 
.A(n_1329),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1331),
.A2(n_1013),
.B1(n_1047),
.B2(n_753),
.Y(n_1456)
);

INVx6_ASAP7_75t_L g1457 ( 
.A(n_1259),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1194),
.B(n_1210),
.Y(n_1458)
);

INVxp33_ASAP7_75t_L g1459 ( 
.A(n_1194),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1283),
.Y(n_1460)
);

AO21x1_ASAP7_75t_L g1461 ( 
.A1(n_1331),
.A2(n_1325),
.B(n_1278),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1203),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1320),
.A2(n_1331),
.B1(n_1242),
.B2(n_1051),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1208),
.B(n_1227),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1225),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1194),
.B(n_1210),
.Y(n_1466)
);

BUFx4f_ASAP7_75t_SL g1467 ( 
.A(n_1195),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1203),
.Y(n_1468)
);

CKINVDCx11_ASAP7_75t_R g1469 ( 
.A(n_1269),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1320),
.A2(n_1331),
.B1(n_1242),
.B2(n_1051),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1225),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1320),
.A2(n_1331),
.B1(n_1242),
.B2(n_1051),
.Y(n_1472)
);

OR2x6_ASAP7_75t_L g1473 ( 
.A(n_1253),
.B(n_1290),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1225),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1203),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1320),
.A2(n_1331),
.B1(n_1242),
.B2(n_1051),
.Y(n_1476)
);

CKINVDCx11_ASAP7_75t_R g1477 ( 
.A(n_1269),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1283),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1194),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1203),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1208),
.B(n_1227),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1194),
.B(n_1210),
.Y(n_1482)
);

CKINVDCx11_ASAP7_75t_R g1483 ( 
.A(n_1269),
.Y(n_1483)
);

BUFx2_ASAP7_75t_SL g1484 ( 
.A(n_1195),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1203),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1285),
.Y(n_1486)
);

BUFx10_ASAP7_75t_L g1487 ( 
.A(n_1211),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1454),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1464),
.B(n_1481),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1423),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1360),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1379),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1360),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1377),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1455),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1377),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1390),
.A2(n_1401),
.B(n_1381),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1351),
.B(n_1375),
.Y(n_1498)
);

AO21x1_ASAP7_75t_SL g1499 ( 
.A1(n_1354),
.A2(n_1351),
.B(n_1356),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1379),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1352),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1369),
.B(n_1384),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1375),
.B(n_1346),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1356),
.B(n_1392),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1453),
.B(n_1456),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1392),
.B(n_1371),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1354),
.A2(n_1371),
.B(n_1359),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1395),
.B(n_1374),
.Y(n_1508)
);

BUFx4f_ASAP7_75t_SL g1509 ( 
.A(n_1454),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1417),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1400),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1397),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1417),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1461),
.A2(n_1343),
.B1(n_1347),
.B2(n_1476),
.Y(n_1514)
);

INVx4_ASAP7_75t_L g1515 ( 
.A(n_1455),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1424),
.Y(n_1516)
);

NAND2x1p5_ASAP7_75t_L g1517 ( 
.A(n_1450),
.B(n_1424),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1420),
.Y(n_1518)
);

NAND2x1_ASAP7_75t_L g1519 ( 
.A(n_1415),
.B(n_1427),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1402),
.Y(n_1520)
);

BUFx2_ASAP7_75t_R g1521 ( 
.A(n_1397),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1404),
.B(n_1343),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1396),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1463),
.B(n_1470),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1400),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1387),
.A2(n_1413),
.B(n_1410),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1387),
.A2(n_1413),
.B(n_1410),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1416),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1424),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1463),
.B(n_1470),
.Y(n_1530)
);

AO21x2_ASAP7_75t_L g1531 ( 
.A1(n_1414),
.A2(n_1362),
.B(n_1361),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1349),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1472),
.B(n_1476),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1416),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1427),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1399),
.B(n_1472),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1408),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_SL g1538 ( 
.A(n_1467),
.B(n_1398),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1485),
.B(n_1459),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1363),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1373),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1349),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1341),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1342),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1429),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1344),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1350),
.Y(n_1547)
);

NAND2x1p5_ASAP7_75t_L g1548 ( 
.A(n_1427),
.B(n_1412),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1430),
.A2(n_1372),
.B(n_1468),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1400),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1355),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1451),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1452),
.Y(n_1553)
);

AO21x2_ASAP7_75t_L g1554 ( 
.A1(n_1448),
.A2(n_1480),
.B(n_1475),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1412),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1462),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1383),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1385),
.Y(n_1558)
);

INVx4_ASAP7_75t_L g1559 ( 
.A(n_1412),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1459),
.B(n_1388),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1386),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1479),
.B(n_1418),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1349),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1473),
.B(n_1368),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1458),
.B(n_1466),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1482),
.B(n_1357),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1412),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1357),
.B(n_1403),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1357),
.B(n_1403),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1432),
.A2(n_1435),
.B(n_1434),
.Y(n_1570)
);

NOR2x1_ASAP7_75t_L g1571 ( 
.A(n_1473),
.B(n_1407),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1370),
.A2(n_1407),
.B1(n_1358),
.B2(n_1403),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1372),
.Y(n_1573)
);

INVx5_ASAP7_75t_SL g1574 ( 
.A(n_1407),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1473),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1378),
.Y(n_1576)
);

AO21x2_ASAP7_75t_L g1577 ( 
.A1(n_1439),
.A2(n_1440),
.B(n_1447),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1419),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1382),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1393),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1409),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1391),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1444),
.A2(n_1443),
.B(n_1442),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1406),
.Y(n_1584)
);

OA21x2_ASAP7_75t_L g1585 ( 
.A1(n_1449),
.A2(n_1421),
.B(n_1438),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1431),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1365),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1365),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1380),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1460),
.A2(n_1478),
.B(n_1446),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1460),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1449),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1478),
.Y(n_1593)
);

AOI21x1_ASAP7_75t_L g1594 ( 
.A1(n_1445),
.A2(n_1433),
.B(n_1370),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1428),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1428),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1428),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1506),
.B(n_1367),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1506),
.B(n_1367),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1535),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1504),
.B(n_1510),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1491),
.B(n_1426),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_SL g1603 ( 
.A(n_1521),
.B(n_1425),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1504),
.B(n_1367),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1531),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1565),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1522),
.A2(n_1503),
.B1(n_1498),
.B2(n_1524),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1491),
.B(n_1345),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1488),
.Y(n_1609)
);

AO21x2_ASAP7_75t_L g1610 ( 
.A1(n_1520),
.A2(n_1474),
.B(n_1353),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1583),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1513),
.B(n_1540),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1563),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1540),
.B(n_1465),
.Y(n_1614)
);

OAI21xp33_ASAP7_75t_L g1615 ( 
.A1(n_1505),
.A2(n_1348),
.B(n_1437),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1563),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1493),
.B(n_1484),
.Y(n_1617)
);

NOR2x1p5_ASAP7_75t_L g1618 ( 
.A(n_1511),
.B(n_1525),
.Y(n_1618)
);

INVxp67_ASAP7_75t_R g1619 ( 
.A(n_1590),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1492),
.Y(n_1620)
);

BUFx4f_ASAP7_75t_SL g1621 ( 
.A(n_1576),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1539),
.B(n_1541),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1523),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1500),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1523),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1579),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1509),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1554),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1502),
.B(n_1353),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1503),
.B(n_1422),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1518),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1554),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1563),
.B(n_1445),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1554),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1493),
.B(n_1494),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1489),
.B(n_1422),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1560),
.B(n_1389),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1499),
.A2(n_1376),
.B1(n_1477),
.B2(n_1364),
.Y(n_1638)
);

NOR2x1_ASAP7_75t_L g1639 ( 
.A(n_1570),
.B(n_1446),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1511),
.B(n_1525),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1519),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1579),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1560),
.B(n_1471),
.Y(n_1643)
);

AND2x4_ASAP7_75t_SL g1644 ( 
.A(n_1495),
.B(n_1487),
.Y(n_1644)
);

NOR2x1_ASAP7_75t_L g1645 ( 
.A(n_1577),
.B(n_1398),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1494),
.B(n_1437),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1583),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1583),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1511),
.B(n_1422),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1501),
.B(n_1467),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1498),
.B(n_1474),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1517),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1514),
.A2(n_1425),
.B1(n_1486),
.B2(n_1457),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1496),
.B(n_1436),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1517),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1524),
.B(n_1389),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1592),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1522),
.B(n_1537),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1530),
.B(n_1474),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1538),
.B(n_1364),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1530),
.B(n_1436),
.Y(n_1661)
);

AOI211xp5_ASAP7_75t_L g1662 ( 
.A1(n_1508),
.A2(n_1405),
.B(n_1376),
.C(n_1483),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1533),
.B(n_1441),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1533),
.B(n_1441),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1496),
.B(n_1487),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1601),
.B(n_1613),
.Y(n_1666)
);

NOR3xp33_ASAP7_75t_L g1667 ( 
.A(n_1653),
.B(n_1594),
.C(n_1571),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1615),
.A2(n_1499),
.B1(n_1578),
.B2(n_1550),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1657),
.B(n_1658),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1616),
.B(n_1529),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1645),
.A2(n_1571),
.B(n_1594),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1616),
.B(n_1529),
.Y(n_1672)
);

AOI211xp5_ASAP7_75t_SL g1673 ( 
.A1(n_1662),
.A2(n_1580),
.B(n_1564),
.C(n_1578),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1622),
.B(n_1562),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1598),
.B(n_1599),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1622),
.B(n_1545),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1638),
.A2(n_1572),
.B(n_1549),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1599),
.B(n_1516),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1642),
.B(n_1536),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1607),
.B(n_1490),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1606),
.A2(n_1584),
.B1(n_1582),
.B2(n_1580),
.C(n_1566),
.Y(n_1681)
);

NOR3xp33_ASAP7_75t_L g1682 ( 
.A(n_1650),
.B(n_1584),
.C(n_1582),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1604),
.B(n_1516),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1604),
.B(n_1516),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1626),
.B(n_1536),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1663),
.A2(n_1550),
.B1(n_1564),
.B2(n_1532),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1637),
.B(n_1497),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1608),
.B(n_1547),
.Y(n_1688)
);

NOR3xp33_ASAP7_75t_L g1689 ( 
.A(n_1629),
.B(n_1542),
.C(n_1532),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1608),
.B(n_1547),
.Y(n_1690)
);

NOR3xp33_ASAP7_75t_L g1691 ( 
.A(n_1660),
.B(n_1542),
.C(n_1559),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_SL g1692 ( 
.A1(n_1644),
.A2(n_1568),
.B(n_1569),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1617),
.B(n_1507),
.C(n_1585),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1617),
.B(n_1507),
.C(n_1585),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1663),
.A2(n_1550),
.B1(n_1507),
.B2(n_1574),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1643),
.B(n_1497),
.Y(n_1696)
);

NAND4xp25_ASAP7_75t_L g1697 ( 
.A(n_1636),
.B(n_1551),
.C(n_1553),
.D(n_1556),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1631),
.B(n_1551),
.Y(n_1698)
);

OAI21xp33_ASAP7_75t_L g1699 ( 
.A1(n_1603),
.A2(n_1566),
.B(n_1553),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_SL g1700 ( 
.A(n_1609),
.B(n_1548),
.C(n_1512),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1618),
.A2(n_1507),
.B(n_1495),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1623),
.Y(n_1702)
);

OA21x2_ASAP7_75t_L g1703 ( 
.A1(n_1628),
.A2(n_1528),
.B(n_1534),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1612),
.B(n_1517),
.Y(n_1704)
);

NAND3xp33_ASAP7_75t_L g1705 ( 
.A(n_1639),
.B(n_1585),
.C(n_1520),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1612),
.B(n_1526),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_SL g1707 ( 
.A1(n_1664),
.A2(n_1574),
.B1(n_1575),
.B2(n_1495),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1623),
.Y(n_1708)
);

AND2x2_ASAP7_75t_SL g1709 ( 
.A(n_1652),
.B(n_1495),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1639),
.A2(n_1549),
.B(n_1590),
.Y(n_1710)
);

OAI21xp33_ASAP7_75t_L g1711 ( 
.A1(n_1664),
.A2(n_1556),
.B(n_1557),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1621),
.A2(n_1574),
.B1(n_1515),
.B2(n_1575),
.Y(n_1712)
);

OAI221xp5_ASAP7_75t_SL g1713 ( 
.A1(n_1665),
.A2(n_1575),
.B1(n_1588),
.B2(n_1591),
.C(n_1589),
.Y(n_1713)
);

NOR3xp33_ASAP7_75t_L g1714 ( 
.A(n_1665),
.B(n_1559),
.C(n_1515),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1640),
.B(n_1490),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1661),
.B(n_1543),
.Y(n_1716)
);

NAND3xp33_ASAP7_75t_L g1717 ( 
.A(n_1632),
.B(n_1585),
.C(n_1573),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1656),
.B(n_1526),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1656),
.B(n_1543),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1659),
.B(n_1544),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1659),
.B(n_1544),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1651),
.B(n_1526),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1618),
.A2(n_1515),
.B(n_1548),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1609),
.A2(n_1574),
.B1(n_1515),
.B2(n_1602),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_L g1725 ( 
.A(n_1632),
.B(n_1573),
.C(n_1593),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1627),
.B(n_1568),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1651),
.A2(n_1561),
.B1(n_1557),
.B2(n_1558),
.C(n_1552),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1630),
.B(n_1527),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1614),
.B(n_1546),
.Y(n_1729)
);

OAI211xp5_ASAP7_75t_L g1730 ( 
.A1(n_1630),
.A2(n_1652),
.B(n_1655),
.C(n_1654),
.Y(n_1730)
);

OAI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1655),
.A2(n_1548),
.B1(n_1581),
.B2(n_1567),
.C(n_1555),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1625),
.B(n_1527),
.Y(n_1732)
);

NAND3xp33_ASAP7_75t_L g1733 ( 
.A(n_1634),
.B(n_1587),
.C(n_1593),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1646),
.A2(n_1586),
.B(n_1567),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_L g1735 ( 
.A(n_1646),
.B(n_1654),
.C(n_1561),
.D(n_1558),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1675),
.B(n_1619),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1675),
.B(n_1619),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1669),
.B(n_1620),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1702),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1670),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1703),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1687),
.B(n_1600),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1687),
.B(n_1600),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1702),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1706),
.B(n_1624),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1708),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1708),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1732),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1703),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1714),
.B(n_1641),
.Y(n_1750)
);

NOR2xp67_ASAP7_75t_L g1751 ( 
.A(n_1693),
.B(n_1611),
.Y(n_1751)
);

BUFx2_ASAP7_75t_L g1752 ( 
.A(n_1709),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1706),
.B(n_1605),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1732),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1696),
.B(n_1666),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1698),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1672),
.B(n_1635),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1704),
.B(n_1641),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1704),
.B(n_1641),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1726),
.B(n_1469),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1676),
.B(n_1647),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1688),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1690),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1678),
.B(n_1683),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1684),
.B(n_1648),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1718),
.B(n_1605),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1722),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1709),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1733),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1728),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1728),
.B(n_1610),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1729),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1719),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1680),
.A2(n_1633),
.B1(n_1640),
.B2(n_1490),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1722),
.B(n_1610),
.Y(n_1775)
);

INVxp67_ASAP7_75t_L g1776 ( 
.A(n_1674),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1694),
.B(n_1648),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1720),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1689),
.B(n_1610),
.Y(n_1779)
);

INVxp67_ASAP7_75t_SL g1780 ( 
.A(n_1751),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1762),
.B(n_1711),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1752),
.B(n_1768),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1739),
.Y(n_1783)
);

AND2x2_ASAP7_75t_SL g1784 ( 
.A(n_1752),
.B(n_1667),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1768),
.B(n_1691),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1760),
.B(n_1469),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1765),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1758),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1762),
.B(n_1711),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1769),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1736),
.B(n_1715),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1741),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1739),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1763),
.B(n_1721),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1769),
.B(n_1716),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1736),
.B(n_1671),
.Y(n_1796)
);

AOI33xp33_ASAP7_75t_L g1797 ( 
.A1(n_1779),
.A2(n_1681),
.A3(n_1695),
.B1(n_1686),
.B2(n_1668),
.B3(n_1727),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1737),
.B(n_1730),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1744),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1737),
.B(n_1758),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1750),
.B(n_1710),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1744),
.Y(n_1802)
);

OR2x6_ASAP7_75t_L g1803 ( 
.A(n_1751),
.B(n_1701),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1758),
.B(n_1723),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1758),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1759),
.B(n_1723),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1741),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1746),
.Y(n_1808)
);

NAND3xp33_ASAP7_75t_L g1809 ( 
.A(n_1779),
.B(n_1682),
.C(n_1673),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1746),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1741),
.Y(n_1811)
);

OAI21xp33_ASAP7_75t_L g1812 ( 
.A1(n_1774),
.A2(n_1699),
.B(n_1735),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1747),
.Y(n_1813)
);

AND2x4_ASAP7_75t_SL g1814 ( 
.A(n_1750),
.B(n_1649),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1763),
.B(n_1685),
.Y(n_1815)
);

AND2x4_ASAP7_75t_SL g1816 ( 
.A(n_1750),
.B(n_1649),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1756),
.B(n_1679),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1747),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1777),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1750),
.B(n_1717),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1759),
.B(n_1701),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1748),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1754),
.Y(n_1823)
);

OR2x6_ASAP7_75t_L g1824 ( 
.A(n_1777),
.B(n_1677),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1759),
.B(n_1734),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1756),
.B(n_1697),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1759),
.B(n_1707),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1766),
.B(n_1705),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1766),
.B(n_1725),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1749),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1753),
.B(n_1634),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1828),
.B(n_1745),
.Y(n_1832)
);

INVxp67_ASAP7_75t_SL g1833 ( 
.A(n_1780),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1826),
.B(n_1772),
.Y(n_1834)
);

NOR3xp33_ASAP7_75t_L g1835 ( 
.A(n_1809),
.B(n_1812),
.C(n_1790),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1782),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1804),
.B(n_1777),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1804),
.B(n_1771),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1783),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1783),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1806),
.B(n_1771),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1806),
.B(n_1775),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1828),
.B(n_1745),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1829),
.B(n_1753),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1792),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1793),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1821),
.B(n_1775),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1793),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1821),
.B(n_1767),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1800),
.B(n_1767),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1781),
.B(n_1772),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1789),
.B(n_1773),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1792),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1795),
.B(n_1773),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1807),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1799),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1829),
.B(n_1767),
.Y(n_1857)
);

AND2x2_ASAP7_75t_SL g1858 ( 
.A(n_1784),
.B(n_1777),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1799),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1802),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1795),
.B(n_1778),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1803),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1800),
.B(n_1770),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1782),
.B(n_1755),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1831),
.B(n_1761),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1827),
.B(n_1755),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1802),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1831),
.B(n_1761),
.Y(n_1868)
);

NOR3xp33_ASAP7_75t_L g1869 ( 
.A(n_1797),
.B(n_1700),
.C(n_1731),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1785),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1785),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1815),
.B(n_1778),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1817),
.B(n_1776),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1808),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1784),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1808),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1807),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1827),
.B(n_1764),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1810),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_SL g1880 ( 
.A(n_1784),
.B(n_1699),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1805),
.B(n_1764),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1805),
.B(n_1742),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1814),
.B(n_1742),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1819),
.B(n_1757),
.Y(n_1884)
);

AOI211xp5_ASAP7_75t_L g1885 ( 
.A1(n_1820),
.A2(n_1724),
.B(n_1712),
.C(n_1692),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1814),
.B(n_1743),
.Y(n_1886)
);

NAND2xp67_ASAP7_75t_L g1887 ( 
.A(n_1816),
.B(n_1477),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1881),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1839),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1839),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1858),
.B(n_1816),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1835),
.B(n_1798),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1884),
.B(n_1824),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1881),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1884),
.B(n_1832),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1869),
.A2(n_1824),
.B1(n_1798),
.B2(n_1803),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1832),
.B(n_1843),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1875),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1840),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1858),
.B(n_1796),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1836),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1845),
.Y(n_1902)
);

NAND3xp33_ASAP7_75t_L g1903 ( 
.A(n_1880),
.B(n_1824),
.C(n_1803),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1845),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1840),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1856),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1878),
.A2(n_1824),
.B1(n_1803),
.B2(n_1796),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1870),
.A2(n_1820),
.B1(n_1713),
.B2(n_1740),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1843),
.B(n_1822),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1878),
.B(n_1788),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1856),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1859),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1864),
.B(n_1866),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1859),
.Y(n_1914)
);

AOI22x1_ASAP7_75t_L g1915 ( 
.A1(n_1833),
.A2(n_1820),
.B1(n_1801),
.B2(n_1788),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1864),
.B(n_1801),
.Y(n_1916)
);

NAND2x1p5_ASAP7_75t_L g1917 ( 
.A(n_1862),
.B(n_1820),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1866),
.B(n_1801),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1862),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1853),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1871),
.B(n_1791),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1853),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1855),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1883),
.B(n_1801),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1855),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1834),
.B(n_1791),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1873),
.B(n_1794),
.Y(n_1927)
);

BUFx3_ASAP7_75t_L g1928 ( 
.A(n_1860),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1844),
.B(n_1822),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1896),
.B(n_1885),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1898),
.B(n_1851),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1903),
.B(n_1837),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1928),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1928),
.Y(n_1934)
);

AOI211x1_ASAP7_75t_L g1935 ( 
.A1(n_1892),
.A2(n_1852),
.B(n_1861),
.C(n_1854),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_SL g1936 ( 
.A(n_1903),
.B(n_1786),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1908),
.A2(n_1896),
.B(n_1900),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1908),
.A2(n_1872),
.B(n_1837),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1928),
.Y(n_1939)
);

INVx2_ASAP7_75t_SL g1940 ( 
.A(n_1891),
.Y(n_1940)
);

OAI211xp5_ASAP7_75t_L g1941 ( 
.A1(n_1915),
.A2(n_1844),
.B(n_1838),
.C(n_1842),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1889),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1895),
.B(n_1897),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1917),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1900),
.A2(n_1837),
.B(n_1846),
.Y(n_1945)
);

INVxp67_ASAP7_75t_L g1946 ( 
.A(n_1919),
.Y(n_1946)
);

AOI21xp33_ASAP7_75t_L g1947 ( 
.A1(n_1915),
.A2(n_1857),
.B(n_1860),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1895),
.B(n_1857),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1901),
.B(n_1863),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1889),
.Y(n_1950)
);

AOI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1891),
.A2(n_1883),
.B1(n_1886),
.B2(n_1863),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1901),
.A2(n_1886),
.B1(n_1841),
.B2(n_1842),
.Y(n_1952)
);

A2O1A1Ixp33_ASAP7_75t_L g1953 ( 
.A1(n_1907),
.A2(n_1919),
.B(n_1893),
.C(n_1897),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1890),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1893),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1913),
.B(n_1838),
.Y(n_1956)
);

AOI22xp33_ASAP7_75t_L g1957 ( 
.A1(n_1921),
.A2(n_1841),
.B1(n_1847),
.B2(n_1849),
.Y(n_1957)
);

OAI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1917),
.A2(n_1847),
.B1(n_1825),
.B2(n_1787),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1890),
.Y(n_1959)
);

AOI211xp5_ASAP7_75t_L g1960 ( 
.A1(n_1918),
.A2(n_1849),
.B(n_1867),
.C(n_1874),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1936),
.Y(n_1961)
);

INVxp33_ASAP7_75t_L g1962 ( 
.A(n_1932),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1943),
.B(n_1917),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1934),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1949),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1934),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1940),
.B(n_1913),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1946),
.B(n_1888),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1946),
.B(n_1888),
.Y(n_1969)
);

NAND2x1_ASAP7_75t_L g1970 ( 
.A(n_1944),
.B(n_1888),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1951),
.B(n_1894),
.Y(n_1971)
);

OAI21xp33_ASAP7_75t_L g1972 ( 
.A1(n_1930),
.A2(n_1926),
.B(n_1918),
.Y(n_1972)
);

OR2x2_ASAP7_75t_L g1973 ( 
.A(n_1948),
.B(n_1894),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1955),
.B(n_1894),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1935),
.B(n_1927),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1952),
.B(n_1910),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1942),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1953),
.B(n_1910),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1957),
.B(n_1924),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1933),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1950),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1957),
.B(n_1924),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1954),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1956),
.B(n_1916),
.Y(n_1984)
);

OAI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1961),
.A2(n_1930),
.B(n_1937),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1967),
.B(n_1939),
.Y(n_1986)
);

OAI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1962),
.A2(n_1938),
.B(n_1941),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1967),
.B(n_1916),
.Y(n_1988)
);

NOR3x1_ASAP7_75t_L g1989 ( 
.A(n_1978),
.B(n_1931),
.C(n_1958),
.Y(n_1989)
);

AOI222xp33_ASAP7_75t_L g1990 ( 
.A1(n_1975),
.A2(n_1959),
.B1(n_1905),
.B2(n_1899),
.C1(n_1914),
.C2(n_1906),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1963),
.A2(n_1947),
.B(n_1945),
.Y(n_1991)
);

A2O1A1Ixp33_ASAP7_75t_L g1992 ( 
.A1(n_1972),
.A2(n_1960),
.B(n_1909),
.C(n_1899),
.Y(n_1992)
);

OAI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1965),
.A2(n_1909),
.B1(n_1787),
.B2(n_1929),
.Y(n_1993)
);

NOR3x1_ASAP7_75t_L g1994 ( 
.A(n_1968),
.B(n_1906),
.C(n_1905),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1974),
.A2(n_1912),
.B(n_1911),
.Y(n_1995)
);

OAI211xp5_ASAP7_75t_SL g1996 ( 
.A1(n_1969),
.A2(n_1483),
.B(n_1912),
.C(n_1911),
.Y(n_1996)
);

NOR3xp33_ASAP7_75t_L g1997 ( 
.A(n_1980),
.B(n_1914),
.C(n_1904),
.Y(n_1997)
);

OAI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1979),
.A2(n_1929),
.B(n_1904),
.Y(n_1998)
);

AOI211xp5_ASAP7_75t_SL g1999 ( 
.A1(n_1964),
.A2(n_1904),
.B(n_1920),
.C(n_1902),
.Y(n_1999)
);

NAND4xp25_ASAP7_75t_L g2000 ( 
.A(n_1985),
.B(n_1979),
.C(n_1982),
.D(n_1971),
.Y(n_2000)
);

NAND4xp75_ASAP7_75t_L g2001 ( 
.A(n_1989),
.B(n_1966),
.C(n_1964),
.D(n_1971),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1986),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1988),
.B(n_1976),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1991),
.B(n_1976),
.Y(n_2004)
);

AND5x1_ASAP7_75t_L g2005 ( 
.A(n_1992),
.B(n_1982),
.C(n_1970),
.D(n_1973),
.E(n_1984),
.Y(n_2005)
);

NAND4xp75_ASAP7_75t_L g2006 ( 
.A(n_1994),
.B(n_1966),
.C(n_1980),
.D(n_1977),
.Y(n_2006)
);

NOR2x1_ASAP7_75t_L g2007 ( 
.A(n_1987),
.B(n_1970),
.Y(n_2007)
);

AOI21xp5_ASAP7_75t_SL g2008 ( 
.A1(n_1993),
.A2(n_1983),
.B(n_1977),
.Y(n_2008)
);

NAND4xp25_ASAP7_75t_L g2009 ( 
.A(n_1990),
.B(n_1984),
.C(n_1981),
.D(n_1973),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1998),
.B(n_1983),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1997),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1996),
.B(n_1887),
.Y(n_2012)
);

NOR2x1_ASAP7_75t_L g2013 ( 
.A(n_2001),
.B(n_1996),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_2003),
.B(n_1995),
.Y(n_2014)
);

NOR3xp33_ASAP7_75t_L g2015 ( 
.A(n_2004),
.B(n_1920),
.C(n_1902),
.Y(n_2015)
);

AOI211xp5_ASAP7_75t_L g2016 ( 
.A1(n_2008),
.A2(n_1999),
.B(n_1902),
.C(n_1922),
.Y(n_2016)
);

NOR3xp33_ASAP7_75t_L g2017 ( 
.A(n_2000),
.B(n_1922),
.C(n_1920),
.Y(n_2017)
);

NOR3xp33_ASAP7_75t_L g2018 ( 
.A(n_2002),
.B(n_1923),
.C(n_1922),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2006),
.Y(n_2019)
);

NAND3xp33_ASAP7_75t_L g2020 ( 
.A(n_2007),
.B(n_1925),
.C(n_1923),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2011),
.B(n_1882),
.Y(n_2021)
);

OAI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_2013),
.A2(n_2012),
.B1(n_2010),
.B2(n_2005),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_2016),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2021),
.Y(n_2024)
);

AOI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_2019),
.A2(n_2009),
.B1(n_1925),
.B2(n_1923),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2020),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2017),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2015),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_2014),
.A2(n_1925),
.B1(n_1882),
.B2(n_1876),
.Y(n_2029)
);

INVxp67_ASAP7_75t_SL g2030 ( 
.A(n_2018),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2023),
.B(n_1848),
.Y(n_2031)
);

AND3x1_ASAP7_75t_L g2032 ( 
.A(n_2025),
.B(n_2027),
.C(n_2026),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2030),
.Y(n_2033)
);

NOR3xp33_ASAP7_75t_L g2034 ( 
.A(n_2022),
.B(n_1877),
.C(n_1874),
.Y(n_2034)
);

NOR4xp75_ASAP7_75t_SL g2035 ( 
.A(n_2028),
.B(n_1887),
.C(n_1738),
.D(n_1877),
.Y(n_2035)
);

NAND2x1p5_ASAP7_75t_L g2036 ( 
.A(n_2024),
.B(n_2029),
.Y(n_2036)
);

NAND3x1_ASAP7_75t_L g2037 ( 
.A(n_2033),
.B(n_1876),
.C(n_1867),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_2031),
.Y(n_2038)
);

NOR2x1p5_ASAP7_75t_L g2039 ( 
.A(n_2032),
.B(n_1879),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_2036),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2037),
.Y(n_2041)
);

OAI222xp33_ASAP7_75t_L g2042 ( 
.A1(n_2041),
.A2(n_2040),
.B1(n_2038),
.B2(n_2035),
.C1(n_2039),
.C2(n_2034),
.Y(n_2042)
);

OA21x2_ASAP7_75t_L g2043 ( 
.A1(n_2042),
.A2(n_1850),
.B(n_1830),
.Y(n_2043)
);

INVx2_ASAP7_75t_SL g2044 ( 
.A(n_2042),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_SL g2045 ( 
.A1(n_2044),
.A2(n_1366),
.B1(n_1394),
.B2(n_1411),
.Y(n_2045)
);

AOI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_2043),
.A2(n_1850),
.B1(n_1787),
.B2(n_1825),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_2045),
.A2(n_2043),
.B1(n_1830),
.B2(n_1811),
.Y(n_2047)
);

AOI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_2046),
.A2(n_1868),
.B(n_1865),
.Y(n_2048)
);

AOI21xp33_ASAP7_75t_L g2049 ( 
.A1(n_2047),
.A2(n_1868),
.B(n_1865),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_SL g2050 ( 
.A1(n_2049),
.A2(n_2048),
.B1(n_1811),
.B2(n_1597),
.Y(n_2050)
);

AOI221xp5_ASAP7_75t_L g2051 ( 
.A1(n_2050),
.A2(n_1818),
.B1(n_1810),
.B2(n_1813),
.C(n_1823),
.Y(n_2051)
);

AOI211xp5_ASAP7_75t_L g2052 ( 
.A1(n_2051),
.A2(n_1597),
.B(n_1595),
.C(n_1596),
.Y(n_2052)
);


endmodule