module real_aes_7516_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_503;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_792;
wire n_1067;
wire n_878;
wire n_665;
wire n_991;
wire n_667;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_979;
wire n_759;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_1089;
wire n_857;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_1034;
wire n_376;
wire n_549;
wire n_571;
wire n_491;
wire n_894;
wire n_923;
wire n_694;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_884;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_1021;
wire n_399;
wire n_700;
wire n_1046;
wire n_958;
wire n_677;
wire n_948;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_815;
wire n_638;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_994;
wire n_495;
wire n_892;
wire n_1072;
wire n_370;
wire n_1078;
wire n_744;
wire n_384;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_1049;
wire n_559;
wire n_872;
wire n_636;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_931;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_962;
wire n_693;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_1017;
wire n_737;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_1006;
wire n_449;
wire n_363;
wire n_607;
wire n_417;
wire n_754;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_1031;
wire n_1037;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_1003;
wire n_533;
wire n_1000;
wire n_1014;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_649;
wire n_358;
wire n_385;
wire n_397;
wire n_749;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_1068;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_653;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_787;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_1102;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1101;
wire n_447;
wire n_603;
wire n_854;
wire n_403;
wire n_1039;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g572 ( .A1(n_0), .A2(n_260), .B1(n_573), .B2(n_574), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g1050 ( .A1(n_1), .A2(n_1051), .B1(n_1052), .B2(n_1068), .Y(n_1050) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_1), .Y(n_1068) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_2), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_3), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_4), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_5), .A2(n_48), .B1(n_744), .B2(n_1003), .Y(n_1002) );
AOI22x1_ASAP7_75t_L g862 ( .A1(n_6), .A2(n_863), .B1(n_895), .B2(n_896), .Y(n_862) );
INVx1_ASAP7_75t_L g895 ( .A(n_6), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_7), .A2(n_124), .B1(n_639), .B2(n_641), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_8), .Y(n_384) );
AO22x2_ASAP7_75t_L g373 ( .A1(n_9), .A2(n_205), .B1(n_374), .B2(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g1047 ( .A(n_9), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_10), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g1015 ( .A(n_11), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_12), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_13), .A2(n_265), .B1(n_497), .B2(n_532), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_14), .A2(n_84), .B1(n_779), .B2(n_905), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_15), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_16), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_17), .A2(n_225), .B1(n_648), .B2(n_649), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_18), .A2(n_142), .B1(n_697), .B2(n_746), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_19), .B(n_627), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_20), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_21), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g995 ( .A(n_22), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_23), .A2(n_328), .B1(n_457), .B2(n_854), .Y(n_1027) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_24), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_25), .Y(n_537) );
AOI222xp33_ASAP7_75t_L g951 ( .A1(n_26), .A2(n_50), .B1(n_314), .B2(n_583), .C1(n_763), .C2(n_952), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_27), .A2(n_112), .B1(n_429), .B2(n_433), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_28), .Y(n_848) );
AO22x2_ASAP7_75t_L g377 ( .A1(n_29), .A2(n_96), .B1(n_374), .B2(n_378), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_30), .A2(n_343), .B1(n_447), .B2(n_450), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_31), .A2(n_227), .B1(n_433), .B2(n_541), .Y(n_949) );
INVx1_ASAP7_75t_L g966 ( .A(n_32), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_33), .A2(n_101), .B1(n_640), .B2(n_657), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_34), .A2(n_148), .B1(n_604), .B2(n_989), .Y(n_988) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_35), .A2(n_251), .B1(n_438), .B2(n_641), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_36), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_37), .B(n_768), .Y(n_767) );
AOI22xp5_ASAP7_75t_SL g577 ( .A1(n_38), .A2(n_578), .B1(n_579), .B2(n_609), .Y(n_577) );
INVx1_ASAP7_75t_L g609 ( .A(n_38), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_39), .A2(n_128), .B1(n_536), .B2(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1096 ( .A(n_40), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_41), .A2(n_269), .B1(n_519), .B2(n_520), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_42), .A2(n_199), .B1(n_418), .B2(n_519), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_43), .A2(n_308), .B1(n_706), .B2(n_975), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_44), .A2(n_224), .B1(n_603), .B2(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_45), .B(n_791), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_46), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_47), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_49), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_51), .A2(n_261), .B1(n_652), .B2(n_655), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g898 ( .A1(n_52), .A2(n_899), .B1(n_924), .B2(n_925), .Y(n_898) );
INVx1_ASAP7_75t_L g924 ( .A(n_52), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_53), .A2(n_117), .B1(n_879), .B2(n_880), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_54), .B(n_627), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_55), .A2(n_294), .B1(n_909), .B2(n_991), .Y(n_990) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_56), .A2(n_618), .B1(n_658), .B2(n_659), .Y(n_617) );
INVx1_ASAP7_75t_L g658 ( .A(n_56), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_57), .A2(n_344), .B1(n_1006), .B2(n_1091), .Y(n_1090) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_58), .A2(n_250), .B1(n_702), .B2(n_703), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_59), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_60), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_61), .A2(n_275), .B1(n_652), .B2(n_872), .Y(n_977) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_62), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_63), .A2(n_90), .B1(n_370), .B2(n_433), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_64), .A2(n_85), .B1(n_854), .B2(n_856), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g1011 ( .A(n_65), .Y(n_1011) );
AOI222xp33_ASAP7_75t_L g743 ( .A1(n_66), .A2(n_255), .B1(n_312), .B2(n_583), .C1(n_627), .C2(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_67), .A2(n_236), .B1(n_519), .B2(n_520), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_68), .A2(n_268), .B1(n_495), .B2(n_498), .Y(n_950) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_69), .A2(n_194), .B1(n_628), .B2(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g662 ( .A(n_70), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g1016 ( .A(n_71), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_72), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_73), .A2(n_119), .B1(n_591), .B2(n_594), .Y(n_1008) );
AO22x2_ASAP7_75t_L g383 ( .A1(n_74), .A2(n_231), .B1(n_374), .B2(n_375), .Y(n_383) );
INVx1_ASAP7_75t_L g1044 ( .A(n_74), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g1056 ( .A(n_75), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_76), .A2(n_77), .B1(n_497), .B2(n_498), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_78), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_79), .A2(n_94), .B1(n_491), .B2(n_650), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_80), .A2(n_211), .B1(n_387), .B2(n_520), .Y(n_560) );
OA22x2_ASAP7_75t_L g504 ( .A1(n_81), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_81), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_82), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_83), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_86), .A2(n_304), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_87), .A2(n_131), .B1(n_393), .B2(n_586), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_88), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_89), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_91), .A2(n_168), .B1(n_524), .B2(n_697), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_92), .A2(n_196), .B1(n_648), .B2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g598 ( .A1(n_93), .A2(n_331), .B1(n_599), .B2(n_600), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_95), .A2(n_136), .B1(n_456), .B2(n_703), .Y(n_801) );
INVx1_ASAP7_75t_L g1048 ( .A(n_96), .Y(n_1048) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_97), .A2(n_153), .B1(n_478), .B2(n_524), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_98), .Y(n_1001) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_99), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_100), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_102), .A2(n_201), .B1(n_450), .B2(n_703), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_103), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_104), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_105), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_106), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_107), .A2(n_264), .B1(n_495), .B2(n_798), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_108), .A2(n_249), .B1(n_599), .B2(n_639), .Y(n_907) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_109), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_110), .A2(n_208), .B1(n_880), .B2(n_909), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_111), .A2(n_121), .B1(n_827), .B2(n_828), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_113), .A2(n_283), .B1(n_431), .B2(n_433), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_114), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_115), .A2(n_163), .B1(n_478), .B2(n_746), .Y(n_1061) );
AOI22xp33_ASAP7_75t_SL g1064 ( .A1(n_116), .A2(n_277), .B1(n_457), .B2(n_497), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_118), .A2(n_307), .B1(n_387), .B2(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_120), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_122), .A2(n_287), .B1(n_418), .B2(n_1021), .Y(n_1020) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_123), .A2(n_300), .B1(n_520), .B2(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_125), .A2(n_305), .B1(n_607), .B2(n_643), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_126), .A2(n_286), .B1(n_773), .B2(n_872), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_127), .A2(n_180), .B1(n_706), .B2(n_774), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_129), .A2(n_187), .B1(n_667), .B2(n_779), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_130), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_132), .B(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_133), .A2(n_184), .B1(n_438), .B2(n_441), .Y(n_437) );
AND2x6_ASAP7_75t_L g353 ( .A(n_134), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g1041 ( .A(n_134), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_135), .A2(n_257), .B1(n_457), .B2(n_643), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_137), .A2(n_218), .B1(n_639), .B2(n_825), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_138), .A2(n_252), .B1(n_393), .B2(n_1006), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_139), .A2(n_161), .B1(n_451), .B2(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g820 ( .A(n_140), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_141), .A2(n_239), .B1(n_491), .B2(n_492), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g1102 ( .A1(n_143), .A2(n_215), .B1(n_230), .B2(n_371), .C1(n_386), .C2(n_418), .Y(n_1102) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_144), .Y(n_838) );
INVx1_ASAP7_75t_L g1076 ( .A(n_145), .Y(n_1076) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_146), .A2(n_237), .B1(n_449), .B2(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_147), .A2(n_169), .B1(n_773), .B2(n_774), .Y(n_772) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_149), .A2(n_254), .B1(n_519), .B2(n_689), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g1024 ( .A(n_150), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_151), .A2(n_282), .B1(n_451), .B2(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g1060 ( .A(n_152), .B(n_738), .Y(n_1060) );
AO22x2_ASAP7_75t_L g381 ( .A1(n_154), .A2(n_220), .B1(n_374), .B2(n_378), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g1045 ( .A(n_154), .B(n_1046), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_155), .B(n_919), .Y(n_918) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_156), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_157), .A2(n_166), .B1(n_643), .B2(n_880), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g1067 ( .A1(n_158), .A2(n_235), .B1(n_536), .B2(n_604), .Y(n_1067) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_159), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g1028 ( .A1(n_160), .A2(n_327), .B1(n_652), .B2(n_655), .Y(n_1028) );
AOI22xp33_ASAP7_75t_SL g1057 ( .A1(n_162), .A2(n_246), .B1(n_520), .B2(n_628), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_164), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_165), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_167), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_170), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_171), .A2(n_207), .B1(n_650), .B2(n_734), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g1066 ( .A1(n_172), .A2(n_183), .B1(n_650), .B2(n_827), .Y(n_1066) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_173), .A2(n_213), .B1(n_497), .B2(n_570), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_174), .A2(n_209), .B1(n_591), .B2(n_594), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g954 ( .A1(n_175), .A2(n_955), .B1(n_978), .B2(n_979), .Y(n_954) );
INVx1_ASAP7_75t_L g978 ( .A(n_175), .Y(n_978) );
AOI22xp33_ASAP7_75t_SL g606 ( .A1(n_176), .A2(n_332), .B1(n_529), .B2(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g584 ( .A(n_177), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_178), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_179), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g953 ( .A(n_181), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_182), .A2(n_338), .B1(n_497), .B2(n_532), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_185), .A2(n_267), .B1(n_531), .B2(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g1098 ( .A(n_186), .Y(n_1098) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_188), .A2(n_276), .B1(n_449), .B2(n_702), .Y(n_800) );
AOI22xp33_ASAP7_75t_SL g1063 ( .A1(n_189), .A2(n_325), .B1(n_447), .B2(n_643), .Y(n_1063) );
CKINVDCx20_ASAP7_75t_R g945 ( .A(n_190), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_191), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g700 ( .A1(n_192), .A2(n_234), .B1(n_433), .B2(n_495), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_193), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_195), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_197), .A2(n_204), .B1(n_628), .B2(n_845), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_198), .A2(n_306), .B1(n_431), .B2(n_603), .Y(n_1029) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_200), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_202), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_203), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_206), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_210), .A2(n_298), .B1(n_497), .B2(n_532), .Y(n_608) );
INVx1_ASAP7_75t_L g1094 ( .A(n_212), .Y(n_1094) );
OA22x2_ASAP7_75t_L g465 ( .A1(n_214), .A2(n_466), .B1(n_467), .B2(n_499), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_214), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_216), .B(n_739), .Y(n_1059) );
XNOR2x2_ASAP7_75t_L g984 ( .A(n_217), .B(n_985), .Y(n_984) );
INVx2_ASAP7_75t_L g358 ( .A(n_219), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_221), .A2(n_233), .B1(n_429), .B2(n_652), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_222), .B(n_594), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_223), .Y(n_916) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_226), .A2(n_346), .B1(n_456), .B2(n_570), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g993 ( .A(n_228), .Y(n_993) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_229), .A2(n_341), .B1(n_641), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_232), .A2(n_319), .B1(n_479), .B2(n_689), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_238), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_240), .A2(n_280), .B1(n_449), .B2(n_649), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_241), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_242), .A2(n_336), .B1(n_643), .B2(n_645), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_243), .B(n_766), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_244), .A2(n_712), .B1(n_747), .B2(n_748), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_244), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_245), .A2(n_342), .B1(n_441), .B2(n_536), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_247), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_248), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_253), .A2(n_278), .B1(n_455), .B2(n_457), .Y(n_454) );
INVx1_ASAP7_75t_L g374 ( .A(n_256), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_256), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_258), .A2(n_340), .B1(n_433), .B2(n_491), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_259), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_262), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_263), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g913 ( .A(n_266), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_270), .Y(n_809) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_271), .A2(n_351), .B(n_359), .C(n_1049), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_272), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_273), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_274), .Y(n_887) );
INVx1_ASAP7_75t_L g912 ( .A(n_279), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_281), .B(n_766), .Y(n_946) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_284), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_285), .A2(n_335), .B1(n_573), .B2(n_574), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_288), .A2(n_303), .B1(n_431), .B2(n_971), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_289), .A2(n_324), .B1(n_495), .B2(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_290), .A2(n_311), .B1(n_395), .B2(n_479), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_291), .Y(n_963) );
INVx1_ASAP7_75t_L g357 ( .A(n_292), .Y(n_357) );
INVx1_ASAP7_75t_L g967 ( .A(n_293), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_295), .Y(n_813) );
INVx1_ASAP7_75t_L g354 ( .A(n_296), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g997 ( .A(n_297), .Y(n_997) );
INVx1_ASAP7_75t_L g1100 ( .A(n_299), .Y(n_1100) );
OA22x2_ASAP7_75t_L g682 ( .A1(n_301), .A2(n_683), .B1(n_684), .B2(n_708), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_301), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_302), .B(n_695), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_309), .Y(n_1019) );
CKINVDCx20_ASAP7_75t_R g998 ( .A(n_310), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_313), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_315), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_316), .Y(n_815) );
INVx1_ASAP7_75t_L g860 ( .A(n_317), .Y(n_860) );
INVx1_ASAP7_75t_L g1086 ( .A(n_318), .Y(n_1086) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_320), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_321), .B(n_393), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_322), .Y(n_922) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_323), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_326), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_329), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_330), .B(n_1089), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_333), .Y(n_719) );
INVx1_ASAP7_75t_L g576 ( .A(n_334), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_337), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_339), .B(n_628), .Y(n_964) );
OA22x2_ASAP7_75t_SL g804 ( .A1(n_345), .A2(n_805), .B1(n_806), .B2(n_832), .Y(n_804) );
INVx1_ASAP7_75t_L g832 ( .A(n_345), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_347), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_348), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g962 ( .A(n_349), .Y(n_962) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_353), .B(n_355), .Y(n_352) );
HB1xp67_ASAP7_75t_L g1040 ( .A(n_354), .Y(n_1040) );
OA21x2_ASAP7_75t_L g1074 ( .A1(n_355), .A2(n_1039), .B(n_1075), .Y(n_1074) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_752), .B1(n_1034), .B2(n_1035), .C(n_1036), .Y(n_359) );
INVx1_ASAP7_75t_L g1034 ( .A(n_360), .Y(n_1034) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B1(n_500), .B2(n_751), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_462), .B2(n_463), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
XOR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_461), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_426), .Y(n_366) );
NOR3xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_399), .C(n_415), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_384), .B1(n_385), .B2(n_391), .C(n_392), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g760 ( .A1(n_369), .A2(n_761), .B(n_762), .Y(n_760) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_SL g888 ( .A(n_370), .Y(n_888) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g517 ( .A(n_371), .Y(n_517) );
INVx4_ASAP7_75t_L g558 ( .A(n_371), .Y(n_558) );
INVx2_ASAP7_75t_L g786 ( .A(n_371), .Y(n_786) );
INVx2_ASAP7_75t_SL g915 ( .A(n_371), .Y(n_915) );
INVx2_ASAP7_75t_L g961 ( .A(n_371), .Y(n_961) );
AND2x6_ASAP7_75t_L g371 ( .A(n_372), .B(n_379), .Y(n_371) );
AND2x4_ASAP7_75t_L g396 ( .A(n_372), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g485 ( .A(n_372), .Y(n_485) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_377), .Y(n_372) );
AND2x2_ASAP7_75t_L g390 ( .A(n_373), .B(n_381), .Y(n_390) );
INVx2_ASAP7_75t_L g406 ( .A(n_373), .Y(n_406) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_376), .Y(n_378) );
OR2x2_ASAP7_75t_L g405 ( .A(n_377), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g414 ( .A(n_377), .B(n_406), .Y(n_414) );
INVx2_ASAP7_75t_L g421 ( .A(n_377), .Y(n_421) );
INVx1_ASAP7_75t_L g460 ( .A(n_377), .Y(n_460) );
AND2x6_ASAP7_75t_L g431 ( .A(n_379), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g440 ( .A(n_379), .B(n_436), .Y(n_440) );
AND2x4_ASAP7_75t_L g449 ( .A(n_379), .B(n_414), .Y(n_449) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
AND2x2_ASAP7_75t_L g408 ( .A(n_380), .B(n_383), .Y(n_408) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g435 ( .A(n_381), .B(n_398), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_381), .B(n_383), .Y(n_444) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g389 ( .A(n_383), .Y(n_389) );
INVx1_ASAP7_75t_L g398 ( .A(n_383), .Y(n_398) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx4f_ASAP7_75t_L g1003 ( .A(n_386), .Y(n_1003) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx12f_ASAP7_75t_L g519 ( .A(n_387), .Y(n_519) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_387), .Y(n_628) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g420 ( .A(n_389), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g419 ( .A(n_390), .B(n_420), .Y(n_419) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_390), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g479 ( .A(n_390), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_SL g520 ( .A(n_396), .Y(n_520) );
BUFx2_ASAP7_75t_SL g763 ( .A(n_396), .Y(n_763) );
BUFx3_ASAP7_75t_L g1091 ( .A(n_396), .Y(n_1091) );
INVx1_ASAP7_75t_L g486 ( .A(n_397), .Y(n_486) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_409), .B2(n_410), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_401), .A2(n_410), .B1(n_883), .B2(n_884), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_401), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g471 ( .A(n_404), .Y(n_471) );
INVx2_ASAP7_75t_L g511 ( .A(n_404), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g671 ( .A1(n_404), .A2(n_412), .B1(n_672), .B2(n_673), .C(n_674), .Y(n_671) );
OR2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
INVx2_ASAP7_75t_L g432 ( .A(n_405), .Y(n_432) );
AND2x2_ASAP7_75t_L g436 ( .A(n_406), .B(n_421), .Y(n_436) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_408), .B(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g456 ( .A(n_408), .B(n_436), .Y(n_456) );
AND2x4_ASAP7_75t_L g593 ( .A(n_408), .B(n_432), .Y(n_593) );
AND2x6_ASAP7_75t_L g595 ( .A(n_408), .B(n_414), .Y(n_595) );
OAI22xp5_ASAP7_75t_SL g509 ( .A1(n_410), .A2(n_510), .B1(n_512), .B2(n_513), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_410), .A2(n_510), .B1(n_621), .B2(n_622), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_410), .A2(n_809), .B1(n_810), .B2(n_811), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_410), .A2(n_838), .B1(n_839), .B2(n_840), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_410), .A2(n_471), .B1(n_958), .B2(n_959), .Y(n_957) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx3_ASAP7_75t_L g1087 ( .A(n_412), .Y(n_1087) );
BUFx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g474 ( .A(n_413), .Y(n_474) );
AND2x2_ASAP7_75t_L g453 ( .A(n_414), .B(n_435), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_414), .B(n_435), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B1(n_422), .B2(n_423), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_418), .Y(n_564) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g492 ( .A(n_419), .Y(n_492) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_419), .Y(n_524) );
BUFx4f_ASAP7_75t_SL g689 ( .A(n_419), .Y(n_689) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_419), .Y(n_746) );
INVx1_ASAP7_75t_L g425 ( .A(n_421), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_423), .A2(n_522), .B1(n_523), .B2(n_525), .Y(n_521) );
BUFx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_424), .A2(n_562), .B1(n_563), .B2(n_565), .Y(n_561) );
INVx4_ASAP7_75t_L g632 ( .A(n_424), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_424), .A2(n_484), .B1(n_741), .B2(n_742), .Y(n_740) );
AND2x2_ASAP7_75t_L g667 ( .A(n_425), .B(n_443), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_445), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_437), .Y(n_427) );
INVx2_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
OAI21xp33_ASAP7_75t_SL g475 ( .A1(n_430), .A2(n_476), .B(n_477), .Y(n_475) );
INVx3_ASAP7_75t_L g599 ( .A(n_430), .Y(n_599) );
INVx4_ASAP7_75t_L g641 ( .A(n_430), .Y(n_641) );
INVx4_ASAP7_75t_L g827 ( .A(n_430), .Y(n_827) );
INVx11_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx11_ASAP7_75t_L g542 ( .A(n_431), .Y(n_542) );
BUFx2_ASAP7_75t_L g903 ( .A(n_433), .Y(n_903) );
INVx1_ASAP7_75t_L g976 ( .A(n_433), .Y(n_976) );
BUFx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g601 ( .A(n_434), .Y(n_601) );
BUFx3_ASAP7_75t_L g650 ( .A(n_434), .Y(n_650) );
BUFx3_ASAP7_75t_L g774 ( .A(n_434), .Y(n_774) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_435), .B(n_436), .Y(n_547) );
AND2x4_ASAP7_75t_L g442 ( .A(n_436), .B(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_L g716 ( .A(n_438), .Y(n_716) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g495 ( .A(n_439), .Y(n_495) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_SL g536 ( .A(n_440), .Y(n_536) );
BUFx2_ASAP7_75t_SL g603 ( .A(n_440), .Y(n_603) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_440), .Y(n_640) );
INVx1_ASAP7_75t_SL g538 ( .A(n_441), .Y(n_538) );
BUFx2_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
BUFx3_ASAP7_75t_L g498 ( .A(n_442), .Y(n_498) );
BUFx2_ASAP7_75t_L g570 ( .A(n_442), .Y(n_570) );
BUFx2_ASAP7_75t_SL g604 ( .A(n_442), .Y(n_604) );
BUFx3_ASAP7_75t_L g657 ( .A(n_442), .Y(n_657) );
BUFx3_ASAP7_75t_L g798 ( .A(n_442), .Y(n_798) );
BUFx3_ASAP7_75t_L g828 ( .A(n_442), .Y(n_828) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x6_ASAP7_75t_L g459 ( .A(n_444), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_454), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g573 ( .A(n_448), .Y(n_573) );
INVx2_ASAP7_75t_L g607 ( .A(n_448), .Y(n_607) );
INVx3_ASAP7_75t_L g706 ( .A(n_448), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_448), .A2(n_545), .B1(n_997), .B2(n_998), .Y(n_996) );
INVx6_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx3_ASAP7_75t_L g491 ( .A(n_449), .Y(n_491) );
BUFx3_ASAP7_75t_L g648 ( .A(n_449), .Y(n_648) );
BUFx3_ASAP7_75t_L g875 ( .A(n_449), .Y(n_875) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g879 ( .A(n_451), .Y(n_879) );
INVx5_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g529 ( .A(n_452), .Y(n_529) );
INVx3_ASAP7_75t_L g574 ( .A(n_452), .Y(n_574) );
BUFx3_ASAP7_75t_L g644 ( .A(n_452), .Y(n_644) );
INVx4_ASAP7_75t_L g702 ( .A(n_452), .Y(n_702) );
INVx8_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx3_ASAP7_75t_L g497 ( .A(n_456), .Y(n_497) );
BUFx3_ASAP7_75t_L g531 ( .A(n_456), .Y(n_531) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_456), .Y(n_654) );
INVx2_ASAP7_75t_L g780 ( .A(n_456), .Y(n_780) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g532 ( .A(n_458), .Y(n_532) );
BUFx2_ASAP7_75t_L g645 ( .A(n_458), .Y(n_645) );
BUFx4f_ASAP7_75t_SL g880 ( .A(n_458), .Y(n_880) );
BUFx2_ASAP7_75t_L g991 ( .A(n_458), .Y(n_991) );
INVx6_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_459), .A2(n_482), .B1(n_483), .B2(n_484), .Y(n_481) );
INVx1_ASAP7_75t_SL g703 ( .A(n_459), .Y(n_703) );
INVx1_ASAP7_75t_L g856 ( .A(n_459), .Y(n_856) );
INVx1_ASAP7_75t_L g480 ( .A(n_460), .Y(n_480) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g499 ( .A(n_467), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_487), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_475), .C(n_481), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_471), .A2(n_554), .B1(n_555), .B2(n_556), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_473), .A2(n_810), .B1(n_912), .B2(n_913), .Y(n_911) );
OA211x2_ASAP7_75t_L g944 ( .A1(n_473), .A2(n_945), .B(n_946), .C(n_947), .Y(n_944) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g556 ( .A(n_474), .Y(n_556) );
INVx2_ASAP7_75t_L g1017 ( .A(n_474), .Y(n_1017) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx3_ASAP7_75t_L g697 ( .A(n_479), .Y(n_697) );
INVx1_ASAP7_75t_L g1007 ( .A(n_479), .Y(n_1007) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_479), .Y(n_1021) );
CKINVDCx16_ASAP7_75t_R g635 ( .A(n_484), .Y(n_635) );
BUFx2_ASAP7_75t_L g821 ( .A(n_484), .Y(n_821) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_493), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_497), .Y(n_869) );
INVxp67_ASAP7_75t_L g1095 ( .A(n_498), .Y(n_1095) );
INVx1_ASAP7_75t_L g751 ( .A(n_500), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_612), .B1(n_749), .B2(n_750), .Y(n_500) );
INVx1_ASAP7_75t_L g749 ( .A(n_501), .Y(n_749) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_548), .B2(n_611), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_526), .Y(n_507) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_514), .C(n_521), .Y(n_508) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g810 ( .A(n_511), .Y(n_810) );
INVx1_ASAP7_75t_SL g839 ( .A(n_511), .Y(n_839) );
OAI21xp33_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_518), .Y(n_514) );
OAI21xp5_ASAP7_75t_SL g675 ( .A1(n_516), .A2(n_676), .B(n_677), .Y(n_675) );
OAI21xp5_ASAP7_75t_SL g686 ( .A1(n_516), .A2(n_687), .B(n_688), .Y(n_686) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g587 ( .A(n_519), .Y(n_587) );
BUFx4f_ASAP7_75t_SL g952 ( .A(n_519), .Y(n_952) );
OAI221xp5_ASAP7_75t_SL g623 ( .A1(n_523), .A2(n_582), .B1(n_624), .B2(n_625), .C(n_626), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_533), .C(n_539), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
INVx1_ASAP7_75t_L g736 ( .A(n_531), .Y(n_736) );
BUFx2_ASAP7_75t_L g825 ( .A(n_531), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_537), .B2(n_538), .Y(n_533) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx5_ASAP7_75t_SL g734 ( .A(n_542), .Y(n_734) );
INVx4_ASAP7_75t_L g773 ( .A(n_542), .Y(n_773) );
OAI221xp5_ASAP7_75t_SL g873 ( .A1(n_545), .A2(n_874), .B1(n_876), .B2(n_877), .C(n_878), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_545), .A2(n_1094), .B1(n_1095), .B2(n_1096), .Y(n_1093) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g729 ( .A(n_546), .Y(n_729) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g611 ( .A(n_548), .Y(n_611) );
OA22x2_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_577), .B2(n_610), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
XOR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_576), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_566), .Y(n_551) );
NOR3xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .C(n_561), .Y(n_552) );
OAI21xp5_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_559), .B(n_560), .Y(n_557) );
INVx4_ASAP7_75t_L g583 ( .A(n_558), .Y(n_583) );
BUFx2_ASAP7_75t_L g843 ( .A(n_558), .Y(n_843) );
OAI221xp5_ASAP7_75t_L g960 ( .A1(n_563), .A2(n_961), .B1(n_962), .B2(n_963), .C(n_964), .Y(n_960) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_SL g886 ( .A(n_564), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_571), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
INVxp67_ASAP7_75t_L g727 ( .A(n_573), .Y(n_727) );
INVx1_ASAP7_75t_L g610 ( .A(n_577), .Y(n_610) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_580), .B(n_596), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_588), .Y(n_580) );
OAI21xp5_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_584), .B(n_585), .Y(n_581) );
OAI221xp5_ASAP7_75t_L g812 ( .A1(n_582), .A2(n_813), .B1(n_814), .B2(n_815), .C(n_816), .Y(n_812) );
OAI21xp33_ASAP7_75t_SL g1018 ( .A1(n_582), .A2(n_1019), .B(n_1020), .Y(n_1018) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx5_ASAP7_75t_L g695 ( .A(n_592), .Y(n_695) );
INVx2_ASAP7_75t_L g766 ( .A(n_592), .Y(n_766) );
INVx2_ASAP7_75t_L g791 ( .A(n_592), .Y(n_791) );
INVx4_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
BUFx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g693 ( .A(n_595), .Y(n_693) );
BUFx2_ASAP7_75t_L g739 ( .A(n_595), .Y(n_739) );
BUFx4f_ASAP7_75t_L g768 ( .A(n_595), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_605), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_602), .Y(n_597) );
INVx1_ASAP7_75t_L g1099 ( .A(n_599), .Y(n_1099) );
BUFx4f_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g750 ( .A(n_612), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_678), .B2(n_679), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_617), .B1(n_660), .B2(n_661), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g659 ( .A(n_618), .Y(n_659) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_636), .Y(n_618) );
NOR3xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_623), .C(n_629), .Y(n_619) );
INVx2_ASAP7_75t_L g890 ( .A(n_627), .Y(n_890) );
BUFx3_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g920 ( .A(n_628), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_633), .B2(n_634), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_631), .A2(n_847), .B1(n_848), .B2(n_849), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_631), .A2(n_821), .B1(n_966), .B2(n_967), .Y(n_965) );
INVx3_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g819 ( .A(n_632), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_634), .A2(n_819), .B1(n_893), .B2(n_894), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_634), .A2(n_819), .B1(n_922), .B2(n_923), .Y(n_921) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g849 ( .A(n_635), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_646), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_642), .Y(n_637) );
BUFx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx3_ASAP7_75t_L g866 ( .A(n_640), .Y(n_866) );
BUFx3_ASAP7_75t_L g971 ( .A(n_640), .Y(n_971) );
BUFx6f_ASAP7_75t_L g989 ( .A(n_640), .Y(n_989) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVxp67_ASAP7_75t_L g723 ( .A(n_645), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_651), .Y(n_646) );
BUFx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx4_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_653), .A2(n_993), .B1(n_994), .B2(n_995), .Y(n_992) );
INVx3_ASAP7_75t_L g1083 ( .A(n_653), .Y(n_1083) );
INVx4_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_656), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_714) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_657), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_660), .A2(n_661), .B1(n_682), .B2(n_709), .Y(n_681) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
XNOR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NOR4xp75_ASAP7_75t_L g663 ( .A(n_664), .B(n_668), .C(n_671), .D(n_675), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI22xp5_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_681), .B1(n_710), .B2(n_711), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g709 ( .A(n_682), .Y(n_709) );
INVx1_ASAP7_75t_L g708 ( .A(n_684), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_698), .Y(n_684) );
NOR2xp67_ASAP7_75t_L g685 ( .A(n_686), .B(n_690), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .C(n_696), .Y(n_690) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_695), .Y(n_738) );
NOR2x1_ASAP7_75t_L g698 ( .A(n_699), .B(n_704), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx2_ASAP7_75t_L g855 ( .A(n_702), .Y(n_855) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_702), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g1101 ( .A(n_706), .Y(n_1101) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g748 ( .A(n_712), .Y(n_748) );
AND4x1_ASAP7_75t_L g712 ( .A(n_713), .B(n_724), .C(n_737), .D(n_743), .Y(n_712) );
NOR2xp33_ASAP7_75t_SL g713 ( .A(n_714), .B(n_718), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B1(n_722), .B2(n_723), .Y(n_718) );
BUFx2_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_730), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_735), .B2(n_736), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g994 ( .A(n_734), .Y(n_994) );
INVx3_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx4_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g814 ( .A(n_746), .Y(n_814) );
BUFx2_ASAP7_75t_L g845 ( .A(n_746), .Y(n_845) );
INVx1_ASAP7_75t_L g1035 ( .A(n_752), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_932), .B1(n_933), .B2(n_1033), .Y(n_752) );
INVx1_ASAP7_75t_L g1033 ( .A(n_753), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_833), .B1(n_930), .B2(n_931), .Y(n_753) );
INVx2_ASAP7_75t_SL g930 ( .A(n_754), .Y(n_930) );
XNOR2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_804), .Y(n_754) );
OAI22x1_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B1(n_782), .B2(n_803), .Y(n_755) );
INVx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
XOR2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_781), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_759), .B(n_770), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_764), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_767), .C(n_769), .Y(n_764) );
NOR2x1_ASAP7_75t_L g770 ( .A(n_771), .B(n_776), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_775), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx3_ASAP7_75t_L g803 ( .A(n_782), .Y(n_803) );
XOR2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_802), .Y(n_782) );
NAND2x1_ASAP7_75t_SL g783 ( .A(n_784), .B(n_794), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_789), .Y(n_784) );
OAI21xp5_ASAP7_75t_SL g785 ( .A1(n_786), .A2(n_787), .B(n_788), .Y(n_785) );
OAI21xp5_ASAP7_75t_SL g1000 ( .A1(n_786), .A2(n_1001), .B(n_1002), .Y(n_1000) );
NAND3xp33_ASAP7_75t_L g789 ( .A(n_790), .B(n_792), .C(n_793), .Y(n_789) );
BUFx2_ASAP7_75t_L g1089 ( .A(n_791), .Y(n_1089) );
NOR2x1_ASAP7_75t_L g794 ( .A(n_795), .B(n_799), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
BUFx2_ASAP7_75t_L g905 ( .A(n_798), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_SL g806 ( .A(n_807), .B(n_822), .Y(n_806) );
NOR3xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_812), .C(n_817), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_819), .B1(n_820), .B2(n_821), .Y(n_817) );
OAI22xp5_ASAP7_75t_SL g1022 ( .A1(n_821), .A2(n_920), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_829), .Y(n_822) );
NAND2xp5_ASAP7_75t_SL g823 ( .A(n_824), .B(n_826), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
INVx1_ASAP7_75t_L g931 ( .A(n_833), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_861), .B1(n_928), .B2(n_929), .Y(n_833) );
INVx1_ASAP7_75t_L g928 ( .A(n_834), .Y(n_928) );
XOR2x2_ASAP7_75t_L g834 ( .A(n_835), .B(n_860), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_850), .Y(n_835) );
NOR3xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_841), .C(n_846), .Y(n_836) );
OAI21xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B(n_844), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_857), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
INVx3_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
INVx1_ASAP7_75t_L g929 ( .A(n_861), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_897), .B1(n_926), .B2(n_927), .Y(n_861) );
INVx2_ASAP7_75t_L g926 ( .A(n_862), .Y(n_926) );
INVx1_ASAP7_75t_SL g896 ( .A(n_863), .Y(n_896) );
AND2x2_ASAP7_75t_SL g863 ( .A(n_864), .B(n_881), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_873), .Y(n_864) );
OAI221xp5_ASAP7_75t_SL g865 ( .A1(n_866), .A2(n_867), .B1(n_868), .B2(n_870), .C(n_871), .Y(n_865) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx3_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NOR3xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_885), .C(n_892), .Y(n_881) );
OAI222xp33_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_887), .B1(n_888), .B2(n_889), .C1(n_890), .C2(n_891), .Y(n_885) );
OAI221xp5_ASAP7_75t_L g914 ( .A1(n_886), .A2(n_915), .B1(n_916), .B2(n_917), .C(n_918), .Y(n_914) );
INVx2_ASAP7_75t_L g927 ( .A(n_897), .Y(n_927) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g925 ( .A(n_899), .Y(n_925) );
AND2x2_ASAP7_75t_SL g899 ( .A(n_900), .B(n_910), .Y(n_899) );
NOR2xp33_ASAP7_75t_SL g900 ( .A(n_901), .B(n_906), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
NOR3xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_914), .C(n_921), .Y(n_910) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
AOI22xp5_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_981), .B1(n_982), .B2(n_1032), .Y(n_933) );
INVx1_ASAP7_75t_SL g1032 ( .A(n_934), .Y(n_1032) );
BUFx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
OAI22xp5_ASAP7_75t_SL g935 ( .A1(n_936), .A2(n_937), .B1(n_954), .B2(n_980), .Y(n_935) );
INVx1_ASAP7_75t_SL g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
XNOR2xp5_ASAP7_75t_L g1009 ( .A(n_938), .B(n_1010), .Y(n_1009) );
INVx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
XOR2x2_ASAP7_75t_L g939 ( .A(n_940), .B(n_953), .Y(n_939) );
NAND4xp75_ASAP7_75t_L g940 ( .A(n_941), .B(n_944), .C(n_948), .D(n_951), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_942), .B(n_943), .Y(n_941) );
AND2x2_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
INVx1_ASAP7_75t_L g980 ( .A(n_954), .Y(n_980) );
INVx2_ASAP7_75t_L g979 ( .A(n_955), .Y(n_979) );
AND2x2_ASAP7_75t_SL g955 ( .A(n_956), .B(n_968), .Y(n_955) );
NOR3xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_960), .C(n_965), .Y(n_956) );
OAI21xp5_ASAP7_75t_SL g1055 ( .A1(n_961), .A2(n_1056), .B(n_1057), .Y(n_1055) );
NOR2xp33_ASAP7_75t_L g968 ( .A(n_969), .B(n_973), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_970), .B(n_972), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_974), .B(n_977), .Y(n_973) );
INVx2_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g983 ( .A1(n_984), .A2(n_1009), .B1(n_1030), .B2(n_1031), .Y(n_983) );
INVx2_ASAP7_75t_L g1030 ( .A(n_984), .Y(n_1030) );
NAND2xp5_ASAP7_75t_SL g985 ( .A(n_986), .B(n_999), .Y(n_985) );
NOR3xp33_ASAP7_75t_L g986 ( .A(n_987), .B(n_992), .C(n_996), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_988), .B(n_990), .Y(n_987) );
NOR2xp33_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1004), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1008), .Y(n_1004) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1009), .Y(n_1031) );
XNOR2x1_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1025), .Y(n_1012) );
NOR3xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1018), .C(n_1022), .Y(n_1013) );
AND4x1_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .C(n_1028), .D(n_1029), .Y(n_1025) );
INVx1_ASAP7_75t_SL g1036 ( .A(n_1037), .Y(n_1036) );
NOR2x1_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1042), .Y(n_1037) );
OR2x2_ASAP7_75t_SL g1105 ( .A(n_1038), .B(n_1043), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1041), .Y(n_1038) );
CKINVDCx20_ASAP7_75t_R g1071 ( .A(n_1039), .Y(n_1071) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_1040), .B(n_1073), .Y(n_1075) );
CKINVDCx16_ASAP7_75t_R g1073 ( .A(n_1041), .Y(n_1073) );
CKINVDCx20_ASAP7_75t_R g1042 ( .A(n_1043), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1048), .Y(n_1046) );
OAI322xp33_ASAP7_75t_L g1049 ( .A1(n_1050), .A2(n_1069), .A3(n_1072), .B1(n_1074), .B2(n_1076), .C1(n_1077), .C2(n_1103), .Y(n_1049) );
CKINVDCx20_ASAP7_75t_R g1051 ( .A(n_1052), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
NAND3x1_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1062), .C(n_1065), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1058), .Y(n_1054) );
NAND3xp33_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1060), .C(n_1061), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1067), .Y(n_1065) );
HB1xp67_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
HB1xp67_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
XOR2x2_ASAP7_75t_L g1079 ( .A(n_1076), .B(n_1080), .Y(n_1079) );
INVx1_ASAP7_75t_SL g1077 ( .A(n_1078), .Y(n_1077) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
NAND4xp75_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1085), .C(n_1092), .D(n_1102), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1084), .Y(n_1081) );
OA211x2_ASAP7_75t_L g1085 ( .A1(n_1086), .A2(n_1087), .B(n_1088), .C(n_1090), .Y(n_1085) );
NOR2xp33_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1097), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_1098), .A2(n_1099), .B1(n_1100), .B2(n_1101), .Y(n_1097) );
CKINVDCx20_ASAP7_75t_R g1103 ( .A(n_1104), .Y(n_1103) );
CKINVDCx20_ASAP7_75t_R g1104 ( .A(n_1105), .Y(n_1104) );
endmodule