module fake_jpeg_28504_n_549 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_549);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_549;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_0),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_54),
.Y(n_168)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_57),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_62),
.Y(n_162)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_21),
.B(n_9),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_68),
.Y(n_115)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_21),
.B(n_9),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

CKINVDCx6p67_ASAP7_75t_R g125 ( 
.A(n_69),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_9),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_86),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g138 ( 
.A(n_76),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_20),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_80),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_20),
.B(n_9),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_10),
.B1(n_17),
.B2(n_16),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_84),
.A2(n_35),
.B1(n_36),
.B2(n_44),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_8),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_40),
.B(n_7),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_105),
.Y(n_126)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_103),
.Y(n_166)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_19),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_54),
.A2(n_38),
.B1(n_91),
.B2(n_37),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_114),
.A2(n_143),
.B1(n_152),
.B2(n_107),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_56),
.A2(n_49),
.B1(n_33),
.B2(n_52),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_116),
.A2(n_144),
.B1(n_0),
.B2(n_1),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_124),
.B(n_127),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_57),
.B(n_42),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_43),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_140),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_43),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_87),
.B(n_42),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_157),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_104),
.A2(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_63),
.B(n_44),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_158),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_67),
.A2(n_74),
.B1(n_58),
.B2(n_62),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_88),
.B(n_35),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_53),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_92),
.B(n_41),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_37),
.Y(n_194)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_171),
.Y(n_261)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_114),
.A2(n_84),
.B1(n_69),
.B2(n_36),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_172),
.B(n_178),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_125),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_173),
.B(n_186),
.Y(n_268)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

AO22x2_ASAP7_75t_SL g177 ( 
.A1(n_116),
.A2(n_94),
.B1(n_97),
.B2(n_99),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_177),
.A2(n_135),
.B(n_136),
.C(n_123),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_119),
.B(n_76),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_128),
.A2(n_31),
.B1(n_53),
.B2(n_41),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_179),
.A2(n_198),
.B1(n_217),
.B2(n_222),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_180),
.A2(n_224),
.B1(n_168),
.B2(n_153),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_76),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_182),
.B(n_191),
.C(n_204),
.Y(n_240)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_112),
.A2(n_77),
.B1(n_64),
.B2(n_71),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_184),
.A2(n_192),
.B1(n_201),
.B2(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_125),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_125),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_187),
.B(n_188),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_137),
.A2(n_75),
.B1(n_83),
.B2(n_85),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_190),
.A2(n_28),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_110),
.B(n_100),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_115),
.A2(n_23),
.B1(n_29),
.B2(n_31),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_126),
.B(n_122),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_215),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_128),
.A2(n_34),
.B1(n_29),
.B2(n_37),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_149),
.A2(n_34),
.B1(n_45),
.B2(n_37),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_200),
.B(n_209),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_143),
.A2(n_154),
.B1(n_121),
.B2(n_136),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_202),
.Y(n_277)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_103),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_52),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_205),
.A2(n_208),
.B(n_129),
.Y(n_242)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_141),
.B(n_52),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_108),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_138),
.Y(n_210)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_108),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_168),
.Y(n_233)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_212),
.Y(n_267)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_121),
.A2(n_52),
.B1(n_32),
.B2(n_45),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_147),
.B(n_45),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_216),
.Y(n_271)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_218),
.A2(n_11),
.B1(n_18),
.B2(n_15),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_150),
.B(n_22),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_219),
.A2(n_220),
.B(n_0),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_155),
.A2(n_45),
.B1(n_22),
.B2(n_28),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_111),
.B(n_45),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_225),
.Y(n_248)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_223),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_138),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_111),
.B(n_45),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_117),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_117),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_133),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_233),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_235),
.B(n_242),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_241),
.A2(n_255),
.B1(n_262),
.B2(n_193),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_178),
.A2(n_129),
.B1(n_159),
.B2(n_138),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_243),
.B(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_177),
.A2(n_123),
.B1(n_162),
.B2(n_164),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_245),
.A2(n_257),
.B1(n_275),
.B2(n_220),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_189),
.A2(n_133),
.B(n_135),
.Y(n_249)
);

OAI31xp33_ASAP7_75t_SL g322 ( 
.A1(n_249),
.A2(n_11),
.A3(n_12),
.B(n_3),
.Y(n_322)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_189),
.B(n_164),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_252),
.B(n_253),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_162),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_177),
.A2(n_22),
.B1(n_102),
.B2(n_28),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_181),
.B(n_22),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_259),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_188),
.B(n_22),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_174),
.A2(n_10),
.B(n_18),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_260),
.B(n_5),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_218),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_200),
.B1(n_185),
.B2(n_199),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_178),
.B(n_28),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_204),
.C(n_202),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_172),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_274),
.B(n_182),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_172),
.A2(n_15),
.B1(n_5),
.B2(n_6),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_197),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_279),
.B(n_309),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_170),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_292),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_281),
.A2(n_320),
.B1(n_254),
.B2(n_251),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_282),
.A2(n_286),
.B1(n_288),
.B2(n_299),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_283),
.A2(n_233),
.B1(n_273),
.B2(n_242),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_284),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_290),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_234),
.A2(n_270),
.B1(n_245),
.B2(n_248),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_291),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_244),
.B(n_225),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_268),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_294),
.Y(n_327)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_236),
.Y(n_295)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_206),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_301),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_234),
.A2(n_172),
.B1(n_221),
.B2(n_195),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g300 ( 
.A1(n_244),
.A2(n_196),
.A3(n_208),
.B1(n_203),
.B2(n_205),
.Y(n_300)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_248),
.B(n_191),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_243),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_302),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_239),
.A2(n_207),
.B1(n_212),
.B2(n_226),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_303),
.A2(n_230),
.B1(n_232),
.B2(n_264),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_270),
.A2(n_208),
.B1(n_205),
.B2(n_191),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_304),
.A2(n_306),
.B1(n_312),
.B2(n_313),
.Y(n_343)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_236),
.Y(n_305)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_305),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_270),
.A2(n_213),
.B1(n_176),
.B2(n_222),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_252),
.B(n_182),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_316),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_235),
.A2(n_229),
.B1(n_228),
.B2(n_227),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_278),
.A2(n_204),
.B1(n_217),
.B2(n_216),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_314),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_175),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_315),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_183),
.C(n_223),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_261),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_317),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_258),
.B(n_171),
.Y(n_319)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_253),
.C(n_259),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_275),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_3),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_240),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_322),
.A2(n_264),
.B(n_256),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_323),
.B(n_301),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_293),
.A2(n_298),
.B(n_249),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_324),
.A2(n_362),
.B(n_313),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_280),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_325),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_328),
.Y(n_397)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_308),
.A2(n_249),
.B1(n_237),
.B2(n_241),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_329),
.A2(n_346),
.B1(n_354),
.B2(n_304),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g330 ( 
.A(n_322),
.B(n_276),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g388 ( 
.A1(n_330),
.A2(n_337),
.B(n_287),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_SL g337 ( 
.A1(n_282),
.A2(n_241),
.B(n_255),
.C(n_265),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_345),
.A2(n_309),
.B1(n_310),
.B2(n_294),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_297),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_355),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_293),
.A2(n_240),
.B(n_247),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_351),
.A2(n_356),
.B(n_360),
.Y(n_381)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_353),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_285),
.A2(n_262),
.B1(n_246),
.B2(n_232),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_315),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_317),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_284),
.Y(n_385)
);

AO22x1_ASAP7_75t_SL g359 ( 
.A1(n_285),
.A2(n_246),
.B1(n_267),
.B2(n_269),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_291),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_293),
.A2(n_298),
.B(n_321),
.Y(n_360)
);

OAI32xp33_ASAP7_75t_L g361 ( 
.A1(n_292),
.A2(n_267),
.A3(n_263),
.B1(n_269),
.B2(n_238),
.Y(n_361)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_298),
.A2(n_321),
.B(n_308),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_279),
.C(n_319),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_372),
.C(n_387),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_364),
.A2(n_382),
.B1(n_343),
.B2(n_332),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_331),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_371),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_366),
.B(n_359),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_340),
.A2(n_288),
.B1(n_299),
.B2(n_307),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_368),
.A2(n_380),
.B1(n_390),
.B2(n_392),
.Y(n_405)
);

AOI221xp5_ASAP7_75t_L g400 ( 
.A1(n_370),
.A2(n_339),
.B1(n_355),
.B2(n_361),
.C(n_332),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_327),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_341),
.B(n_352),
.Y(n_372)
);

OAI21xp33_ASAP7_75t_SL g425 ( 
.A1(n_373),
.A2(n_388),
.B(n_337),
.Y(n_425)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_324),
.A2(n_316),
.B(n_312),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_375),
.A2(n_378),
.B(n_393),
.Y(n_407)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_356),
.A2(n_306),
.B(n_283),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_340),
.A2(n_307),
.B1(n_310),
.B2(n_286),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_346),
.A2(n_320),
.B1(n_300),
.B2(n_289),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_395),
.Y(n_414)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_335),
.Y(n_384)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_384),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_385),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_296),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_341),
.B(n_311),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_323),
.B(n_271),
.C(n_318),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_328),
.C(n_362),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_348),
.A2(n_314),
.B1(n_284),
.B2(n_271),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_326),
.B(n_314),
.Y(n_391)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_391),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_348),
.A2(n_266),
.B1(n_305),
.B2(n_295),
.Y(n_392)
);

XOR2x2_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_266),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_326),
.B(n_238),
.Y(n_394)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_394),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_350),
.B(n_263),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_343),
.A2(n_317),
.B1(n_231),
.B2(n_261),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_396),
.A2(n_344),
.B1(n_357),
.B2(n_336),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_400),
.A2(n_426),
.B1(n_427),
.B2(n_365),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_404),
.A2(n_408),
.B1(n_417),
.B2(n_423),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_364),
.A2(n_337),
.B1(n_339),
.B2(n_360),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_412),
.C(n_413),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_381),
.A2(n_333),
.B(n_334),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_411),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_328),
.C(n_342),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_342),
.C(n_357),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_415),
.B(n_419),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_382),
.A2(n_337),
.B1(n_354),
.B2(n_338),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_418),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_363),
.Y(n_419)
);

NAND3xp33_ASAP7_75t_L g420 ( 
.A(n_367),
.B(n_330),
.C(n_358),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_370),
.Y(n_439)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_359),
.Y(n_422)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_369),
.A2(n_337),
.B1(n_338),
.B2(n_347),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_379),
.B(n_347),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_424),
.B(n_376),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_378),
.B1(n_373),
.B2(n_375),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_369),
.A2(n_344),
.B1(n_349),
.B2(n_336),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_395),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_429),
.B(n_391),
.Y(n_431)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_431),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_418),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_432),
.B(n_442),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_434),
.A2(n_438),
.B1(n_455),
.B2(n_405),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_393),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_440),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_417),
.A2(n_368),
.B1(n_380),
.B2(n_390),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_439),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_393),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_389),
.C(n_387),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_444),
.C(n_449),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_421),
.B(n_394),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_381),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_415),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_366),
.C(n_397),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_424),
.Y(n_445)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_445),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_383),
.Y(n_446)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_446),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_401),
.B(n_392),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_423),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_397),
.C(n_396),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_406),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_385),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_451),
.A2(n_404),
.B1(n_428),
.B2(n_403),
.Y(n_472)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_398),
.Y(n_454)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_454),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_408),
.A2(n_397),
.B1(n_377),
.B2(n_388),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_433),
.A2(n_438),
.B1(n_445),
.B2(n_405),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_458),
.A2(n_471),
.B1(n_451),
.B2(n_436),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_474),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_472),
.Y(n_491)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_467),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_429),
.Y(n_468)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_468),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_452),
.A2(n_431),
.B(n_446),
.Y(n_470)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_470),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_403),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_430),
.B(n_407),
.C(n_428),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_449),
.C(n_441),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_440),
.B(n_407),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_477),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_443),
.B(n_411),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_398),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_437),
.B(n_427),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_448),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_484),
.C(n_488),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_482),
.A2(n_377),
.B1(n_399),
.B2(n_384),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_430),
.C(n_444),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_465),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_448),
.C(n_436),
.Y(n_488)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_489),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_434),
.C(n_433),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_496),
.C(n_476),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_388),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_497),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_474),
.A2(n_450),
.B(n_402),
.Y(n_493)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_493),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_459),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_457),
.B(n_416),
.C(n_414),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_414),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_501),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_477),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_509),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_491),
.B(n_485),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_495),
.A2(n_471),
.B1(n_474),
.B2(n_463),
.Y(n_502)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_502),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_481),
.A2(n_461),
.B1(n_462),
.B2(n_464),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_503),
.B(n_377),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_486),
.A2(n_468),
.B(n_472),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_505),
.A2(n_496),
.B(n_399),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_12),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_480),
.B(n_416),
.C(n_422),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_509),
.C(n_498),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_490),
.A2(n_470),
.B(n_473),
.Y(n_511)
);

AOI21x1_ASAP7_75t_L g518 ( 
.A1(n_511),
.A2(n_512),
.B(n_497),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_487),
.A2(n_426),
.B(n_402),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_513),
.A2(n_231),
.B1(n_11),
.B2(n_12),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_514),
.B(n_523),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_518),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_484),
.C(n_488),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_501),
.C(n_500),
.Y(n_532)
);

AOI21xp33_ASAP7_75t_L g519 ( 
.A1(n_504),
.A2(n_483),
.B(n_492),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_519),
.A2(n_522),
.B(n_526),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_508),
.A2(n_374),
.B(n_349),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_525),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_12),
.Y(n_526)
);

A2O1A1Ixp33_ASAP7_75t_L g529 ( 
.A1(n_520),
.A2(n_507),
.B(n_512),
.C(n_502),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_529),
.B(n_532),
.Y(n_537)
);

NOR2xp67_ASAP7_75t_SL g531 ( 
.A(n_516),
.B(n_503),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_531),
.A2(n_521),
.B(n_524),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_498),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_533),
.A2(n_535),
.B(n_515),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_517),
.B(n_499),
.C(n_505),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_536),
.B(n_538),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_528),
.A2(n_523),
.B(n_521),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_539),
.B(n_540),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_534),
.B(n_4),
.Y(n_540)
);

OAI31xp33_ASAP7_75t_SL g541 ( 
.A1(n_537),
.A2(n_529),
.A3(n_527),
.B(n_530),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_541),
.B(n_542),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_533),
.C(n_527),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_544),
.B(n_545),
.C(n_4),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_4),
.C(n_371),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_4),
.Y(n_548)
);

BUFx24_ASAP7_75t_SL g549 ( 
.A(n_548),
.Y(n_549)
);


endmodule