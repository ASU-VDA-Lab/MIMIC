module fake_jpeg_31618_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx4_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_19),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_17),
.B(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_24),
.Y(n_26)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

AO22x2_ASAP7_75t_SL g24 ( 
.A1(n_13),
.A2(n_8),
.B1(n_11),
.B2(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_9),
.Y(n_30)
);

AOI322xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_24),
.A3(n_10),
.B1(n_11),
.B2(n_18),
.C1(n_20),
.C2(n_23),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.C(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_24),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_36),
.B(n_33),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_29),
.B1(n_28),
.B2(n_3),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_39),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_35),
.B(n_7),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_11),
.C(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_0),
.B(n_1),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_7),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_0),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_49),
.B(n_4),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_4),
.B1(n_5),
.B2(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_48),
.Y(n_51)
);


endmodule