module fake_jpeg_16734_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_0),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_SL g7 ( 
.A(n_0),
.B(n_1),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_8),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_15)
);

OAI32xp33_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_19),
.A3(n_23),
.B1(n_13),
.B2(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_18),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_6),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_7),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_11),
.A2(n_14),
.B1(n_9),
.B2(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx24_ASAP7_75t_SL g33 ( 
.A(n_26),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_11),
.B1(n_30),
.B2(n_27),
.Y(n_36)
);

AOI322xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_22),
.A3(n_15),
.B1(n_20),
.B2(n_18),
.C1(n_16),
.C2(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_35),
.B(n_28),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_38),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_32),
.B1(n_11),
.B2(n_27),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.B(n_38),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_39),
.B(n_31),
.Y(n_44)
);


endmodule