module real_jpeg_12316_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_4),
.A2(n_22),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_4),
.A2(n_22),
.B1(n_29),
.B2(n_30),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_4),
.A2(n_22),
.B1(n_40),
.B2(n_42),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_4),
.B(n_27),
.C(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_4),
.B(n_28),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_4),
.B(n_45),
.C(n_52),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_4),
.B(n_37),
.C(n_42),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_4),
.B(n_117),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_6),
.A2(n_40),
.B1(n_42),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_90),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_88),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_70),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_14),
.B(n_70),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_56),
.C(n_67),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_15),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_32),
.B2(n_33),
.Y(n_15)
);

AOI211xp5_ASAP7_75t_SL g73 ( 
.A1(n_16),
.A2(n_35),
.B(n_74),
.C(n_75),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_16),
.A2(n_17),
.B1(n_48),
.B2(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_49),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_23),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_22),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_22),
.B(n_61),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

AO22x1_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_30),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_30),
.B(n_98),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_32),
.A2(n_33),
.B1(n_94),
.B2(n_95),
.Y(n_132)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_34),
.B(n_49),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_34),
.A2(n_35),
.B1(n_78),
.B2(n_82),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_34),
.A2(n_49),
.B(n_94),
.C(n_99),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_34),
.A2(n_35),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_34),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_34),
.A2(n_35),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_34),
.A2(n_35),
.B1(n_111),
.B2(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_35),
.B(n_66),
.C(n_115),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_35),
.B(n_101),
.C(n_105),
.Y(n_140)
);

OA21x2_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_43),
.B(n_47),
.Y(n_35)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

AO22x1_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g42 ( 
.A(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_40),
.B(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_61),
.Y(n_62)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OA22x2_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_46),
.B1(n_52),
.B2(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_45),
.B(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_66),
.C(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_48),
.A2(n_49),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_55),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_56),
.A2(n_57),
.B1(n_67),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_58),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_66),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_58),
.A2(n_66),
.B1(n_114),
.B2(n_118),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_58),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_62),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_66),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_66),
.B(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_66),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_66),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_83),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_136),
.B(n_141),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_107),
.B(n_135),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_100),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_131),
.B(n_134),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_119),
.B(n_130),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_140),
.Y(n_141)
);


endmodule