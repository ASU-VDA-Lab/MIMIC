module fake_jpeg_19084_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_21),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_17),
.B(n_27),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_55),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_51),
.B1(n_57),
.B2(n_18),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_32),
.B1(n_24),
.B2(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_32),
.B1(n_23),
.B2(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_71),
.B(n_73),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_18),
.B1(n_30),
.B2(n_21),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_72),
.A2(n_86),
.B1(n_25),
.B2(n_66),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_74),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_17),
.B(n_27),
.C(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_82),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_63),
.B1(n_56),
.B2(n_31),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_81),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_45),
.B1(n_44),
.B2(n_41),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_97),
.B1(n_98),
.B2(n_102),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_30),
.B1(n_23),
.B2(n_25),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_35),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_93),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_40),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_26),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_62),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_45),
.B1(n_44),
.B2(n_41),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_1),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_31),
.Y(n_144)
);

AOI22x1_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_69),
.B1(n_80),
.B2(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_98),
.B1(n_84),
.B2(n_102),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_130),
.B1(n_78),
.B2(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_63),
.B1(n_43),
.B2(n_31),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_127),
.B1(n_74),
.B2(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_20),
.B1(n_16),
.B2(n_22),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_31),
.B1(n_19),
.B2(n_20),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_132),
.A2(n_140),
.B1(n_149),
.B2(n_106),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_138),
.B1(n_145),
.B2(n_146),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_135),
.B(n_150),
.Y(n_194)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_139),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_96),
.B1(n_74),
.B2(n_78),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_75),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_91),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_148),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_70),
.B1(n_95),
.B2(n_87),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_70),
.B1(n_90),
.B2(n_94),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_79),
.B1(n_85),
.B2(n_92),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_158),
.B1(n_162),
.B2(n_2),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_83),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_79),
.B1(n_85),
.B2(n_19),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_89),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_20),
.C(n_16),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_155),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_19),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_152),
.B(n_161),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_20),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_105),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_19),
.C(n_22),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_22),
.C(n_15),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_11),
.Y(n_180)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_104),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_158)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_128),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_15),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_104),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_113),
.B(n_112),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_108),
.B(n_118),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_171),
.B(n_173),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_108),
.B1(n_118),
.B2(n_109),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_179),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_106),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_170),
.A2(n_182),
.B(n_197),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_109),
.B(n_107),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_174),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_113),
.B(n_129),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_180),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_137),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_135),
.A2(n_105),
.B1(n_112),
.B2(n_124),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_183),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_124),
.Y(n_182)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_107),
.A3(n_119),
.B1(n_110),
.B2(n_14),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_185),
.A2(n_133),
.B1(n_137),
.B2(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_133),
.B(n_110),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_188),
.B1(n_154),
.B2(n_160),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_13),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_3),
.C(n_5),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_156),
.B(n_13),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_193),
.B(n_6),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_132),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_149),
.B1(n_151),
.B2(n_134),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_163),
.A2(n_10),
.B1(n_12),
.B2(n_5),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_163),
.B(n_158),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_197),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_162),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_198),
.A2(n_199),
.B(n_210),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_201),
.A2(n_207),
.B1(n_214),
.B2(n_195),
.Y(n_241)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_209),
.A2(n_164),
.B1(n_170),
.B2(n_182),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_170),
.A2(n_139),
.B(n_160),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_212),
.A2(n_225),
.B(n_175),
.Y(n_245)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_180),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_223),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_174),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_167),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_179),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_168),
.A2(n_6),
.B(n_7),
.Y(n_225)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_178),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_231),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_185),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_238),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_178),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_176),
.B1(n_184),
.B2(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_173),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_233),
.B(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_192),
.Y(n_237)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_172),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_240),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_205),
.A2(n_165),
.B1(n_169),
.B2(n_190),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_207),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_188),
.B1(n_168),
.B2(n_181),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_244),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_190),
.B1(n_191),
.B2(n_166),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_245),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_196),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_246),
.B(n_198),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_189),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_251),
.A2(n_241),
.B1(n_230),
.B2(n_206),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_203),
.B1(n_219),
.B2(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_253),
.B(n_239),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_255),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_220),
.C(n_212),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_257),
.C(n_263),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_222),
.C(n_221),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_217),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_226),
.B(n_200),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_264),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_217),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_240),
.C(n_244),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_262),
.Y(n_269)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_275),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_249),
.B1(n_266),
.B2(n_243),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_272),
.A2(n_247),
.B1(n_238),
.B2(n_225),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_235),
.B(n_236),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_278),
.Y(n_289)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_R g279 ( 
.A(n_259),
.B(n_235),
.C(n_199),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_263),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_282),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_265),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_258),
.A2(n_228),
.B(n_227),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_284),
.A2(n_198),
.B(n_245),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_288),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_257),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_261),
.C(n_256),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_297),
.C(n_278),
.Y(n_300)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_293),
.A2(n_270),
.B1(n_274),
.B2(n_276),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_279),
.B(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_281),
.B(n_250),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_261),
.C(n_250),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_273),
.A2(n_253),
.B1(n_214),
.B2(n_218),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_303),
.C(n_291),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_269),
.B(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_277),
.C(n_284),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_306),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_305),
.A2(n_307),
.B(n_286),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_285),
.A2(n_275),
.B(n_7),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_287),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_313),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_299),
.B(n_301),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_305),
.A2(n_289),
.B(n_290),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_315),
.B(n_300),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_290),
.Y(n_315)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_310),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_309),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_318),
.C(n_313),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_320),
.B(n_319),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_295),
.B(n_297),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_8),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_9),
.C(n_296),
.Y(n_327)
);


endmodule