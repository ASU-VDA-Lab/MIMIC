module fake_jpeg_26376_n_298 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_298);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_288;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_12),
.B(n_9),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

HAxp5_ASAP7_75t_SL g35 ( 
.A(n_12),
.B(n_11),
.CON(n_35),
.SN(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_21),
.B1(n_15),
.B2(n_12),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_53),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_30),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_15),
.B1(n_21),
.B2(n_24),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_24),
.B1(n_25),
.B2(n_20),
.Y(n_87)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_27),
.B1(n_32),
.B2(n_29),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_27),
.B1(n_46),
.B2(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_40),
.B(n_15),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_39),
.B1(n_40),
.B2(n_27),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_75),
.B1(n_81),
.B2(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_33),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_39),
.B1(n_29),
.B2(n_32),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_26),
.C(n_34),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_31),
.C(n_34),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_87),
.A2(n_24),
.B1(n_61),
.B2(n_20),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_92),
.B1(n_99),
.B2(n_110),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_63),
.B(n_48),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_107),
.B(n_109),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_90),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_48),
.B1(n_64),
.B2(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_95),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_56),
.B1(n_61),
.B2(n_66),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_108),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_104),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_52),
.B1(n_17),
.B2(n_60),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_52),
.B1(n_17),
.B2(n_35),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_26),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_26),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_38),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_17),
.B1(n_34),
.B2(n_13),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_82),
.B1(n_76),
.B2(n_77),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_25),
.B(n_23),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_23),
.B1(n_25),
.B2(n_13),
.Y(n_108)
);

OA21x2_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_77),
.B(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_26),
.B1(n_16),
.B2(n_13),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_111),
.A2(n_84),
.B1(n_70),
.B2(n_76),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_115),
.B(n_119),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_118),
.B1(n_122),
.B2(n_140),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_85),
.B1(n_87),
.B2(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_84),
.B(n_69),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_100),
.B(n_102),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_69),
.B1(n_70),
.B2(n_83),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_19),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_131),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_136),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_69),
.B(n_11),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_139),
.B(n_108),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_22),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_26),
.C(n_38),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_19),
.C(n_18),
.Y(n_168)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_137),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_105),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_80),
.B1(n_57),
.B2(n_18),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_80),
.B1(n_18),
.B2(n_16),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_89),
.A2(n_8),
.B(n_9),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_91),
.A2(n_93),
.B1(n_105),
.B2(n_101),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_134),
.A3(n_123),
.B1(n_137),
.B2(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_145),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_89),
.B(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_163),
.Y(n_180)
);

AOI32xp33_ASAP7_75t_SL g156 ( 
.A1(n_129),
.A2(n_107),
.A3(n_88),
.B1(n_110),
.B2(n_96),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_112),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_98),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_162),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_80),
.B1(n_16),
.B2(n_13),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_22),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_122),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_80),
.B1(n_18),
.B2(n_16),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_164),
.A2(n_22),
.B1(n_19),
.B2(n_2),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_8),
.B(n_9),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_167),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_115),
.A2(n_7),
.B(n_9),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_124),
.C(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_193),
.C(n_168),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_144),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_186),
.Y(n_204)
);

XOR2x2_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_130),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_156),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_182),
.B1(n_197),
.B2(n_159),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_130),
.B1(n_112),
.B2(n_114),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_22),
.Y(n_192)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_80),
.C(n_19),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_171),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_194),
.B(n_154),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_206),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_219),
.B(n_198),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_158),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_170),
.C(n_169),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_214),
.C(n_218),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_209),
.A2(n_165),
.B1(n_173),
.B2(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_213),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_157),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_212),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_143),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_153),
.Y(n_218)
);

OAI22x1_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_148),
.B1(n_165),
.B2(n_166),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_150),
.C(n_149),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_185),
.C(n_178),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_229),
.B1(n_237),
.B2(n_181),
.Y(n_241)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_184),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_228),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_212),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_219),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_173),
.B1(n_179),
.B2(n_184),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_233),
.B(n_235),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_178),
.C(n_200),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_251),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_207),
.C(n_208),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_242),
.B(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_226),
.C(n_185),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_246),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_205),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_249),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_211),
.C(n_191),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_214),
.C(n_181),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_226),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_188),
.B1(n_195),
.B2(n_176),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_197),
.B1(n_144),
.B2(n_189),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_252),
.A2(n_228),
.B1(n_227),
.B2(n_225),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_264),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_232),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_254),
.B(n_256),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_248),
.A2(n_236),
.B(n_224),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_6),
.B(n_1),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_221),
.B1(n_223),
.B2(n_186),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_262),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_221),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_257),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_189),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_0),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_243),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_270),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_260),
.A2(n_244),
.B1(n_240),
.B2(n_167),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_0),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_164),
.B1(n_6),
.B2(n_19),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_271),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_SL g271 ( 
.A(n_264),
.B(n_19),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_6),
.B(n_1),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_0),
.B(n_1),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_0),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_6),
.C(n_1),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_279),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_283),
.B(n_2),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_0),
.B(n_2),
.Y(n_282)
);

OAI321xp33_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_284),
.A3(n_271),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_2),
.B(n_3),
.Y(n_284)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_3),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_272),
.B(n_273),
.C(n_5),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_277),
.C(n_4),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.C(n_285),
.Y(n_294)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_280),
.B(n_286),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_293),
.A2(n_294),
.B1(n_3),
.B2(n_4),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_3),
.C(n_4),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_4),
.C(n_5),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_5),
.Y(n_298)
);


endmodule