module fake_jpeg_2424_n_187 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_187);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_64),
.B1(n_53),
.B2(n_60),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_57),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_64),
.B1(n_53),
.B2(n_61),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_53),
.B1(n_61),
.B2(n_55),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_55),
.B1(n_59),
.B2(n_63),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_85),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_72),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_90),
.Y(n_102)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_72),
.C(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_0),
.Y(n_106)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_56),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_65),
.C(n_78),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_65),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_7),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_32),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_70),
.B1(n_68),
.B2(n_81),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_121),
.B1(n_85),
.B2(n_25),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_109),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_70),
.B(n_58),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_115),
.Y(n_124)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_58),
.B1(n_2),
.B2(n_3),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_4),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_134),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_112),
.C(n_105),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_118),
.C(n_111),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_8),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_139),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_140),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_124),
.B1(n_133),
.B2(n_129),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_151),
.B1(n_29),
.B2(n_30),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_139),
.A2(n_114),
.B(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_149),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_118),
.B1(n_13),
.B2(n_21),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_17),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_125),
.B1(n_23),
.B2(n_27),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_162),
.B(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_22),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_165),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_28),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_155),
.B1(n_145),
.B2(n_152),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_164),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_33),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_149),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_169),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_154),
.C(n_153),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_153),
.C(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_163),
.C(n_157),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_176),
.Y(n_180)
);

AOI31xp67_ASAP7_75t_SL g181 ( 
.A1(n_180),
.A2(n_171),
.A3(n_174),
.B(n_173),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_179),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_172),
.C(n_35),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_46),
.C(n_39),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_34),
.C(n_40),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_41),
.B(n_42),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_45),
.Y(n_187)
);


endmodule