module fake_jpeg_3093_n_171 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_42),
.Y(n_71)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_75),
.Y(n_87)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_82),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_56),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_85),
.C(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_44),
.C(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_91),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_50),
.C(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_47),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_43),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_101),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_64),
.B1(n_51),
.B2(n_47),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_83),
.B1(n_90),
.B2(n_86),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_57),
.A3(n_54),
.B1(n_52),
.B2(n_65),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_7),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_51),
.C(n_65),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_62),
.C(n_60),
.Y(n_116)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_0),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_113),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_62),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_115),
.Y(n_136)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_55),
.B(n_1),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_120),
.B(n_107),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_121),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_0),
.B(n_1),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_2),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_129),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_24),
.C(n_40),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_103),
.C(n_27),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_131),
.B(n_19),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_8),
.B(n_9),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_116),
.B1(n_23),
.B2(n_25),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_146),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_26),
.C(n_39),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_141),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_143),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_132),
.B1(n_115),
.B2(n_120),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_20),
.Y(n_146)
);

AOI221xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_130),
.B1(n_126),
.B2(n_123),
.C(n_117),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_155),
.B1(n_137),
.B2(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_147),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_156),
.B(n_158),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_140),
.C(n_134),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_160),
.B(n_151),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_136),
.B(n_153),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_149),
.B(n_152),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_164),
.A2(n_165),
.B(n_163),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_156),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_144),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_144),
.C(n_28),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_21),
.A3(n_29),
.B1(n_30),
.B2(n_31),
.C1(n_32),
.C2(n_34),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_35),
.B(n_36),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_38),
.Y(n_171)
);


endmodule