module fake_jpeg_943_n_480 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_480);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_480;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_46),
.Y(n_156)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_47),
.Y(n_138)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_65),
.Y(n_120)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_13),
.Y(n_64)
);

CKINVDCx12_ASAP7_75t_R g118 ( 
.A(n_64),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_38),
.B(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_78),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_15),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_38),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_83),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_22),
.B(n_6),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_36),
.B(n_4),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_89),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_12),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_15),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_98),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_103),
.B(n_114),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_41),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_34),
.B1(n_43),
.B2(n_45),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_39),
.B1(n_44),
.B2(n_89),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_52),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_37),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_146),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_57),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_74),
.B(n_26),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_18),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_71),
.B(n_26),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_54),
.B(n_37),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_56),
.B(n_41),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_159),
.Y(n_237)
);

INVx5_ASAP7_75t_SL g161 ( 
.A(n_118),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_131),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_98),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_133),
.C(n_138),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_134),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_172),
.B(n_182),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_70),
.B1(n_97),
.B2(n_90),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_139),
.B1(n_150),
.B2(n_129),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_22),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_177),
.Y(n_209)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_126),
.B(n_44),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_186),
.Y(n_212)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_181),
.A2(n_185),
.B1(n_188),
.B2(n_193),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_134),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_184),
.A2(n_195),
.B1(n_201),
.B2(n_204),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_121),
.A2(n_42),
.B1(n_45),
.B2(n_30),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_121),
.B(n_120),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_190),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_42),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_191),
.B(n_192),
.Y(n_228)
);

CKINVDCx12_ASAP7_75t_R g192 ( 
.A(n_145),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_196),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_146),
.A2(n_66),
.B1(n_86),
.B2(n_81),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_197),
.A2(n_199),
.B1(n_156),
.B2(n_137),
.Y(n_232)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_200),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_106),
.B(n_40),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_102),
.A2(n_77),
.B1(n_69),
.B2(n_63),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_203),
.Y(n_227)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_142),
.A2(n_45),
.B1(n_30),
.B2(n_40),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_139),
.B1(n_129),
.B2(n_60),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_213),
.B1(n_217),
.B2(n_222),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_171),
.C(n_175),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_119),
.C(n_155),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_214),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_151),
.C(n_148),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_138),
.B1(n_127),
.B2(n_153),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_131),
.B1(n_84),
.B2(n_147),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_160),
.B(n_133),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_232),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_189),
.A2(n_55),
.B1(n_49),
.B2(n_113),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_242),
.Y(n_290)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_161),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_227),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_249),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_209),
.B(n_177),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_254),
.Y(n_269)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_212),
.A2(n_231),
.B(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_223),
.Y(n_250)
);

NAND2xp33_ASAP7_75t_SL g277 ( 
.A(n_250),
.B(n_260),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_189),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_253),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_171),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_210),
.B(n_164),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_255),
.A2(n_257),
.B1(n_261),
.B2(n_238),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_227),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_256),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_180),
.B(n_101),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_258),
.A2(n_263),
.B(n_264),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_218),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_223),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_218),
.B(n_169),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_226),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_208),
.A2(n_203),
.B(n_165),
.Y(n_263)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_186),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_205),
.B(n_179),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_266),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_232),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_276),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_246),
.A2(n_236),
.B1(n_213),
.B2(n_222),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_272),
.A2(n_273),
.B1(n_279),
.B2(n_281),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_252),
.A2(n_256),
.B1(n_241),
.B2(n_240),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_205),
.C(n_237),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_221),
.B1(n_206),
.B2(n_207),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_240),
.A2(n_206),
.B1(n_221),
.B2(n_228),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_287),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_241),
.A2(n_183),
.B1(n_191),
.B2(n_163),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_254),
.A2(n_188),
.B1(n_200),
.B2(n_162),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_255),
.Y(n_303)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_229),
.C(n_220),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_220),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_255),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_294),
.Y(n_312)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_299),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_SL g300 ( 
.A1(n_274),
.A2(n_251),
.B(n_253),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_300),
.A2(n_302),
.B(n_287),
.Y(n_328)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_301),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_268),
.A2(n_258),
.B(n_250),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_311),
.Y(n_337)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_304),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_277),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_286),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_285),
.B(n_247),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_306),
.B(n_314),
.Y(n_331)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_307),
.Y(n_323)
);

BUFx8_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_290),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_264),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_276),
.C(n_271),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_230),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_283),
.A2(n_257),
.B1(n_248),
.B2(n_243),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_294),
.B1(n_281),
.B2(n_272),
.Y(n_349)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_319),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_268),
.B(n_257),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_317),
.B(n_318),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_261),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_287),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_285),
.B(n_260),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_288),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_324),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_320),
.A2(n_286),
.B1(n_269),
.B2(n_274),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_325),
.A2(n_340),
.B1(n_299),
.B2(n_279),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_312),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_335),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_328),
.A2(n_333),
.B(n_310),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_317),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_307),
.B(n_269),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_338),
.B(n_309),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_339),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_320),
.A2(n_297),
.B1(n_299),
.B2(n_303),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_318),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_341),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_313),
.B(n_273),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_344),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_315),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_345),
.A2(n_349),
.B1(n_278),
.B2(n_248),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_346),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_305),
.Y(n_348)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_348),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_350),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_361),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_357),
.A2(n_370),
.B(n_328),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_342),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_358),
.B(n_375),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_338),
.B(n_296),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_323),
.B(n_267),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_374),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_364),
.A2(n_365),
.B1(n_368),
.B2(n_330),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_340),
.A2(n_302),
.B1(n_321),
.B2(n_310),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_325),
.A2(n_321),
.B1(n_295),
.B2(n_298),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_329),
.Y(n_369)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_369),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g370 ( 
.A(n_324),
.B(n_304),
.Y(n_370)
);

AO22x1_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_311),
.B1(n_282),
.B2(n_290),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_371),
.Y(n_390)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_372),
.Y(n_376)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_334),
.Y(n_373)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_282),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_326),
.Y(n_379)
);

NAND3xp33_ASAP7_75t_L g408 ( 
.A(n_379),
.B(n_392),
.C(n_215),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_380),
.A2(n_394),
.B1(n_397),
.B2(n_353),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_371),
.Y(n_381)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_381),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_350),
.C(n_336),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_386),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_357),
.A2(n_336),
.B(n_335),
.Y(n_385)
);

OAI321xp33_ASAP7_75t_L g401 ( 
.A1(n_385),
.A2(n_352),
.A3(n_359),
.B1(n_360),
.B2(n_355),
.C(n_370),
.Y(n_401)
);

NOR2x1_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_342),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_356),
.A2(n_349),
.B1(n_337),
.B2(n_343),
.Y(n_387)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_365),
.A2(n_337),
.B(n_343),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_389),
.B(n_393),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_366),
.B(n_347),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_362),
.B(n_327),
.C(n_347),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_L g394 ( 
.A1(n_368),
.A2(n_327),
.B1(n_346),
.B2(n_278),
.Y(n_394)
);

OA22x2_ASAP7_75t_L g396 ( 
.A1(n_364),
.A2(n_198),
.B1(n_243),
.B2(n_242),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_238),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_358),
.A2(n_261),
.B1(n_242),
.B2(n_229),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_361),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_403),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_385),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_408),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_401),
.A2(n_381),
.B(n_389),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_391),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_410),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_395),
.A2(n_363),
.B1(n_353),
.B2(n_354),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_407),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_261),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_409),
.B(n_411),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_377),
.B(n_215),
.C(n_233),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_414),
.Y(n_426)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_388),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_233),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_415),
.B(n_416),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_382),
.B(n_202),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_417),
.A2(n_157),
.B1(n_123),
.B2(n_98),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_386),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_422),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_405),
.A2(n_395),
.B(n_390),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_421),
.A2(n_181),
.B(n_72),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_394),
.C(n_396),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_396),
.C(n_383),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_425),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_396),
.C(n_383),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_412),
.A2(n_376),
.B1(n_390),
.B2(n_397),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_429),
.B(n_431),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_404),
.A2(n_376),
.B1(n_196),
.B2(n_176),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_170),
.C(n_154),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_433),
.C(n_34),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_415),
.C(n_407),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_420),
.A2(n_406),
.B1(n_410),
.B2(n_197),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_436),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_19),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_420),
.A2(n_19),
.B1(n_28),
.B2(n_18),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_438),
.B(n_440),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_96),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_34),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_441),
.A2(n_438),
.B(n_46),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_443),
.A2(n_447),
.B(n_46),
.Y(n_456)
);

INVx6_ASAP7_75t_L g444 ( 
.A(n_430),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_444),
.B(n_422),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_433),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_SL g450 ( 
.A(n_445),
.B(n_446),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_157),
.C(n_123),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_424),
.A2(n_157),
.B(n_96),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_452),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_423),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_451),
.A2(n_456),
.B(n_449),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_430),
.C(n_425),
.Y(n_452)
);

OAI221xp5_ASAP7_75t_L g453 ( 
.A1(n_437),
.A2(n_426),
.B1(n_428),
.B2(n_8),
.C(n_3),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_453),
.A2(n_435),
.B(n_446),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_455),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_457),
.B(n_458),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_442),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_459),
.A2(n_462),
.B(n_465),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_454),
.B(n_439),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_463),
.B(n_466),
.Y(n_468)
);

OAI21xp33_ASAP7_75t_L g465 ( 
.A1(n_451),
.A2(n_4),
.B(n_7),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_450),
.B(n_4),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_464),
.A2(n_13),
.B(n_7),
.Y(n_467)
);

AOI21x1_ASAP7_75t_L g474 ( 
.A1(n_467),
.A2(n_1),
.B(n_2),
.Y(n_474)
);

A2O1A1O1Ixp25_ASAP7_75t_L g470 ( 
.A1(n_460),
.A2(n_461),
.B(n_7),
.C(n_11),
.D(n_13),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g472 ( 
.A(n_470),
.B(n_0),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_464),
.B(n_7),
.C(n_1),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_471),
.B(n_0),
.C(n_1),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_472),
.A2(n_469),
.B(n_468),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_473),
.B(n_474),
.Y(n_476)
);

BUFx24_ASAP7_75t_SL g477 ( 
.A(n_475),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_477),
.B(n_476),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_478),
.B(n_2),
.Y(n_479)
);

BUFx24_ASAP7_75t_SL g480 ( 
.A(n_479),
.Y(n_480)
);


endmodule