module fake_netlist_1_2488_n_704 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_704);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_704;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_27), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_45), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_43), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_72), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_13), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_17), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_61), .Y(n_85) );
BUFx3_ASAP7_75t_L g86 ( .A(n_12), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_59), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_75), .Y(n_88) );
BUFx2_ASAP7_75t_SL g89 ( .A(n_23), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_54), .Y(n_90) );
INVx1_ASAP7_75t_SL g91 ( .A(n_55), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_73), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_78), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_46), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_22), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_40), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_38), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_57), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_53), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_66), .Y(n_100) );
CKINVDCx14_ASAP7_75t_R g101 ( .A(n_8), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_52), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_10), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_58), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_28), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_31), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_26), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_15), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_39), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_49), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_77), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_20), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_70), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_24), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_5), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_69), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_11), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_47), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_8), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_48), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_29), .Y(n_124) );
OR2x2_ASAP7_75t_L g125 ( .A(n_32), .B(n_17), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_68), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_87), .Y(n_127) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_79), .A2(n_33), .B(n_74), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_105), .B(n_103), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_86), .B(n_0), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_114), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
NOR2x1_ASAP7_75t_L g139 ( .A(n_86), .B(n_0), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_88), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_90), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_103), .B(n_1), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_93), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_113), .B(n_2), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_117), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_107), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_96), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_97), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_113), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_97), .Y(n_155) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_98), .A2(n_34), .B(n_71), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_117), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_126), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_98), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_99), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_126), .B(n_3), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_107), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_101), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_107), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_82), .B(n_3), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_99), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_107), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_115), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_115), .Y(n_169) );
INVx2_ASAP7_75t_SL g170 ( .A(n_163), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_161), .B(n_83), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_163), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_130), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_147), .Y(n_174) );
BUFx10_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_130), .A2(n_120), .B1(n_84), .B2(n_112), .Y(n_176) );
OR2x6_ASAP7_75t_L g177 ( .A(n_147), .B(n_89), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_161), .B(n_108), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_154), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_161), .B(n_168), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_127), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_154), .B(n_100), .Y(n_182) );
OR2x2_ASAP7_75t_L g183 ( .A(n_143), .B(n_109), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_147), .A2(n_119), .B1(n_84), .B2(n_112), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_161), .A2(n_109), .B1(n_118), .B2(n_125), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_161), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_129), .B(n_104), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_129), .B(n_106), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_136), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_136), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_131), .B(n_92), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_168), .B(n_111), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_131), .B(n_118), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_133), .B(n_124), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_133), .B(n_102), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_168), .B(n_123), .Y(n_198) );
INVx4_ASAP7_75t_L g199 ( .A(n_136), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_169), .A2(n_125), .B1(n_89), .B2(n_121), .Y(n_200) );
NAND2xp33_ASAP7_75t_SL g201 ( .A(n_134), .B(n_110), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_168), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_134), .B(n_110), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_169), .B(n_95), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_135), .B(n_95), .Y(n_205) );
INVx5_ASAP7_75t_L g206 ( .A(n_127), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_166), .Y(n_207) );
INVx5_ASAP7_75t_L g208 ( .A(n_127), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_166), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_169), .B(n_91), .Y(n_210) );
INVxp33_ASAP7_75t_L g211 ( .A(n_143), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_166), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_135), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_127), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_127), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_127), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_138), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_138), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_140), .B(n_116), .Y(n_219) );
OAI22xp5_ASAP7_75t_SL g220 ( .A1(n_139), .A2(n_122), .B1(n_165), .B2(n_145), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_140), .A2(n_94), .B1(n_80), .B2(n_6), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_128), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_141), .B(n_155), .Y(n_223) );
OR2x2_ASAP7_75t_L g224 ( .A(n_141), .B(n_4), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_144), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_127), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_144), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_145), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_164), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_146), .B(n_4), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_146), .B(n_35), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_132), .Y(n_232) );
BUFx10_ASAP7_75t_L g233 ( .A(n_151), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_233), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_233), .Y(n_235) );
NAND2xp33_ASAP7_75t_L g236 ( .A(n_179), .B(n_152), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_211), .B(n_152), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_233), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_211), .B(n_153), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_173), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_189), .B(n_153), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_224), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_193), .B(n_151), .Y(n_243) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_180), .A2(n_155), .B(n_160), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_195), .B(n_159), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_185), .A2(n_159), .B1(n_160), .B2(n_139), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_172), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_176), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_203), .B(n_157), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_205), .B(n_157), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_175), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_225), .B(n_157), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_175), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_177), .A2(n_149), .B1(n_132), .B2(n_137), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_232), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_174), .B(n_149), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_183), .B(n_149), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_171), .B(n_132), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_182), .B(n_137), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_199), .B(n_137), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_232), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_182), .B(n_148), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_171), .B(n_148), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_202), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_214), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_171), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_204), .B(n_213), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_204), .B(n_148), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_214), .Y(n_269) );
INVxp67_ASAP7_75t_L g270 ( .A(n_170), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_217), .B(n_158), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_219), .B(n_158), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_184), .B(n_158), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_218), .B(n_156), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_227), .B(n_156), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_199), .B(n_167), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_186), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_228), .B(n_156), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_188), .B(n_167), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_207), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_177), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_219), .B(n_156), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_200), .B(n_156), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_180), .B(n_128), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_178), .A2(n_142), .B(n_150), .C(n_162), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_177), .B(n_128), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_187), .B(n_128), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_209), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_187), .B(n_128), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_196), .B(n_162), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_196), .B(n_162), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_197), .B(n_162), .Y(n_292) );
OAI22xp5_ASAP7_75t_SL g293 ( .A1(n_220), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_212), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_230), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_201), .A2(n_150), .B1(n_142), .B2(n_167), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_197), .B(n_150), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_192), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_192), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_178), .B(n_150), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_240), .B(n_190), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_298), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g303 ( .A1(n_246), .A2(n_223), .B(n_191), .C(n_210), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_286), .A2(n_222), .B(n_223), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_235), .B(n_210), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_266), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_235), .B(n_221), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_237), .B(n_198), .Y(n_308) );
NOR2xp33_ASAP7_75t_R g309 ( .A(n_247), .B(n_248), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_247), .Y(n_310) );
AO32x1_ASAP7_75t_L g311 ( .A1(n_287), .A2(n_222), .A3(n_181), .B1(n_226), .B2(n_216), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_241), .A2(n_194), .B(n_198), .C(n_231), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_248), .A2(n_194), .B1(n_231), .B2(n_142), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_236), .A2(n_142), .B1(n_226), .B2(n_216), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_284), .A2(n_215), .B(n_181), .Y(n_315) );
OR2x6_ASAP7_75t_L g316 ( .A(n_281), .B(n_164), .Y(n_316) );
AOI21x1_ASAP7_75t_L g317 ( .A1(n_283), .A2(n_215), .B(n_229), .Y(n_317) );
OA22x2_ASAP7_75t_L g318 ( .A1(n_293), .A2(n_7), .B1(n_9), .B2(n_10), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_245), .B(n_206), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_245), .B(n_206), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_270), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_274), .A2(n_229), .B(n_208), .Y(n_322) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_235), .B(n_208), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_299), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_242), .B(n_9), .Y(n_325) );
INVx4_ASAP7_75t_L g326 ( .A(n_235), .Y(n_326) );
INVx3_ASAP7_75t_SL g327 ( .A(n_251), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_234), .B(n_208), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_273), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_275), .A2(n_208), .B(n_206), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_278), .A2(n_206), .B(n_167), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_239), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_295), .B(n_11), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_289), .A2(n_167), .B(n_164), .Y(n_334) );
NOR3xp33_ASAP7_75t_SL g335 ( .A(n_257), .B(n_243), .C(n_272), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_264), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_236), .B(n_12), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_238), .B(n_13), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_252), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_251), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_276), .A2(n_167), .B(n_164), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_276), .A2(n_167), .B(n_164), .Y(n_342) );
NAND3xp33_ASAP7_75t_SL g343 ( .A(n_254), .B(n_14), .C(n_16), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_253), .B(n_164), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_253), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_280), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_277), .B(n_14), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g349 ( .A1(n_258), .A2(n_164), .B1(n_16), .B2(n_19), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_294), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_272), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_244), .B(n_18), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_SL g353 ( .A1(n_352), .A2(n_282), .B(n_268), .C(n_249), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_329), .A2(n_263), .B1(n_258), .B2(n_267), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_310), .Y(n_355) );
AOI21xp5_ASAP7_75t_SL g356 ( .A1(n_316), .A2(n_282), .B(n_263), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_335), .A2(n_250), .B(n_262), .C(n_259), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_327), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_321), .B(n_260), .Y(n_359) );
INVxp67_ASAP7_75t_L g360 ( .A(n_325), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_325), .Y(n_361) );
AO31x2_ASAP7_75t_L g362 ( .A1(n_352), .A2(n_271), .A3(n_297), .B(n_292), .Y(n_362) );
AO31x2_ASAP7_75t_L g363 ( .A1(n_334), .A2(n_291), .A3(n_290), .B(n_255), .Y(n_363) );
O2A1O1Ixp33_ASAP7_75t_L g364 ( .A1(n_333), .A2(n_256), .B(n_260), .C(n_300), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_332), .A2(n_339), .B1(n_351), .B2(n_346), .Y(n_365) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_318), .A2(n_261), .B1(n_296), .B2(n_256), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_304), .A2(n_279), .B(n_269), .Y(n_367) );
INVx4_ASAP7_75t_L g368 ( .A(n_326), .Y(n_368) );
A2O1A1Ixp33_ASAP7_75t_L g369 ( .A1(n_303), .A2(n_285), .B(n_279), .C(n_269), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_346), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_SL g371 ( .A1(n_307), .A2(n_265), .B(n_244), .C(n_30), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_333), .A2(n_265), .B1(n_25), .B2(n_36), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_337), .A2(n_21), .B1(n_37), .B2(n_41), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_L g374 ( .A1(n_343), .A2(n_42), .B(n_44), .C(n_50), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_301), .B(n_76), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_348), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g377 ( .A1(n_347), .A2(n_51), .B(n_56), .C(n_60), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_301), .B(n_62), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
O2A1O1Ixp5_ASAP7_75t_L g380 ( .A1(n_331), .A2(n_63), .B(n_64), .C(n_65), .Y(n_380) );
OR2x6_ASAP7_75t_L g381 ( .A(n_316), .B(n_67), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_336), .Y(n_382) );
NOR2xp67_ASAP7_75t_SL g383 ( .A(n_326), .B(n_345), .Y(n_383) );
AO31x2_ASAP7_75t_L g384 ( .A1(n_322), .A2(n_315), .A3(n_311), .B(n_341), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_340), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_355), .B(n_309), .Y(n_386) );
OA21x2_ASAP7_75t_L g387 ( .A1(n_380), .A2(n_317), .B(n_342), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_381), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g389 ( .A1(n_357), .A2(n_312), .B(n_320), .C(n_319), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_376), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_375), .B(n_306), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_361), .B(n_308), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_366), .B(n_349), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_353), .A2(n_311), .B(n_330), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_360), .B(n_318), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_371), .A2(n_311), .B(n_305), .Y(n_396) );
AO31x2_ASAP7_75t_L g397 ( .A1(n_372), .A2(n_338), .A3(n_324), .B(n_302), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_365), .B(n_345), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_367), .A2(n_319), .B(n_320), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_356), .A2(n_344), .B(n_328), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_358), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_354), .B(n_340), .Y(n_403) );
A2O1A1Ixp33_ASAP7_75t_L g404 ( .A1(n_374), .A2(n_313), .B(n_314), .C(n_340), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_369), .A2(n_316), .B(n_323), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_358), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_364), .A2(n_323), .B(n_345), .Y(n_407) );
OAI21xp5_ASAP7_75t_L g408 ( .A1(n_382), .A2(n_378), .B(n_359), .Y(n_408) );
OAI21x1_ASAP7_75t_L g409 ( .A1(n_373), .A2(n_384), .B(n_370), .Y(n_409) );
BUFx12f_ASAP7_75t_L g410 ( .A(n_368), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_375), .Y(n_411) );
OAI21x1_ASAP7_75t_L g412 ( .A1(n_384), .A2(n_363), .B(n_362), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_381), .A2(n_377), .B(n_362), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_412), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_389), .B(n_362), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_388), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_390), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_412), .Y(n_418) );
OR2x6_ASAP7_75t_L g419 ( .A(n_388), .B(n_381), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_409), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_402), .Y(n_421) );
OA21x2_ASAP7_75t_L g422 ( .A1(n_394), .A2(n_384), .B(n_363), .Y(n_422) );
NOR2xp67_ASAP7_75t_L g423 ( .A(n_388), .B(n_368), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_388), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_395), .B(n_363), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_389), .A2(n_383), .B1(n_385), .B2(n_392), .C(n_411), .Y(n_426) );
INVx3_ASAP7_75t_L g427 ( .A(n_410), .Y(n_427) );
AOI21xp5_ASAP7_75t_SL g428 ( .A1(n_391), .A2(n_413), .B(n_398), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_391), .B(n_386), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_410), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_403), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_409), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_399), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_401), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_387), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_391), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_393), .A2(n_408), .B1(n_401), .B2(n_406), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_397), .B(n_393), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_400), .Y(n_439) );
AO21x2_ASAP7_75t_L g440 ( .A1(n_396), .A2(n_405), .B(n_404), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_397), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_397), .B(n_404), .Y(n_442) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_407), .A2(n_397), .B(n_387), .Y(n_443) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_387), .A2(n_394), .B(n_396), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_388), .B(n_409), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_388), .B(n_412), .Y(n_446) );
OR2x6_ASAP7_75t_L g447 ( .A(n_388), .B(n_413), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_395), .A2(n_293), .B1(n_335), .B2(n_236), .C(n_357), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_412), .Y(n_449) );
OAI211xp5_ASAP7_75t_SL g450 ( .A1(n_448), .A2(n_429), .B(n_427), .C(n_421), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_425), .B(n_446), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_425), .B(n_431), .Y(n_452) );
INVx5_ASAP7_75t_SL g453 ( .A(n_419), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_425), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_430), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_417), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_441), .Y(n_457) );
NOR2xp33_ASAP7_75t_SL g458 ( .A(n_430), .B(n_427), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_419), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_441), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_431), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_427), .B(n_430), .Y(n_462) );
INVx5_ASAP7_75t_L g463 ( .A(n_419), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_427), .B(n_429), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_419), .Y(n_465) );
INVx5_ASAP7_75t_L g466 ( .A(n_419), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_434), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_446), .B(n_438), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_446), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_433), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_438), .B(n_421), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_424), .B(n_434), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_438), .B(n_417), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_414), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_433), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_436), .B(n_437), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_419), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_436), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_414), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_424), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_423), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_415), .B(n_437), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_442), .B(n_445), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_427), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_414), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_418), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_418), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_418), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_449), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_442), .B(n_445), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_442), .B(n_445), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_416), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_449), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_445), .B(n_422), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_445), .B(n_447), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_422), .B(n_415), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_448), .B(n_416), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_449), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_471), .B(n_439), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_452), .B(n_422), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_462), .B(n_428), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_456), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_451), .B(n_447), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_461), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_461), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_452), .B(n_422), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_471), .B(n_426), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_469), .B(n_447), .Y(n_510) );
BUFx3_ASAP7_75t_L g511 ( .A(n_485), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_473), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_473), .B(n_426), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_469), .B(n_447), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_451), .B(n_447), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_468), .B(n_447), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_468), .B(n_422), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_455), .B(n_432), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_481), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_479), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_464), .B(n_432), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_450), .B(n_458), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_457), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_457), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_454), .B(n_440), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_460), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_460), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_454), .B(n_440), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_483), .B(n_440), .Y(n_529) );
BUFx2_ASAP7_75t_L g530 ( .A(n_487), .Y(n_530) );
NAND3x1_ASAP7_75t_L g531 ( .A(n_496), .B(n_440), .C(n_444), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_484), .B(n_440), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_474), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_499), .A2(n_420), .B1(n_444), .B2(n_443), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_494), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_497), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_484), .B(n_420), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_483), .B(n_420), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_470), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_492), .B(n_435), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_467), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_497), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_497), .B(n_435), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_493), .B(n_476), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_498), .B(n_444), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_493), .B(n_443), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_470), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_475), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_475), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_498), .B(n_444), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_496), .B(n_443), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_482), .B(n_443), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_474), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_486), .B(n_443), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_486), .B(n_500), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_478), .B(n_463), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_472), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_485), .B(n_477), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_517), .B(n_459), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_523), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_517), .B(n_459), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_541), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_530), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_546), .B(n_465), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_535), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_533), .Y(n_566) );
INVx4_ASAP7_75t_L g567 ( .A(n_511), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_524), .Y(n_568) );
INVx4_ASAP7_75t_L g569 ( .A(n_511), .Y(n_569) );
NAND2x1_ASAP7_75t_L g570 ( .A(n_556), .B(n_465), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_557), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_501), .B(n_463), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_526), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_533), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_546), .B(n_488), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_551), .B(n_488), .Y(n_576) );
OAI22xp33_ASAP7_75t_SL g577 ( .A1(n_503), .A2(n_463), .B1(n_466), .B2(n_478), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_551), .B(n_500), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_540), .B(n_495), .Y(n_579) );
INVx3_ASAP7_75t_SL g580 ( .A(n_556), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_512), .B(n_472), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_544), .B(n_495), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_527), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_556), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_540), .B(n_491), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_544), .B(n_491), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_504), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_539), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_547), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_506), .B(n_453), .Y(n_590) );
INVx3_ASAP7_75t_L g591 ( .A(n_543), .Y(n_591) );
INVx4_ASAP7_75t_L g592 ( .A(n_543), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_507), .B(n_453), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_553), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_550), .B(n_480), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_555), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_548), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_532), .B(n_489), .Y(n_598) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_555), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_550), .B(n_490), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_522), .B(n_463), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_502), .B(n_453), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_553), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_519), .Y(n_604) );
NAND2xp33_ASAP7_75t_SL g605 ( .A(n_502), .B(n_453), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_520), .B(n_463), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_549), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_565), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_576), .B(n_528), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_596), .B(n_528), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_599), .B(n_525), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_571), .B(n_525), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_562), .B(n_545), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_587), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_604), .Y(n_615) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_601), .A2(n_552), .B(n_558), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_576), .B(n_537), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_563), .B(n_534), .C(n_518), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_575), .B(n_513), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_582), .Y(n_620) );
CKINVDCx16_ASAP7_75t_R g621 ( .A(n_567), .Y(n_621) );
INVx2_ASAP7_75t_SL g622 ( .A(n_580), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_582), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_586), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_575), .B(n_509), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_586), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_578), .B(n_508), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_567), .B(n_529), .C(n_521), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_560), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_578), .B(n_537), .Y(n_630) );
CKINVDCx16_ASAP7_75t_R g631 ( .A(n_567), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_560), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_595), .Y(n_633) );
INVxp67_ASAP7_75t_SL g634 ( .A(n_595), .Y(n_634) );
BUFx2_ASAP7_75t_L g635 ( .A(n_580), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_559), .B(n_516), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_559), .B(n_516), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_568), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_580), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_598), .B(n_508), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_572), .A2(n_510), .B1(n_514), .B2(n_515), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_568), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_573), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_606), .Y(n_644) );
AOI222xp33_ASAP7_75t_L g645 ( .A1(n_623), .A2(n_561), .B1(n_564), .B2(n_581), .C1(n_605), .C2(n_598), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_627), .Y(n_646) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_633), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_627), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_613), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_621), .A2(n_561), .B1(n_564), .B2(n_592), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_608), .A2(n_616), .B1(n_624), .B2(n_618), .C(n_644), .Y(n_651) );
OAI211xp5_ASAP7_75t_L g652 ( .A1(n_635), .A2(n_569), .B(n_570), .C(n_592), .Y(n_652) );
AOI221xp5_ASAP7_75t_SL g653 ( .A1(n_639), .A2(n_577), .B1(n_584), .B2(n_505), .C(n_515), .Y(n_653) );
OAI211xp5_ASAP7_75t_L g654 ( .A1(n_635), .A2(n_569), .B(n_570), .C(n_592), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_628), .A2(n_569), .B(n_602), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_633), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_609), .B(n_585), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_640), .B(n_585), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_619), .A2(n_583), .B1(n_597), .B2(n_589), .C(n_588), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_609), .B(n_579), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_629), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_632), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_622), .B(n_542), .Y(n_663) );
NAND2x1p5_ASAP7_75t_L g664 ( .A(n_622), .B(n_466), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_631), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_634), .A2(n_505), .B1(n_602), .B2(n_593), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_625), .B(n_536), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_665), .Y(n_668) );
OAI22xp5_ASAP7_75t_SL g669 ( .A1(n_650), .A2(n_641), .B1(n_466), .B2(n_626), .Y(n_669) );
OAI32xp33_ASAP7_75t_L g670 ( .A1(n_646), .A2(n_620), .A3(n_611), .B1(n_610), .B2(n_612), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_652), .A2(n_630), .B1(n_617), .B2(n_636), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_654), .A2(n_614), .B(n_615), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_648), .Y(n_673) );
OAI322xp33_ASAP7_75t_L g674 ( .A1(n_649), .A2(n_529), .A3(n_643), .B1(n_642), .B2(n_638), .C1(n_600), .C2(n_607), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_SL g675 ( .A1(n_647), .A2(n_591), .B(n_590), .C(n_600), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_655), .A2(n_531), .B(n_630), .Y(n_676) );
BUFx2_ASAP7_75t_L g677 ( .A(n_663), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g678 ( .A1(n_666), .A2(n_466), .B1(n_591), .B2(n_542), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_651), .B(n_617), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_653), .A2(n_637), .B(n_636), .C(n_591), .Y(n_680) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_645), .A2(n_573), .B(n_589), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_679), .B(n_659), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_676), .A2(n_656), .B(n_662), .Y(n_683) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_671), .A2(n_664), .B(n_666), .Y(n_684) );
NAND4xp25_ASAP7_75t_L g685 ( .A(n_681), .B(n_663), .C(n_667), .D(n_536), .Y(n_685) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_677), .B(n_661), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_673), .Y(n_687) );
NOR2x1_ASAP7_75t_SL g688 ( .A(n_675), .B(n_658), .Y(n_688) );
OAI211xp5_ASAP7_75t_L g689 ( .A1(n_668), .A2(n_466), .B(n_660), .C(n_657), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_682), .A2(n_670), .B1(n_674), .B2(n_672), .C(n_669), .Y(n_690) );
NOR5xp2_ASAP7_75t_L g691 ( .A(n_684), .B(n_680), .C(n_678), .D(n_583), .E(n_607), .Y(n_691) );
NOR2x1_ASAP7_75t_L g692 ( .A(n_686), .B(n_678), .Y(n_692) );
NOR5xp2_ASAP7_75t_L g693 ( .A(n_683), .B(n_597), .C(n_588), .D(n_531), .E(n_637), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_692), .B(n_688), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_690), .B(n_685), .C(n_689), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_691), .B(n_687), .C(n_542), .Y(n_696) );
AO22x2_ASAP7_75t_L g697 ( .A1(n_694), .A2(n_693), .B1(n_536), .B2(n_574), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_696), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_698), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_699), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_695), .B(n_697), .Y(n_701) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_701), .A2(n_697), .B(n_554), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_702), .A2(n_538), .B1(n_603), .B2(n_574), .Y(n_703) );
AOI222xp33_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_603), .B1(n_594), .B2(n_566), .C1(n_554), .C2(n_579), .Y(n_704) );
endmodule