module fake_aes_6850_n_14 (n_1, n_2, n_4, n_3, n_0, n_14);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
AO21x2_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_4), .B(n_0), .Y(n_5) );
CKINVDCx5p33_ASAP7_75t_R g6 ( .A(n_1), .Y(n_6) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_6), .B(n_2), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
INVx1_ASAP7_75t_SL g9 ( .A(n_8), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_9), .B(n_5), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
INVxp67_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
INVx1_ASAP7_75t_SL g14 ( .A(n_13), .Y(n_14) );
endmodule