module fake_ariane_3132_n_1342 (n_295, n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_289, n_288, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_294, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_274, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_281, n_209, n_49, n_262, n_291, n_20, n_292, n_174, n_275, n_100, n_17, n_283, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_290, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_286, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_287, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_284, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_278, n_122, n_268, n_257, n_266, n_198, n_282, n_148, n_232, n_164, n_52, n_277, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_293, n_171, n_228, n_15, n_118, n_93, n_121, n_276, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_279, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_280, n_215, n_252, n_142, n_251, n_161, n_285, n_14, n_163, n_88, n_186, n_141, n_296, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_273, n_54, n_25, n_1342);

input n_295;
input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_289;
input n_288;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_294;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_274;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_281;
input n_209;
input n_49;
input n_262;
input n_291;
input n_20;
input n_292;
input n_174;
input n_275;
input n_100;
input n_17;
input n_283;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_290;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_286;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_287;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_284;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_278;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_282;
input n_148;
input n_232;
input n_164;
input n_52;
input n_277;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_293;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_276;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_279;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_280;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_285;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_296;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_273;
input n_54;
input n_25;

output n_1342;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_302;
wire n_380;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_337;
wire n_967;
wire n_1083;
wire n_746;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1266;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1341;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_203),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_26),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_119),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_142),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_296),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_218),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_292),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_288),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_58),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_242),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_22),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_75),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_117),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_32),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_267),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_109),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_85),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_183),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_243),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_17),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_233),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_144),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_27),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_206),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_134),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_3),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_257),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_285),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_89),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_132),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_232),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_95),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_215),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_237),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_143),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_157),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_275),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_253),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_64),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_115),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_26),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_55),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_208),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_163),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_216),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_29),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_147),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_295),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_169),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_214),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_140),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_235),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_190),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_256),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_236),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_27),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_234),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_164),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_80),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_84),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_239),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g364 ( 
.A(n_213),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_200),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_230),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_284),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_228),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_217),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_15),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_241),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_137),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_248),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_196),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_50),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_34),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_88),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_219),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_171),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_197),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_165),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_258),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_61),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_192),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_199),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_153),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_4),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_87),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_62),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_126),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_6),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_286),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_53),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_210),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_67),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_123),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_91),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_90),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_112),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_73),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_120),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_6),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_201),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_191),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_231),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_152),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_162),
.Y(n_407)
);

BUFx8_ASAP7_75t_SL g408 ( 
.A(n_150),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_46),
.B(n_250),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_76),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_57),
.B(n_125),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_39),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_254),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_269),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_82),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_175),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_44),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_68),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_34),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_16),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_98),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_240),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_225),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_97),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_15),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_9),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_266),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_50),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_13),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_0),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_265),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_178),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_23),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_22),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_207),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_223),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_283),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_246),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_179),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_259),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_37),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_110),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_11),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_146),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_280),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_124),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_184),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_77),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_8),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_211),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_122),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_291),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_187),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_31),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_72),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_202),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_205),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_224),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_36),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_29),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_39),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_244),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_114),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_263),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_145),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_1),
.B(n_281),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_116),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_103),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_138),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_108),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_161),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_238),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_226),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_245),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_31),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_10),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_7),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_59),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_273),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_194),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_209),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_289),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_227),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_222),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_156),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_9),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_133),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_1),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_180),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_130),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_12),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_141),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_188),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_65),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_182),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_189),
.Y(n_496)
);

BUFx10_ASAP7_75t_L g497 ( 
.A(n_270),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_3),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_185),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_35),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_118),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_274),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_28),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_252),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_21),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_177),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_293),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_271),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_264),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_92),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_52),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_5),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_2),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_186),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_46),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_212),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_13),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_131),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_96),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_94),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_204),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_86),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_44),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_0),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_370),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_488),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_488),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_368),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_408),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_368),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_470),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_312),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_312),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_428),
.B(n_7),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_340),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_391),
.Y(n_536)
);

BUFx12f_ASAP7_75t_L g537 ( 
.A(n_320),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_470),
.Y(n_538)
);

AOI22x1_ASAP7_75t_SL g539 ( 
.A1(n_376),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

OA21x2_ASAP7_75t_L g541 ( 
.A1(n_299),
.A2(n_14),
.B(n_16),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_398),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_523),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_391),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_298),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_322),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_404),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_425),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_425),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_348),
.B(n_14),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_404),
.Y(n_551)
);

INVx6_ASAP7_75t_L g552 ( 
.A(n_320),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_306),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_302),
.A2(n_17),
.B(n_18),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_306),
.A2(n_56),
.B(n_54),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_463),
.Y(n_556)
);

BUFx8_ASAP7_75t_SL g557 ( 
.A(n_387),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_470),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_323),
.B(n_60),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_507),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_330),
.Y(n_561)
);

OA21x2_ASAP7_75t_L g562 ( 
.A1(n_309),
.A2(n_18),
.B(n_19),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_427),
.B(n_19),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_323),
.B(n_385),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_507),
.Y(n_565)
);

OAI21x1_ASAP7_75t_L g566 ( 
.A1(n_385),
.A2(n_66),
.B(n_63),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_524),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_403),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_409),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_503),
.B(n_20),
.Y(n_570)
);

OA21x2_ASAP7_75t_L g571 ( 
.A1(n_310),
.A2(n_24),
.B(n_25),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_330),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_403),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_343),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_311),
.B(n_24),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_463),
.B(n_25),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_325),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_319),
.B(n_28),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_358),
.B(n_30),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_507),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_412),
.B(n_419),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_343),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_507),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_410),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_383),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_426),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_449),
.B(n_30),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_313),
.B(n_32),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_459),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_432),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_383),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_473),
.Y(n_592)
);

AND2x2_ASAP7_75t_SL g593 ( 
.A(n_466),
.B(n_33),
.Y(n_593)
);

BUFx12f_ASAP7_75t_L g594 ( 
.A(n_473),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_315),
.B(n_33),
.Y(n_595)
);

BUFx8_ASAP7_75t_SL g596 ( 
.A(n_483),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_432),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_461),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_318),
.B(n_35),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_497),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_522),
.B(n_36),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_462),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_477),
.B(n_37),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_462),
.Y(n_604)
);

BUFx8_ASAP7_75t_SL g605 ( 
.A(n_341),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_321),
.B(n_324),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_497),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_342),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_512),
.B(n_38),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_373),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_307),
.B(n_38),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_508),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_515),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_508),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_326),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_347),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_375),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_333),
.Y(n_619)
);

AOI22x1_ASAP7_75t_SL g620 ( 
.A1(n_430),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_334),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_335),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_510),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_402),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_517),
.B(n_40),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_417),
.B(n_41),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_510),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_345),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_346),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_349),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_350),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_420),
.B(n_42),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_351),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_429),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_354),
.B(n_357),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_365),
.Y(n_636)
);

OA21x2_ASAP7_75t_L g637 ( 
.A1(n_371),
.A2(n_43),
.B(n_45),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_372),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_433),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_374),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_434),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_297),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_382),
.Y(n_643)
);

OA21x2_ASAP7_75t_L g644 ( 
.A1(n_400),
.A2(n_43),
.B(n_45),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_441),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_423),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_435),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_443),
.Y(n_648)
);

OA21x2_ASAP7_75t_L g649 ( 
.A1(n_436),
.A2(n_47),
.B(n_48),
.Y(n_649)
);

BUFx12f_ASAP7_75t_L g650 ( 
.A(n_454),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_437),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_300),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_438),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_440),
.B(n_47),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_460),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_475),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_369),
.B(n_69),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_448),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_476),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_453),
.Y(n_660)
);

OAI22x1_ASAP7_75t_R g661 ( 
.A1(n_486),
.A2(n_49),
.B1(n_51),
.B2(n_70),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_458),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_465),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_467),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_378),
.B(n_71),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_469),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_472),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_474),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_479),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_491),
.B(n_498),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_500),
.Y(n_671)
);

BUFx12f_ASAP7_75t_L g672 ( 
.A(n_505),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_480),
.B(n_74),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_485),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_487),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_490),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_513),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_499),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_501),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_596),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_526),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_565),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_535),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_584),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_529),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_605),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_557),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_531),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_584),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_584),
.Y(n_690)
);

XOR2xp5_ASAP7_75t_L g691 ( 
.A(n_618),
.B(n_301),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_531),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_597),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_642),
.B(n_317),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_574),
.B(n_600),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g696 ( 
.A(n_606),
.B(n_506),
.C(n_502),
.Y(n_696)
);

AND2x6_ASAP7_75t_L g697 ( 
.A(n_550),
.B(n_509),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_R g698 ( 
.A(n_645),
.B(n_303),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_597),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_597),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_624),
.Y(n_701)
);

AO21x2_ASAP7_75t_L g702 ( 
.A1(n_575),
.A2(n_514),
.B(n_511),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_528),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_543),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_565),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_531),
.Y(n_706)
);

CKINVDCx16_ASAP7_75t_R g707 ( 
.A(n_537),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_574),
.B(n_411),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_642),
.B(n_652),
.Y(n_709)
);

XNOR2xp5_ASAP7_75t_L g710 ( 
.A(n_593),
.B(n_337),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_671),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_552),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_639),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_650),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_672),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_546),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_577),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_538),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_594),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_552),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_R g721 ( 
.A(n_545),
.B(n_304),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_538),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_652),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_574),
.B(n_519),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_602),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_572),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_617),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_602),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_R g729 ( 
.A(n_641),
.B(n_521),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_R g730 ( 
.A(n_641),
.B(n_305),
.Y(n_730)
);

NOR2x1p5_ASAP7_75t_L g731 ( 
.A(n_585),
.B(n_308),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_582),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_592),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_602),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_604),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_607),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_538),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_677),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_604),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_600),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_540),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_600),
.Y(n_742)
);

NOR2xp67_ASAP7_75t_L g743 ( 
.A(n_591),
.B(n_464),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_634),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_655),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_659),
.Y(n_746)
);

AND3x2_ASAP7_75t_L g747 ( 
.A(n_534),
.B(n_384),
.C(n_355),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_670),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_604),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_613),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_R g751 ( 
.A(n_648),
.B(n_314),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_561),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_616),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_R g754 ( 
.A(n_648),
.B(n_520),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_621),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_540),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_591),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_638),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_R g759 ( 
.A(n_550),
.B(n_316),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_613),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_608),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_527),
.B(n_397),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_R g763 ( 
.A(n_628),
.B(n_327),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_530),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_R g765 ( 
.A(n_628),
.B(n_518),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_SL g766 ( 
.A1(n_569),
.A2(n_525),
.B1(n_656),
.B2(n_661),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_613),
.Y(n_767)
);

CKINVDCx16_ASAP7_75t_R g768 ( 
.A(n_661),
.Y(n_768)
);

AOI21x1_ASAP7_75t_L g769 ( 
.A1(n_553),
.A2(n_364),
.B(n_329),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_608),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_R g771 ( 
.A(n_563),
.B(n_328),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_608),
.B(n_401),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_540),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_610),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_615),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_542),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_630),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_615),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_615),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_R g780 ( 
.A(n_640),
.B(n_516),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_610),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_716),
.B(n_717),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_712),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_748),
.B(n_563),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_777),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_682),
.B(n_576),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_748),
.B(n_709),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_777),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_764),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_703),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_L g791 ( 
.A(n_766),
.B(n_569),
.C(n_656),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_681),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_698),
.B(n_570),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_684),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_682),
.B(n_610),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_689),
.Y(n_796)
);

BUFx5_ASAP7_75t_L g797 ( 
.A(n_697),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_688),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_705),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_776),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_688),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_705),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_716),
.B(n_547),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_762),
.B(n_612),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_723),
.B(n_612),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_690),
.Y(n_806)
);

AO221x1_ASAP7_75t_L g807 ( 
.A1(n_717),
.A2(n_620),
.B1(n_539),
.B2(n_525),
.C(n_640),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_753),
.B(n_570),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_691),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_693),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_699),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_694),
.B(n_755),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_758),
.B(n_551),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_700),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_697),
.B(n_556),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_688),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_732),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_725),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_768),
.B(n_595),
.C(n_575),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_728),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_772),
.B(n_663),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_763),
.B(n_611),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_721),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_765),
.B(n_780),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_724),
.B(n_664),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_733),
.B(n_664),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_741),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_SL g828 ( 
.A(n_711),
.B(n_625),
.Y(n_828)
);

BUFx5_ASAP7_75t_L g829 ( 
.A(n_697),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_734),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_685),
.B(n_619),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_736),
.B(n_635),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_727),
.B(n_626),
.Y(n_833)
);

OR2x6_ASAP7_75t_L g834 ( 
.A(n_695),
.B(n_586),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_697),
.B(n_622),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_735),
.Y(n_836)
);

OR2x6_ASAP7_75t_L g837 ( 
.A(n_731),
.B(n_589),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_702),
.B(n_629),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_739),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_740),
.B(n_632),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_738),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_708),
.B(n_647),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_729),
.B(n_578),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_749),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_750),
.Y(n_845)
);

BUFx6f_ASAP7_75t_SL g846 ( 
.A(n_686),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_759),
.B(n_601),
.C(n_588),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_742),
.B(n_653),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_744),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_760),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_696),
.B(n_658),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_761),
.B(n_660),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_L g853 ( 
.A(n_730),
.B(n_595),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_745),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_751),
.B(n_754),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_746),
.B(n_599),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_720),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_726),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_743),
.B(n_662),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_770),
.B(n_578),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_767),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_774),
.B(n_579),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_775),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_778),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_779),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_781),
.B(n_667),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_771),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_747),
.B(n_668),
.Y(n_868)
);

BUFx5_ASAP7_75t_L g869 ( 
.A(n_769),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_710),
.B(n_669),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_757),
.B(n_630),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_713),
.B(n_579),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_692),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_706),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_718),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_722),
.B(n_623),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_787),
.B(n_587),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_821),
.B(n_587),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_792),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_802),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_846),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_806),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_818),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_785),
.Y(n_884)
);

NOR3xp33_ASAP7_75t_SL g885 ( 
.A(n_784),
.B(n_654),
.C(n_687),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_858),
.Y(n_886)
);

BUFx8_ASAP7_75t_L g887 ( 
.A(n_841),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_826),
.B(n_714),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_788),
.Y(n_889)
);

INVx4_ASAP7_75t_L g890 ( 
.A(n_797),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_812),
.B(n_603),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_782),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_SL g893 ( 
.A(n_817),
.B(n_704),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_849),
.B(n_707),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_823),
.B(n_752),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_786),
.A2(n_673),
.B(n_599),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_783),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_847),
.A2(n_564),
.B1(n_609),
.B2(n_603),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_854),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_820),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_795),
.A2(n_566),
.B(n_555),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_832),
.B(n_609),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_857),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_867),
.B(n_715),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_825),
.B(n_631),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_830),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_834),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_803),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_809),
.B(n_683),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_793),
.B(n_701),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_790),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_791),
.A2(n_564),
.B1(n_623),
.B2(n_631),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_L g913 ( 
.A(n_870),
.B(n_719),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_837),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_794),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_831),
.B(n_631),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_851),
.B(n_633),
.Y(n_917)
);

AND2x6_ASAP7_75t_L g918 ( 
.A(n_835),
.B(n_581),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_861),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_863),
.Y(n_920)
);

NOR2x1_ASAP7_75t_L g921 ( 
.A(n_855),
.B(n_457),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_871),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_853),
.A2(n_856),
.B1(n_833),
.B2(n_843),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_828),
.A2(n_564),
.B1(n_332),
.B2(n_336),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_865),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_796),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_SL g927 ( 
.A(n_819),
.B(n_680),
.C(n_539),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_L g928 ( 
.A(n_824),
.B(n_620),
.C(n_633),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_813),
.B(n_536),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_799),
.B(n_840),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_808),
.B(n_636),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_876),
.Y(n_932)
);

INVxp67_ASAP7_75t_SL g933 ( 
.A(n_797),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_810),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_811),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_789),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_814),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_838),
.A2(n_564),
.B1(n_623),
.B2(n_636),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_836),
.Y(n_939)
);

INVx5_ASAP7_75t_L g940 ( 
.A(n_834),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_800),
.B(n_544),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_797),
.B(n_636),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_839),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_845),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_850),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_798),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_868),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_798),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_822),
.A2(n_338),
.B1(n_339),
.B2(n_331),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_864),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_860),
.B(n_598),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_799),
.B(n_643),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_872),
.B(n_614),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_804),
.A2(n_554),
.B(n_541),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_862),
.A2(n_562),
.B1(n_571),
.B2(n_541),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_798),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_805),
.B(n_848),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_873),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_801),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_807),
.A2(n_646),
.B1(n_651),
.B2(n_643),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_874),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_797),
.A2(n_352),
.B1(n_353),
.B2(n_344),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_875),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_852),
.B(n_544),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_844),
.B(n_643),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_829),
.A2(n_359),
.B1(n_360),
.B2(n_356),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_801),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_815),
.A2(n_651),
.B1(n_666),
.B2(n_646),
.Y(n_968)
);

XOR2xp5_ASAP7_75t_L g969 ( 
.A(n_866),
.B(n_646),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_859),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_842),
.B(n_651),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_829),
.B(n_666),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_829),
.B(n_674),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_SL g974 ( 
.A(n_869),
.B(n_362),
.C(n_361),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_SL g975 ( 
.A1(n_928),
.A2(n_571),
.B1(n_637),
.B2(n_562),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_952),
.A2(n_930),
.B(n_896),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_882),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_901),
.A2(n_644),
.B(n_637),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_923),
.A2(n_877),
.B(n_902),
.C(n_891),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_878),
.A2(n_869),
.B(n_649),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_892),
.A2(n_568),
.B(n_573),
.C(n_553),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_903),
.Y(n_982)
);

O2A1O1Ixp5_ASAP7_75t_L g983 ( 
.A1(n_957),
.A2(n_756),
.B(n_773),
.C(n_737),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_880),
.A2(n_573),
.B(n_590),
.C(n_568),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_940),
.B(n_567),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_886),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_909),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_922),
.B(n_674),
.Y(n_988)
);

AO32x2_ASAP7_75t_L g989 ( 
.A1(n_955),
.A2(n_869),
.A3(n_644),
.B1(n_649),
.B2(n_678),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_SL g990 ( 
.A1(n_931),
.A2(n_533),
.B(n_548),
.C(n_532),
.Y(n_990)
);

BUFx8_ASAP7_75t_SL g991 ( 
.A(n_881),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_898),
.A2(n_366),
.B1(n_367),
.B2(n_363),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_887),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_909),
.B(n_532),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_899),
.A2(n_377),
.B1(n_380),
.B2(n_379),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_R g996 ( 
.A(n_893),
.B(n_801),
.Y(n_996)
);

OR2x6_ASAP7_75t_L g997 ( 
.A(n_907),
.B(n_533),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_897),
.B(n_940),
.Y(n_998)
);

AOI22x1_ASAP7_75t_L g999 ( 
.A1(n_932),
.A2(n_954),
.B1(n_933),
.B2(n_883),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_936),
.A2(n_627),
.B(n_549),
.C(n_567),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_972),
.A2(n_869),
.B(n_386),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_895),
.B(n_816),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_929),
.B(n_674),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_964),
.B(n_675),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_900),
.A2(n_549),
.B(n_676),
.C(n_675),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_924),
.B(n_827),
.Y(n_1006)
);

BUFx4f_ASAP7_75t_L g1007 ( 
.A(n_894),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_905),
.A2(n_388),
.B(n_381),
.Y(n_1008)
);

AOI22x1_ASAP7_75t_L g1009 ( 
.A1(n_906),
.A2(n_827),
.B1(n_816),
.B2(n_676),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_890),
.A2(n_390),
.B(n_389),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_910),
.A2(n_452),
.B1(n_392),
.B2(n_393),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_890),
.A2(n_456),
.B1(n_394),
.B2(n_395),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_L g1013 ( 
.A(n_888),
.B(n_399),
.C(n_396),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_919),
.A2(n_481),
.B1(n_405),
.B2(n_406),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_911),
.B(n_908),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_913),
.B(n_816),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_970),
.B(n_675),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_887),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_960),
.A2(n_879),
.B1(n_925),
.B2(n_920),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_962),
.A2(n_478),
.B1(n_407),
.B2(n_431),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_915),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_934),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_969),
.B(n_676),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_914),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_951),
.A2(n_679),
.B1(n_678),
.B2(n_559),
.Y(n_1025)
);

NAND3xp33_ASAP7_75t_SL g1026 ( 
.A(n_885),
.B(n_414),
.C(n_413),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_941),
.A2(n_679),
.B(n_415),
.C(n_484),
.Y(n_1027)
);

BUFx10_ASAP7_75t_L g1028 ( 
.A(n_951),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_973),
.A2(n_418),
.B(n_416),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_949),
.B(n_827),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_937),
.A2(n_679),
.B1(n_559),
.B2(n_665),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_946),
.Y(n_1032)
);

NAND2xp33_ASAP7_75t_SL g1033 ( 
.A(n_974),
.B(n_421),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_942),
.A2(n_424),
.B(n_422),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_939),
.A2(n_559),
.B1(n_665),
.B2(n_657),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_917),
.B(n_559),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_904),
.B(n_439),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_943),
.A2(n_657),
.B1(n_665),
.B2(n_492),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_947),
.B(n_657),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_953),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_944),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_912),
.B(n_657),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_971),
.B(n_665),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_918),
.B(n_442),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_L g1045 ( 
.A(n_921),
.B(n_741),
.Y(n_1045)
);

NOR2xp67_ASAP7_75t_L g1046 ( 
.A(n_961),
.B(n_444),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_967),
.A2(n_446),
.B(n_445),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_884),
.B(n_447),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_945),
.B(n_450),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_965),
.A2(n_468),
.B(n_451),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_889),
.A2(n_495),
.B(n_471),
.C(n_482),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_950),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_966),
.A2(n_504),
.B1(n_489),
.B2(n_493),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_918),
.B(n_494),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_1032),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_1032),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_999),
.A2(n_963),
.B(n_935),
.Y(n_1057)
);

AO21x2_ASAP7_75t_L g1058 ( 
.A1(n_978),
.A2(n_980),
.B(n_1001),
.Y(n_1058)
);

BUFx2_ASAP7_75t_SL g1059 ( 
.A(n_993),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_991),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_979),
.A2(n_938),
.B1(n_926),
.B2(n_959),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_994),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_982),
.Y(n_1063)
);

OR2x6_ASAP7_75t_L g1064 ( 
.A(n_994),
.B(n_916),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_977),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_976),
.A2(n_958),
.B(n_968),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1022),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_983),
.A2(n_1009),
.B(n_1036),
.Y(n_1068)
);

INVx5_ASAP7_75t_L g1069 ( 
.A(n_987),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1006),
.A2(n_948),
.B(n_946),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1002),
.B(n_948),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_1016),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_986),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_1018),
.B(n_948),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_1028),
.Y(n_1075)
);

AO21x2_ASAP7_75t_L g1076 ( 
.A1(n_1043),
.A2(n_927),
.B(n_956),
.Y(n_1076)
);

BUFx5_ASAP7_75t_L g1077 ( 
.A(n_1041),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1021),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1052),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_988),
.B(n_1019),
.Y(n_1080)
);

AO21x2_ASAP7_75t_L g1081 ( 
.A1(n_1030),
.A2(n_959),
.B(n_956),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_1007),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_984),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_1017),
.A2(n_956),
.B(n_959),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1015),
.B(n_496),
.Y(n_1085)
);

INVx6_ASAP7_75t_SL g1086 ( 
.A(n_997),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_1023),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1045),
.A2(n_1042),
.B(n_1004),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1003),
.A2(n_364),
.B(n_78),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_1024),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_987),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1005),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1049),
.B(n_364),
.Y(n_1093)
);

OA21x2_ASAP7_75t_L g1094 ( 
.A1(n_981),
.A2(n_364),
.B(n_558),
.Y(n_1094)
);

BUFx2_ASAP7_75t_SL g1095 ( 
.A(n_985),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_998),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_1040),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_975),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1039),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_1044),
.Y(n_1100)
);

AO21x2_ASAP7_75t_L g1101 ( 
.A1(n_990),
.A2(n_364),
.B(n_560),
.Y(n_1101)
);

INVx8_ASAP7_75t_L g1102 ( 
.A(n_996),
.Y(n_1102)
);

AO21x1_ASAP7_75t_L g1103 ( 
.A1(n_1033),
.A2(n_364),
.B(n_79),
.Y(n_1103)
);

BUFx5_ASAP7_75t_L g1104 ( 
.A(n_989),
.Y(n_1104)
);

BUFx2_ASAP7_75t_SL g1105 ( 
.A(n_1046),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1011),
.B(n_560),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_989),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_1048),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_989),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1054),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1014),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1000),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1051),
.A2(n_81),
.B(n_83),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1025),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1035),
.A2(n_93),
.B(n_99),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_1026),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_1098),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1079),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1082),
.B(n_1037),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_1060),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_1086),
.Y(n_1121)
);

INVx6_ASAP7_75t_L g1122 ( 
.A(n_1102),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1069),
.B(n_1013),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1108),
.B(n_995),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1078),
.Y(n_1125)
);

INVx6_ASAP7_75t_L g1126 ( 
.A(n_1102),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1067),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1065),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1067),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1102),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1111),
.A2(n_1027),
.B1(n_1031),
.B2(n_1038),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1098),
.A2(n_992),
.B1(n_1053),
.B2(n_1020),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_1063),
.Y(n_1133)
);

NAND2x1p5_ASAP7_75t_L g1134 ( 
.A(n_1055),
.B(n_1047),
.Y(n_1134)
);

BUFx10_ASAP7_75t_L g1135 ( 
.A(n_1073),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_1087),
.B(n_1012),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1057),
.A2(n_1050),
.B(n_1008),
.Y(n_1137)
);

BUFx4f_ASAP7_75t_SL g1138 ( 
.A(n_1086),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_1056),
.B(n_1010),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1112),
.A2(n_1080),
.B1(n_1107),
.B2(n_1109),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1077),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1081),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1112),
.A2(n_1029),
.B1(n_1034),
.B2(n_583),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_SL g1144 ( 
.A1(n_1087),
.A2(n_583),
.B1(n_580),
.B2(n_102),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1081),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1077),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1077),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1077),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_SL g1149 ( 
.A(n_1113),
.B(n_100),
.C(n_101),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1099),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_1070),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1068),
.A2(n_583),
.B(n_580),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1100),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1110),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1099),
.Y(n_1155)
);

CKINVDCx14_ASAP7_75t_R g1156 ( 
.A(n_1090),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1062),
.A2(n_580),
.B1(n_105),
.B2(n_106),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1099),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1066),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_1058),
.A2(n_104),
.B(n_107),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1071),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1072),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1114),
.A2(n_111),
.B1(n_113),
.B2(n_121),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1073),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1064),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1114),
.A2(n_135),
.B1(n_136),
.B2(n_139),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1083),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_1063),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1097),
.B(n_148),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1105),
.A2(n_149),
.B1(n_151),
.B2(n_154),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1088),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1118),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1132),
.A2(n_1149),
.B(n_1113),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1127),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1117),
.B(n_1091),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1124),
.B(n_1064),
.Y(n_1176)
);

NAND2xp33_ASAP7_75t_R g1177 ( 
.A(n_1121),
.B(n_1096),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1117),
.A2(n_1116),
.B1(n_1076),
.B2(n_1093),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1125),
.Y(n_1179)
);

NOR3xp33_ASAP7_75t_SL g1180 ( 
.A(n_1120),
.B(n_1085),
.C(n_1116),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1161),
.B(n_1129),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1119),
.B(n_1069),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1120),
.Y(n_1183)
);

NAND2xp33_ASAP7_75t_L g1184 ( 
.A(n_1132),
.B(n_1116),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1156),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1128),
.B(n_1095),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1154),
.B(n_1096),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1158),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1136),
.B(n_1076),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1167),
.B(n_1107),
.Y(n_1190)
);

CKINVDCx16_ASAP7_75t_R g1191 ( 
.A(n_1130),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_1138),
.Y(n_1192)
);

OR2x6_ASAP7_75t_L g1193 ( 
.A(n_1150),
.B(n_1059),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1122),
.Y(n_1194)
);

INVx2_ASAP7_75t_R g1195 ( 
.A(n_1141),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1164),
.B(n_1074),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_1130),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1123),
.B(n_1075),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1130),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1168),
.B(n_1106),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1162),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1153),
.A2(n_1104),
.B1(n_1061),
.B2(n_1092),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1133),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1122),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1159),
.A2(n_1140),
.A3(n_1143),
.B(n_1103),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1135),
.B(n_1104),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1155),
.B(n_1126),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1140),
.A2(n_1092),
.A3(n_1104),
.B(n_1058),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_SL g1209 ( 
.A1(n_1144),
.A2(n_1166),
.B1(n_1163),
.B2(n_1165),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1169),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1134),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1134),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1147),
.B(n_1084),
.Y(n_1213)
);

AND2x4_ASAP7_75t_SL g1214 ( 
.A(n_1193),
.B(n_1180),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1210),
.B(n_1148),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1176),
.B(n_1146),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1188),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1175),
.B(n_1160),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1208),
.Y(n_1219)
);

AOI221xp5_ASAP7_75t_L g1220 ( 
.A1(n_1173),
.A2(n_1131),
.B1(n_1143),
.B2(n_1166),
.C(n_1163),
.Y(n_1220)
);

AOI33xp33_ASAP7_75t_L g1221 ( 
.A1(n_1202),
.A2(n_1144),
.A3(n_1170),
.B1(n_1157),
.B2(n_1131),
.B3(n_1139),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1189),
.B(n_1142),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1174),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1172),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1182),
.B(n_1145),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1208),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1186),
.B(n_1151),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1184),
.B(n_1139),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1206),
.B(n_1145),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1181),
.B(n_1171),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1213),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1208),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1200),
.B(n_1094),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1199),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1187),
.B(n_1101),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1190),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1211),
.A2(n_1152),
.A3(n_1137),
.B(n_1089),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1190),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1201),
.B(n_1115),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1179),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1212),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1213),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1205),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1205),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1205),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1195),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1194),
.B(n_155),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1191),
.B(n_158),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1207),
.B(n_159),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1196),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1194),
.B(n_160),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1203),
.B(n_166),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1198),
.B(n_167),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1178),
.B(n_168),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1199),
.B(n_170),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1220),
.A2(n_1209),
.B1(n_1204),
.B2(n_1185),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1224),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1217),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1241),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1242),
.B(n_1197),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1231),
.B(n_1227),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1231),
.B(n_1197),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1223),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1218),
.B(n_1183),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1238),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1236),
.B(n_1192),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1238),
.B(n_172),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1245),
.B(n_173),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1245),
.B(n_174),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1241),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1215),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1230),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1225),
.B(n_1177),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1240),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1222),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1233),
.B(n_176),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1229),
.B(n_181),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1272),
.B(n_1235),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1261),
.B(n_1246),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1259),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1271),
.B(n_1216),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1257),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1264),
.B(n_1243),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1259),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1263),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1275),
.B(n_1250),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1270),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1273),
.B(n_1244),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1258),
.B(n_1219),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1260),
.B(n_1219),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1262),
.B(n_1214),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1273),
.B(n_1226),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1291),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1283),
.A2(n_1256),
.B1(n_1228),
.B2(n_1214),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1278),
.B(n_1266),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1280),
.Y(n_1296)
);

INVxp67_ASAP7_75t_SL g1297 ( 
.A(n_1289),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1280),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1282),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1281),
.A2(n_1269),
.B1(n_1268),
.B2(n_1248),
.Y(n_1300)
);

AO221x1_ASAP7_75t_L g1301 ( 
.A1(n_1285),
.A2(n_1265),
.B1(n_1234),
.B2(n_1226),
.C(n_1232),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1296),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1301),
.A2(n_1288),
.B1(n_1292),
.B2(n_1254),
.Y(n_1303)
);

AOI211xp5_ASAP7_75t_SL g1304 ( 
.A1(n_1293),
.A2(n_1291),
.B(n_1290),
.C(n_1279),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1300),
.A2(n_1221),
.B(n_1276),
.C(n_1277),
.Y(n_1305)
);

OAI211xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1295),
.A2(n_1221),
.B(n_1252),
.C(n_1286),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1294),
.A2(n_1232),
.B1(n_1274),
.B2(n_1284),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1298),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1299),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_1297),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1309),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1309),
.Y(n_1312)
);

AOI211x1_ASAP7_75t_SL g1313 ( 
.A1(n_1305),
.A2(n_1253),
.B(n_1234),
.C(n_1284),
.Y(n_1313)
);

AOI21xp33_ASAP7_75t_L g1314 ( 
.A1(n_1306),
.A2(n_1249),
.B(n_1267),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1310),
.A2(n_1247),
.B(n_1251),
.C(n_1255),
.Y(n_1315)
);

NOR3xp33_ASAP7_75t_L g1316 ( 
.A(n_1302),
.B(n_1308),
.C(n_1239),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1303),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1311),
.Y(n_1318)
);

NOR3x1_ASAP7_75t_L g1319 ( 
.A(n_1317),
.B(n_1304),
.C(n_1307),
.Y(n_1319)
);

NOR2x1_ASAP7_75t_SL g1320 ( 
.A(n_1312),
.B(n_1287),
.Y(n_1320)
);

NOR2x1_ASAP7_75t_L g1321 ( 
.A(n_1318),
.B(n_1315),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1319),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1321),
.B(n_1316),
.Y(n_1323)
);

AOI31xp33_ASAP7_75t_L g1324 ( 
.A1(n_1322),
.A2(n_1314),
.A3(n_1320),
.B(n_1313),
.Y(n_1324)
);

OAI221xp5_ASAP7_75t_L g1325 ( 
.A1(n_1322),
.A2(n_1237),
.B1(n_193),
.B2(n_195),
.C(n_198),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1323),
.Y(n_1326)
);

NOR2xp67_ASAP7_75t_L g1327 ( 
.A(n_1325),
.B(n_1324),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1327),
.A2(n_1237),
.B1(n_220),
.B2(n_221),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1326),
.B(n_290),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1329),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1328),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1330),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1331),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1332),
.B(n_229),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1333),
.Y(n_1335)
);

OAI22x1_ASAP7_75t_L g1336 ( 
.A1(n_1335),
.A2(n_247),
.B1(n_249),
.B2(n_251),
.Y(n_1336)
);

NAND2xp33_ASAP7_75t_R g1337 ( 
.A(n_1334),
.B(n_255),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1336),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1338),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1339),
.A2(n_1337),
.B1(n_260),
.B2(n_261),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1340),
.B(n_272),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1341),
.A2(n_277),
.B1(n_278),
.B2(n_282),
.Y(n_1342)
);


endmodule