module real_jpeg_33560_n_7 (n_5, n_4, n_0, n_1, n_26, n_2, n_27, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_26;
input n_2;
input n_27;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_23;
wire n_11;
wire n_14;
wire n_22;
wire n_18;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

OAI221xp5_ASAP7_75t_L g10 ( 
.A1(n_0),
.A2(n_11),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_10)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g7 ( 
.A1(n_1),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_2),
.B(n_26),
.Y(n_13)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_6),
.C(n_12),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

INVxp33_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.C(n_15),
.Y(n_12)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_27),
.Y(n_14)
);


endmodule