module fake_jpeg_7781_n_335 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_25),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_27),
.B1(n_18),
.B2(n_22),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_48),
.A2(n_38),
.B1(n_46),
.B2(n_26),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_65),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_27),
.B1(n_22),
.B2(n_30),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_22),
.B1(n_30),
.B2(n_17),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_16),
.Y(n_95)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_49),
.B(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_79),
.Y(n_105)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_93),
.Y(n_128)
);

NAND2x1_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_44),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_89),
.C(n_90),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_44),
.C(n_39),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_44),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_47),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_40),
.B1(n_66),
.B2(n_58),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_14),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_97),
.B1(n_21),
.B2(n_20),
.Y(n_111)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_53),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_46),
.B1(n_38),
.B2(n_71),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_112),
.B1(n_98),
.B2(n_83),
.Y(n_133)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_106),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_36),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_111),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_39),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_110),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_39),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_46),
.B1(n_38),
.B2(n_40),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_119),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_87),
.B1(n_76),
.B2(n_46),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_118),
.B1(n_40),
.B2(n_84),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_46),
.B1(n_38),
.B2(n_53),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_74),
.B(n_38),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_91),
.B1(n_40),
.B2(n_90),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_127),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_87),
.A2(n_40),
.B1(n_29),
.B2(n_17),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_86),
.B(n_93),
.Y(n_139)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_36),
.CI(n_44),
.CON(n_127),
.SN(n_127)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_133),
.B1(n_123),
.B2(n_118),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_122),
.A2(n_91),
.B1(n_40),
.B2(n_90),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_131),
.A2(n_134),
.B(n_139),
.Y(n_179)
);

OAI31xp33_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_96),
.A3(n_90),
.B(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_145),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_141),
.B1(n_146),
.B2(n_124),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_79),
.B1(n_42),
.B2(n_47),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_36),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_147),
.B(n_121),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_120),
.B(n_116),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_36),
.B(n_23),
.Y(n_180)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_77),
.B1(n_52),
.B2(n_56),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_36),
.B(n_95),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_79),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_153),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_101),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_156),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_36),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_106),
.C(n_103),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_43),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_43),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_43),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_110),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_147),
.B(n_179),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_128),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_160),
.C(n_162),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_161),
.B(n_180),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_99),
.C(n_115),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_183),
.B1(n_185),
.B2(n_151),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_112),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_181),
.C(n_162),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_178),
.B1(n_132),
.B2(n_148),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_174),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_114),
.B1(n_52),
.B2(n_60),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_173),
.A2(n_184),
.B1(n_42),
.B2(n_100),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_108),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_149),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_114),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_177),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_133),
.A2(n_126),
.B1(n_80),
.B2(n_17),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_80),
.C(n_92),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_155),
.A2(n_47),
.B1(n_43),
.B2(n_42),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_47),
.B1(n_43),
.B2(n_42),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_42),
.B1(n_35),
.B2(n_33),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_195),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_197),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_202),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_199),
.B1(n_161),
.B2(n_180),
.Y(n_215)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NOR2x1_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_134),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_203),
.C(n_204),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_139),
.B(n_130),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_201),
.B(n_207),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_143),
.A3(n_154),
.B1(n_138),
.B2(n_145),
.C1(n_148),
.C2(n_135),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_143),
.C(n_135),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_154),
.C(n_125),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_177),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_183),
.B1(n_164),
.B2(n_185),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_82),
.C(n_36),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_184),
.C(n_174),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_32),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_157),
.B(n_29),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_212),
.A2(n_176),
.B1(n_171),
.B2(n_25),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_214),
.A2(n_224),
.B1(n_233),
.B2(n_236),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_190),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_197),
.A2(n_171),
.B1(n_178),
.B2(n_182),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_226),
.B1(n_204),
.B2(n_25),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_172),
.B1(n_175),
.B2(n_169),
.Y(n_218)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_228),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_229),
.C(n_237),
.Y(n_244)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

AO22x2_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_158),
.B1(n_32),
.B2(n_33),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_82),
.C(n_23),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_230),
.B(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_187),
.A2(n_35),
.B1(n_32),
.B2(n_33),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_238),
.B1(n_239),
.B2(n_206),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_23),
.C(n_28),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_188),
.B1(n_194),
.B2(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_260),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_209),
.B1(n_196),
.B2(n_212),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_246),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_189),
.C(n_210),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_253),
.C(n_255),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_221),
.A2(n_196),
.B1(n_192),
.B2(n_199),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g252 ( 
.A1(n_220),
.A2(n_189),
.B(n_25),
.C(n_163),
.D(n_23),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_214),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_28),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_254),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_23),
.C(n_28),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_220),
.B(n_23),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_257),
.B(n_251),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_223),
.C(n_228),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_261),
.C(n_235),
.Y(n_270)
);

FAx1_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_23),
.CI(n_34),
.CON(n_260),
.SN(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_225),
.C(n_216),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_240),
.A2(n_226),
.B1(n_227),
.B2(n_231),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_262),
.A2(n_276),
.B1(n_260),
.B2(n_255),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_236),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_271),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_224),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_278),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_244),
.C(n_249),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_233),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_9),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_0),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_16),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_0),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_289),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_261),
.B(n_241),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_294),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_259),
.B(n_244),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_286),
.C(n_279),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_257),
.B1(n_260),
.B2(n_252),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_273),
.B1(n_263),
.B2(n_262),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_269),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_290),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_253),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_269),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_11),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_34),
.C(n_16),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_293),
.C(n_12),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_14),
.C(n_13),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_270),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_302),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_272),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_297),
.B(n_283),
.Y(n_311)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_277),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_297),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_317)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_276),
.B1(n_264),
.B2(n_274),
.Y(n_299)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_304),
.C(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_12),
.C(n_11),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_281),
.B(n_10),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_10),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_314),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_311),
.A2(n_3),
.B(n_6),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_312),
.B(n_317),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_10),
.C(n_1),
.Y(n_314)
);

AOI221xp5_ASAP7_75t_L g316 ( 
.A1(n_296),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_302),
.B(n_307),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_303),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_321),
.B(n_323),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_301),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_318),
.B1(n_316),
.B2(n_321),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_2),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_313),
.C(n_7),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_6),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_6),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_329),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_319),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_328),
.B(n_7),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_332),
.B(n_330),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_7),
.B1(n_8),
.B2(n_326),
.Y(n_335)
);


endmodule