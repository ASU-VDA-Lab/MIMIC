module fake_jpeg_8088_n_34 (n_3, n_2, n_1, n_0, n_4, n_5, n_34);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_3),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_5),
.Y(n_7)
);

INVx2_ASAP7_75t_SL g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

OR2x2_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_8),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_6),
.C(n_9),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_15),
.B(n_9),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.C(n_24),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_21),
.B1(n_8),
.B2(n_11),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_28),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_17),
.C(n_19),
.Y(n_28)
);

AOI322xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_16),
.A3(n_13),
.B1(n_14),
.B2(n_10),
.C1(n_11),
.C2(n_5),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B(n_8),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_10),
.B(n_8),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B(n_4),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_2),
.B(n_4),
.Y(n_33)
);


endmodule