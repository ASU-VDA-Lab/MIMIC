module fake_jpeg_4279_n_114 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

INVx6_ASAP7_75t_SL g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_13),
.B1(n_14),
.B2(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_9),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_19),
.C(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_23),
.C(n_18),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_14),
.B(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_46),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_28),
.B1(n_26),
.B2(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_29),
.B1(n_26),
.B2(n_28),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_43),
.Y(n_51)
);

BUFx24_ASAP7_75t_SL g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_26),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_57),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_50),
.A3(n_48),
.B1(n_45),
.B2(n_44),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_26),
.B(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_9),
.Y(n_66)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_28),
.Y(n_59)
);

NOR3xp33_ASAP7_75t_SL g61 ( 
.A(n_59),
.B(n_20),
.C(n_22),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_28),
.B1(n_16),
.B2(n_9),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_66),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_21),
.A3(n_22),
.B1(n_20),
.B2(n_29),
.C1(n_30),
.C2(n_16),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_30),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_13),
.B(n_14),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_71),
.B(n_17),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_8),
.B(n_7),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_70),
.B(n_8),
.Y(n_81)
);

AOI322xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_16),
.A3(n_9),
.B1(n_21),
.B2(n_29),
.C1(n_8),
.C2(n_5),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_13),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_77),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_58),
.B(n_57),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_67),
.B1(n_15),
.B2(n_12),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_81),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_30),
.C(n_42),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_79),
.C(n_82),
.Y(n_84)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_72),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_30),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_17),
.B(n_12),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_69),
.C(n_65),
.Y(n_82)
);

AOI322xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_65),
.A3(n_67),
.B1(n_15),
.B2(n_17),
.C1(n_12),
.C2(n_5),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_85),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_79),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_15),
.B1(n_12),
.B2(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_75),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_15),
.C(n_1),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_82),
.C(n_1),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_93),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_96),
.C(n_84),
.Y(n_98)
);

AOI31xp67_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_90),
.A3(n_85),
.B(n_87),
.Y(n_97)
);

NAND2xp67_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_91),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_84),
.C(n_88),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_101),
.B(n_0),
.C(n_3),
.Y(n_107)
);

NOR2xp67_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_94),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_107),
.B(n_0),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_15),
.B1(n_1),
.B2(n_3),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_106),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_0),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_107),
.C(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_0),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_4),
.C(n_6),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_112),
.B(n_109),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_4),
.Y(n_114)
);


endmodule