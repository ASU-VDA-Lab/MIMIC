module fake_jpeg_32189_n_484 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_484);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_484;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

BUFx12f_ASAP7_75t_SL g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_53),
.B(n_58),
.Y(n_122)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_20),
.A2(n_6),
.B(n_11),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_64),
.B(n_65),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_18),
.B(n_6),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_75),
.Y(n_160)
);

NAND2x1_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_9),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_76),
.B(n_0),
.Y(n_127)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_41),
.B(n_9),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_80),
.B(n_84),
.Y(n_153)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_18),
.B(n_4),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_4),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_92),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_10),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_16),
.Y(n_93)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_26),
.B(n_10),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_96),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_26),
.B(n_10),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

BUFx4f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_99),
.Y(n_129)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_27),
.B(n_10),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_33),
.Y(n_121)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_27),
.B(n_11),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_39),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_112),
.B(n_121),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_152),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_143),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_80),
.A2(n_15),
.B1(n_49),
.B2(n_48),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_140),
.B1(n_151),
.B2(n_46),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_83),
.A2(n_49),
.B1(n_30),
.B2(n_32),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_67),
.A2(n_49),
.B1(n_42),
.B2(n_32),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_141),
.A2(n_144),
.B1(n_98),
.B2(n_87),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_76),
.A2(n_16),
.B(n_22),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_77),
.A2(n_102),
.B1(n_73),
.B2(n_104),
.Y(n_144)
);

BUFx10_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_148),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_35),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_60),
.A2(n_39),
.B1(n_47),
.B2(n_33),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_70),
.B(n_28),
.Y(n_152)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_117),
.A2(n_159),
.B1(n_107),
.B2(n_126),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_166),
.A2(n_197),
.B1(n_138),
.B2(n_144),
.Y(n_214)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

AO22x2_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_42),
.B1(n_66),
.B2(n_74),
.Y(n_170)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_170),
.B(n_42),
.Y(n_245)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_172),
.B(n_191),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_153),
.C(n_146),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_174),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_37),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_142),
.A2(n_71),
.B1(n_55),
.B2(n_103),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_179),
.A2(n_210),
.B1(n_211),
.B2(n_161),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_183),
.Y(n_215)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_135),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_192),
.Y(n_247)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

BUFx24_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_116),
.B(n_28),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_195),
.B(n_198),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_131),
.B(n_68),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_132),
.B(n_47),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_148),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_201),
.Y(n_223)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_133),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_122),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_203),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_204),
.A2(n_207),
.B1(n_209),
.B2(n_129),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_122),
.B(n_40),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_213),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_120),
.B(n_89),
.C(n_88),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_129),
.B(n_123),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_139),
.Y(n_207)
);

AO22x1_ASAP7_75t_L g208 ( 
.A1(n_140),
.A2(n_75),
.B1(n_62),
.B2(n_91),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_141),
.B(n_161),
.C(n_46),
.Y(n_235)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_133),
.A2(n_86),
.B1(n_62),
.B2(n_32),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_114),
.B(n_40),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_214),
.A2(n_218),
.B1(n_179),
.B2(n_211),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_138),
.B1(n_157),
.B2(n_137),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_219),
.A2(n_238),
.B1(n_184),
.B2(n_210),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_51),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_228),
.B(n_232),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_51),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_235),
.B(n_183),
.Y(n_261)
);

OAI22x1_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_123),
.B1(n_160),
.B2(n_155),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_157),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_246),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_170),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_174),
.B(n_137),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_196),
.B1(n_166),
.B2(n_170),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_251),
.A2(n_245),
.B1(n_233),
.B2(n_229),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_173),
.C(n_206),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_230),
.C(n_235),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_246),
.B(n_170),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_255),
.B(n_259),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_256),
.A2(n_264),
.B(n_274),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_220),
.B(n_177),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_262),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_238),
.B1(n_264),
.B2(n_263),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_191),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_261),
.B(n_265),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_169),
.Y(n_262)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_239),
.B(n_168),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_217),
.B(n_175),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_267),
.B(n_275),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_223),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_269),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_270),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_186),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_215),
.A2(n_181),
.B(n_113),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_232),
.B(n_35),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_245),
.A2(n_162),
.B1(n_111),
.B2(n_201),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_277),
.A2(n_229),
.B1(n_241),
.B2(n_245),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_215),
.B(n_167),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_234),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_243),
.B(n_45),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_224),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_285),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_286),
.B(n_265),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_301),
.C(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_290),
.B(n_259),
.Y(n_319)
);

XOR2x2_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_245),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_252),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_270),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_294),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_296),
.A2(n_299),
.B1(n_251),
.B2(n_253),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_300),
.B1(n_308),
.B2(n_277),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_270),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_298),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_251),
.A2(n_255),
.B1(n_256),
.B2(n_279),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_249),
.C(n_244),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_265),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_265),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_252),
.B(n_249),
.C(n_244),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_256),
.A2(n_224),
.B1(n_194),
.B2(n_241),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_309),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_293),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_316),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_312),
.A2(n_292),
.B1(n_300),
.B2(n_301),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_297),
.A2(n_278),
.B1(n_258),
.B2(n_268),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_315),
.B(n_321),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_278),
.B1(n_256),
.B2(n_261),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_281),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_283),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_327),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_328),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_276),
.Y(n_320)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_284),
.A2(n_274),
.B(n_278),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_322),
.A2(n_324),
.B1(n_329),
.B2(n_254),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_323),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_299),
.A2(n_289),
.B1(n_284),
.B2(n_304),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_287),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_326),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_305),
.B(n_257),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_292),
.A2(n_265),
.B1(n_275),
.B2(n_271),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_293),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_333),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_332),
.B(n_247),
.Y(n_362)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_280),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_286),
.C(n_291),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_273),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_295),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_336),
.A2(n_339),
.B1(n_343),
.B2(n_347),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_341),
.C(n_344),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_312),
.A2(n_288),
.B1(n_283),
.B2(n_302),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_288),
.C(n_290),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_313),
.A2(n_315),
.B1(n_327),
.B2(n_323),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_253),
.C(n_303),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_307),
.C(n_303),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_352),
.C(n_355),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_311),
.A2(n_307),
.B1(n_302),
.B2(n_298),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_320),
.A2(n_331),
.B1(n_309),
.B2(n_322),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_348),
.A2(n_212),
.B1(n_109),
.B2(n_154),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_266),
.C(n_272),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_353),
.A2(n_333),
.B1(n_326),
.B2(n_319),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_294),
.C(n_281),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_321),
.A2(n_295),
.B(n_231),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_357),
.A2(n_314),
.B(n_330),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_317),
.B(n_260),
.Y(n_358)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_324),
.B(n_247),
.C(n_221),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_240),
.C(n_190),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_314),
.B(n_330),
.Y(n_361)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_361),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_362),
.B(n_329),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_310),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_365),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_335),
.Y(n_366)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_366),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_336),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_357),
.A2(n_316),
.B(n_318),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_368),
.A2(n_338),
.B(n_346),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_370),
.A2(n_375),
.B1(n_388),
.B2(n_347),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_356),
.B(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_371),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g372 ( 
.A(n_362),
.B(n_222),
.CI(n_225),
.CON(n_372),
.SN(n_372)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_372),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_353),
.A2(n_260),
.B1(n_236),
.B2(n_221),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_236),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_360),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_361),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_378),
.A2(n_380),
.B1(n_386),
.B2(n_389),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_381),
.C(n_385),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_342),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_240),
.C(n_204),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_351),
.B(n_237),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_358),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_200),
.C(n_145),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_338),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_0),
.Y(n_387)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_387),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_359),
.A2(n_45),
.B1(n_37),
.B2(n_22),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_390),
.A2(n_377),
.B1(n_363),
.B2(n_389),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_397),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_396),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_355),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_406),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_341),
.C(n_352),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_400),
.C(n_403),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_381),
.B(n_337),
.C(n_343),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_369),
.B(n_350),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_385),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_346),
.C(n_350),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_376),
.B(n_339),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_366),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_407),
.B(n_410),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_356),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_367),
.C(n_379),
.Y(n_421)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_409),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_413),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_393),
.A2(n_370),
.B1(n_374),
.B2(n_384),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_401),
.A2(n_375),
.B1(n_359),
.B2(n_382),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_418),
.Y(n_436)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_392),
.Y(n_417)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_363),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_405),
.A2(n_382),
.B1(n_368),
.B2(n_377),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_421),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_216),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_365),
.C(n_372),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_424),
.B(n_400),
.C(n_403),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_SL g425 ( 
.A1(n_407),
.A2(n_349),
.B(n_354),
.C(n_372),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_425),
.A2(n_419),
.B1(n_422),
.B2(n_411),
.Y(n_433)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

NAND3xp33_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_349),
.C(n_340),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_429),
.B(n_434),
.Y(n_450)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_430),
.Y(n_445)
);

FAx1_ASAP7_75t_SL g431 ( 
.A(n_425),
.B(n_424),
.CI(n_394),
.CON(n_431),
.SN(n_431)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_426),
.Y(n_444)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_433),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_414),
.A2(n_406),
.B(n_398),
.Y(n_434)
);

AOI21x1_ASAP7_75t_L g435 ( 
.A1(n_425),
.A2(n_387),
.B(n_408),
.Y(n_435)
);

AOI21xp33_ASAP7_75t_L g453 ( 
.A1(n_435),
.A2(n_17),
.B(n_13),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_395),
.C(n_399),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_437),
.B(n_438),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_420),
.A2(n_397),
.B(n_410),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_421),
.A2(n_216),
.B(n_237),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_439),
.B(n_415),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_440),
.A2(n_442),
.B1(n_428),
.B2(n_443),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_216),
.C(n_237),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_441),
.B(n_415),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_216),
.B(n_13),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_442),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_13),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_456),
.Y(n_465)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_447),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_449),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_437),
.B(n_212),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_434),
.B(n_431),
.Y(n_451)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_451),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_453),
.B(n_455),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_17),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_432),
.A2(n_429),
.B1(n_433),
.B2(n_431),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_445),
.A2(n_441),
.B1(n_428),
.B2(n_440),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_458),
.B(n_459),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_32),
.C(n_57),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_463),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_450),
.B(n_32),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_61),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_457),
.B(n_455),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_466),
.A2(n_452),
.B(n_1),
.Y(n_472)
);

NOR2x1_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_446),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_468),
.A2(n_472),
.B(n_474),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_471),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_470),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_465),
.B(n_444),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_467),
.A2(n_452),
.B(n_1),
.Y(n_474)
);

A2O1A1O1Ixp25_ASAP7_75t_L g476 ( 
.A1(n_473),
.A2(n_462),
.B(n_466),
.C(n_464),
.D(n_0),
.Y(n_476)
);

AO21x1_ASAP7_75t_L g480 ( 
.A1(n_476),
.A2(n_1),
.B(n_2),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_478),
.B(n_473),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_479),
.A2(n_480),
.B(n_475),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_481),
.B(n_477),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_482),
.A2(n_1),
.B(n_2),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_483),
.A2(n_2),
.B(n_361),
.Y(n_484)
);


endmodule