module real_jpeg_26266_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_0),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.Y(n_103)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_2),
.B(n_69),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_2),
.B(n_36),
.C(n_38),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_72),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_2),
.B(n_41),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_72),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_2),
.B(n_49),
.C(n_52),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_2),
.A2(n_83),
.B(n_171),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_4),
.A2(n_27),
.B1(n_62),
.B2(n_67),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_4),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_4),
.A2(n_27),
.B1(n_49),
.B2(n_53),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_7),
.A2(n_28),
.B1(n_31),
.B2(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_7),
.A2(n_43),
.B1(n_49),
.B2(n_53),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_49),
.B1(n_53),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_10),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_87),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_12),
.A2(n_49),
.B1(n_53),
.B2(n_91),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_12),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_13),
.A2(n_49),
.B1(n_53),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_14),
.A2(n_58),
.B1(n_71),
.B2(n_77),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_28),
.B1(n_31),
.B2(n_58),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_14),
.A2(n_49),
.B1(n_53),
.B2(n_58),
.Y(n_140)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_15),
.Y(n_138)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_15),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_128),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_20),
.B(n_104),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_95),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_21),
.A2(n_22),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_59),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_25),
.B(n_44),
.C(n_59),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_26),
.Y(n_97)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_28),
.A2(n_31),
.B1(n_65),
.B2(n_66),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_28),
.A2(n_65),
.B(n_73),
.C(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_28),
.B(n_134),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_SL g94 ( 
.A(n_31),
.B(n_66),
.C(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_32),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_33),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_33),
.A2(n_110),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_40),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_34),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_36),
.B1(n_51),
.B2(n_52),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_36),
.B(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_41),
.B(n_99),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_42),
.Y(n_109)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B(n_54),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_46),
.A2(n_48),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_48),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_48),
.A2(n_54),
.B(n_143),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_48),
.B(n_72),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_84),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_53),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_55),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_57),
.B(n_145),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_70),
.B(n_75),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_112),
.B(n_114),
.Y(n_111)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_73),
.Y(n_70)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_72),
.B(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_78),
.A2(n_79),
.B1(n_95),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_92),
.B2(n_93),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_92),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_88),
.B2(n_90),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_82),
.A2(n_183),
.B1(n_185),
.B2(n_187),
.Y(n_182)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_86),
.B1(n_89),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_89),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_83),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_84),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_89),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_95),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_102),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_96),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_116),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_125),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_123),
.A2(n_159),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_212),
.B(n_218),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_160),
.B(n_211),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_149),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_131),
.B(n_149),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_141),
.C(n_146),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_132),
.B(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_135),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B(n_139),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_139),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_140),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_141),
.A2(n_146),
.B1(n_147),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_150),
.B(n_156),
.C(n_157),
.Y(n_217)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_205),
.B(n_210),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_180),
.B(n_204),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_174),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_174),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_190),
.B(n_203),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_188),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_194),
.B(n_195),
.Y(n_193)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_196),
.B(n_202),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_209),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_217),
.Y(n_218)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);


endmodule