module real_jpeg_23329_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_1),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_1),
.A2(n_22),
.B1(n_27),
.B2(n_87),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_1),
.A2(n_63),
.B1(n_65),
.B2(n_87),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_1),
.A2(n_54),
.B1(n_58),
.B2(n_87),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_30),
.B1(n_80),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_2),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_2),
.A2(n_22),
.B1(n_27),
.B2(n_121),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_2),
.A2(n_63),
.B1(n_65),
.B2(n_121),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_2),
.A2(n_54),
.B1(n_58),
.B2(n_121),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_3),
.B(n_30),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_3),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_3),
.B(n_21),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_3),
.B(n_63),
.C(n_93),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_3),
.A2(n_22),
.B1(n_27),
.B2(n_222),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_3),
.B(n_136),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_3),
.A2(n_63),
.B1(n_65),
.B2(n_222),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_3),
.B(n_54),
.C(n_68),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_3),
.A2(n_53),
.B(n_284),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_7),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_7),
.A2(n_63),
.B1(n_65),
.B2(n_97),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_7),
.A2(n_32),
.B1(n_80),
.B2(n_97),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_7),
.A2(n_54),
.B1(n_58),
.B2(n_97),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_9),
.A2(n_42),
.B1(n_63),
.B2(n_65),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_9),
.A2(n_42),
.B1(n_54),
.B2(n_58),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_9),
.A2(n_22),
.B1(n_27),
.B2(n_42),
.Y(n_138)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_11),
.A2(n_30),
.B1(n_81),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_11),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_11),
.A2(n_22),
.B1(n_27),
.B2(n_170),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_11),
.A2(n_63),
.B1(n_65),
.B2(n_170),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_11),
.A2(n_54),
.B1(n_58),
.B2(n_170),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_12),
.A2(n_22),
.B1(n_27),
.B2(n_62),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_12),
.A2(n_30),
.B1(n_62),
.B2(n_81),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_12),
.A2(n_54),
.B1(n_58),
.B2(n_62),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_13),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_13),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_13),
.A2(n_22),
.B1(n_27),
.B2(n_82),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_13),
.A2(n_63),
.B1(n_65),
.B2(n_82),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_13),
.A2(n_54),
.B1(n_58),
.B2(n_82),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_15),
.A2(n_35),
.B1(n_54),
.B2(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_15),
.A2(n_35),
.B1(n_63),
.B2(n_65),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_15),
.A2(n_22),
.B1(n_27),
.B2(n_35),
.Y(n_158)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_16),
.Y(n_199)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_16),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_16),
.A2(n_195),
.B1(n_296),
.B2(n_298),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_45),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_43),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_34),
.Y(n_20)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_21),
.A2(n_28),
.B1(n_34),
.B2(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_21),
.A2(n_28),
.B1(n_120),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_21),
.A2(n_28),
.B1(n_41),
.B2(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_22),
.A2(n_27),
.B1(n_93),
.B2(n_94),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g193 ( 
.A(n_22),
.B(n_26),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_22),
.B(n_247),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g191 ( 
.A1(n_25),
.A2(n_27),
.A3(n_80),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_28),
.B(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_28),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_28),
.A2(n_124),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_33),
.A2(n_78),
.B(n_83),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_33),
.B(n_85),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_33),
.A2(n_78),
.B1(n_122),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_33),
.A2(n_122),
.B1(n_144),
.B2(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_33),
.A2(n_83),
.B(n_185),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_SL g221 ( 
.A1(n_36),
.A2(n_222),
.B(n_223),
.Y(n_221)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_40),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_40),
.B(n_356),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_355),
.B(n_357),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_343),
.B(n_354),
.Y(n_46)
);

OAI31xp33_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_146),
.A3(n_160),
.B(n_340),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_125),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_49),
.B(n_125),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_88),
.C(n_104),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_50),
.A2(n_88),
.B1(n_89),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_50),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_74),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_51),
.A2(n_52),
.B(n_76),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_52),
.A2(n_59),
.B1(n_60),
.B2(n_75),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_56),
.B(n_57),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_53),
.A2(n_57),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_53),
.A2(n_55),
.B1(n_109),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_53),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_53),
.A2(n_197),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_53),
.B(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_53),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_58),
.B1(n_68),
.B2(n_70),
.Y(n_71)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_55),
.Y(n_252)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_56),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_56),
.B(n_222),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_58),
.B(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_61),
.A2(n_66),
.B1(n_73),
.B2(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_63),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_65),
.B1(n_68),
.B2(n_70),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_65),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_63),
.B(n_292),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_66),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_66),
.A2(n_73),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_66),
.B(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_66),
.A2(n_73),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_71),
.A2(n_100),
.B1(n_115),
.B2(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_71),
.A2(n_180),
.B(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_71),
.A2(n_218),
.B(n_257),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_71),
.B(n_222),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_73),
.B(n_219),
.Y(n_272)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B(n_103),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_98),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_91),
.A2(n_92),
.B1(n_138),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_91),
.A2(n_187),
.B(n_189),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_91),
.A2(n_189),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_92),
.A2(n_117),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_92),
.A2(n_173),
.B(n_227),
.Y(n_226)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_100),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_100),
.A2(n_272),
.B(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_102),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_104),
.A2(n_105),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.C(n_118),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_106),
.A2(n_107),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_108),
.A2(n_112),
.B1(n_113),
.B2(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_108),
.Y(n_182)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_116),
.B(n_118),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B(n_123),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_128),
.C(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_143),
.B2(n_145),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_140),
.C(n_143),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_135),
.A2(n_136),
.B1(n_188),
.B2(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_135),
.A2(n_136),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_136),
.B(n_174),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_140),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_140),
.B(n_153),
.C(n_157),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_143),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_145),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_143),
.B(n_149),
.C(n_152),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_147),
.A2(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_159),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_148),
.B(n_159),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_154),
.Y(n_350)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_158),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_333),
.B(n_339),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_207),
.B(n_332),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_200),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_163),
.B(n_200),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_181),
.C(n_183),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_164),
.A2(n_165),
.B1(n_181),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_175),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_171),
.C(n_175),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_176),
.B(n_179),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_181),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_183),
.B(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_190),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_186),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_190),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_194),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_199),
.A2(n_297),
.B(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_202),
.B(n_203),
.C(n_206),
.Y(n_338)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_239),
.B(n_326),
.C(n_331),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_233),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_233),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_224),
.C(n_225),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_210),
.A2(n_211),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_220),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_216),
.C(n_220),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_224),
.B(n_225),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.C(n_230),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_320),
.B(n_325),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_273),
.B(n_319),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_262),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_244),
.B(n_262),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_255),
.C(n_259),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_245),
.B(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_248),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B(n_253),
.Y(n_248)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_253),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_254),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_255),
.A2(n_259),
.B1(n_260),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_267),
.B2(n_268),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_263),
.B(n_269),
.C(n_270),
.Y(n_324)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_313),
.B(n_318),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_293),
.B(n_312),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_287),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_287),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_317)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_301),
.B(n_311),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_299),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_299),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_306),
.B(n_310),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_304),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_317),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_324),
.Y(n_325)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_338),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_338),
.Y(n_339)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_345),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_353),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_349),
.B1(n_351),
.B2(n_352),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_347),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_349),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_351),
.C(n_353),
.Y(n_356)
);


endmodule