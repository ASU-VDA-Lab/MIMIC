module real_jpeg_15457_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_566),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_0),
.B(n_567),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_1),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_1),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_2),
.A2(n_9),
.B1(n_47),
.B2(n_51),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_2),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_2),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_2),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_2),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_2),
.B(n_73),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_2),
.B(n_336),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_2),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_2),
.B(n_384),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_3),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_3),
.Y(n_281)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_3),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_4),
.B(n_67),
.Y(n_66)
);

AND2x4_ASAP7_75t_SL g82 ( 
.A(n_4),
.B(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_4),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_4),
.B(n_140),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_4),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_4),
.B(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_4),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_4),
.B(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_5),
.Y(n_123)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_5),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_5),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_5),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_6),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_6),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_6),
.B(n_73),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_6),
.B(n_496),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_6),
.B(n_510),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_7),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_7),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_7),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_7),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_7),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_7),
.B(n_513),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_7),
.B(n_560),
.Y(n_559)
);

NAND2x1_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_8),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_8),
.B(n_85),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_8),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_8),
.B(n_78),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_8),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_8),
.B(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_9),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_9),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_9),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_9),
.B(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_9),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_9),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_9),
.B(n_481),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_9),
.B(n_520),
.Y(n_519)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_10),
.Y(n_193)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_11),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_12),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_12),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_12),
.B(n_126),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_12),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_12),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_12),
.B(n_143),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_12),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_12),
.B(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_13),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_13),
.Y(n_246)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_13),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_14),
.Y(n_141)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_14),
.Y(n_208)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_14),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_15),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_15),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_15),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_15),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_15),
.B(n_205),
.Y(n_378)
);

BUFx2_ASAP7_75t_R g398 ( 
.A(n_15),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_17),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_17),
.B(n_75),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_17),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_17),
.B(n_47),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_17),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_17),
.B(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g117 ( 
.A(n_18),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g522 ( 
.A(n_18),
.Y(n_522)
);

BUFx5_ASAP7_75t_L g562 ( 
.A(n_18),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_549),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_436),
.B(n_544),
.Y(n_22)
);

AO21x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_265),
.B(n_433),
.Y(n_23)
);

NOR2xp67_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_216),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_172),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_26),
.B(n_172),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_95),
.Y(n_26)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_27),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_70),
.C(n_87),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_29),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_45),
.C(n_56),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_30),
.B(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

MAJx2_ASAP7_75t_L g461 ( 
.A(n_31),
.B(n_166),
.C(n_258),
.Y(n_461)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_33),
.B(n_38),
.C(n_41),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_33),
.B(n_166),
.Y(n_255)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_36),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_40),
.Y(n_405)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_44),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_45),
.A2(n_46),
.B1(n_56),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_46),
.A2(n_284),
.B(n_288),
.Y(n_283)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_53),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_55),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_55),
.Y(n_229)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_56),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.C(n_66),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_58),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_57),
.A2(n_58),
.B1(n_66),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_58),
.B(n_100),
.C(n_107),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_62),
.B(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_66),
.Y(n_187)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_69),
.Y(n_274)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_69),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_70),
.A2(n_87),
.B1(n_88),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_70),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_81),
.C(n_83),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_71),
.B(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.C(n_77),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_72),
.A2(n_77),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_72),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_72),
.B(n_331),
.Y(n_330)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_74),
.B(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_77),
.Y(n_296)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_79),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_83),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_86),
.Y(n_287)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_86),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2x1_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_90),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_90),
.B(n_271),
.C(n_277),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_90),
.A2(n_162),
.B1(n_277),
.B2(n_278),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_94),
.B(n_161),
.C(n_162),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_131),
.B1(n_170),
.B2(n_171),
.Y(n_95)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_96),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_112),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_97),
.B(n_113),
.C(n_119),
.Y(n_261)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_106),
.B1(n_107),
.B2(n_111),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_100),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_100),
.A2(n_111),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_101),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_101),
.B(n_557),
.Y(n_556)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_105),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_107),
.B1(n_118),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_114),
.C(n_118),
.Y(n_113)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_111),
.B(n_222),
.C(n_232),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_119),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_120),
.B(n_125),
.C(n_128),
.Y(n_238)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_159),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_132),
.B(n_160),
.C(n_163),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.C(n_151),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_136),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.C(n_147),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_137),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_142),
.A2(n_147),
.B1(n_148),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_147),
.B(n_304),
.C(n_307),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_147),
.A2(n_148),
.B1(n_304),
.B2(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_149),
.Y(n_334)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_154),
.C(n_158),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_157),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_164),
.B(n_169),
.C(n_260),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_166),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_170),
.B(n_263),
.C(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_178),
.C(n_181),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_178),
.Y(n_324)
);

XOR2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_182),
.B(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_209),
.C(n_213),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_183),
.B(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_198),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_185),
.B(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_188),
.B(n_198),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_189),
.B(n_195),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.C(n_204),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_199),
.A2(n_203),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_199),
.Y(n_300)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_203),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_203),
.B(n_375),
.C(n_377),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_203),
.A2(n_301),
.B1(n_377),
.B2(n_378),
.Y(n_388)
);

XOR2x1_ASAP7_75t_L g298 ( 
.A(n_204),
.B(n_299),
.Y(n_298)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_210),
.B(n_213),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_216),
.A2(n_434),
.B(n_435),
.Y(n_433)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_262),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_217),
.B(n_262),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_218),
.B(n_220),
.C(n_252),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_252),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_237),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_221),
.B(n_238),
.C(n_239),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_231),
.A2(n_232),
.B1(n_465),
.B2(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_SL g487 ( 
.A(n_232),
.B(n_465),
.C(n_467),
.Y(n_487)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_240),
.B(n_242),
.C(n_247),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_247),
.Y(n_241)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_261),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_259),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_254),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_256),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_259),
.B(n_537),
.C(n_538),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_261),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_429),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_320),
.C(n_325),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_312),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_268),
.B(n_312),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_297),
.C(n_310),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_269),
.B(n_427),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_282),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_270),
.B(n_283),
.C(n_293),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_271),
.B(n_419),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

XNOR2x1_ASAP7_75t_SL g364 ( 
.A(n_272),
.B(n_275),
.Y(n_364)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_272),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_272),
.A2(n_382),
.B1(n_383),
.B2(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_293),
.Y(n_282)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_287),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_295),
.B(n_332),
.C(n_335),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_297),
.B(n_310),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_302),
.C(n_308),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_298),
.B(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_303),
.B(n_309),
.Y(n_414)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_304),
.Y(n_360)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_306),
.Y(n_452)
);

XOR2x2_ASAP7_75t_SL g358 ( 
.A(n_307),
.B(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_318),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_315),
.C(n_318),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_321),
.Y(n_431)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_322),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_424),
.B(n_428),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_410),
.B(n_423),
.Y(n_326)
);

OAI21x1_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_369),
.B(n_409),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_355),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_329),
.B(n_355),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_339),
.C(n_346),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_339),
.A2(n_340),
.B1(n_346),
.B2(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_341),
.B(n_345),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

AO22x1_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_350),
.B1(n_353),
.B2(n_354),
.Y(n_346)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_350),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_353),
.Y(n_362)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_351),
.Y(n_385)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_402),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_361),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_358),
.C(n_361),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_364),
.C(n_365),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_379),
.B(n_408),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_374),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_374),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_375),
.A2(n_376),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_380),
.A2(n_389),
.B(n_407),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_386),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_386),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_401),
.B(n_406),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_399),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_399),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_398),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_398),
.B(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_422),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_422),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_415),
.B2(n_416),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_417),
.C(n_421),
.Y(n_425)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_420),
.B2(n_421),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_425),
.B(n_426),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.C(n_432),
.Y(n_429)
);

NOR3xp33_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_525),
.C(n_539),
.Y(n_436)
);

OAI21x1_ASAP7_75t_SL g544 ( 
.A1(n_437),
.A2(n_545),
.B(n_548),
.Y(n_544)
);

NOR2x1_ASAP7_75t_R g437 ( 
.A(n_438),
.B(n_501),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_438),
.B(n_501),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_462),
.C(n_475),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_439),
.B(n_528),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_442),
.C(n_461),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_441),
.B(n_533),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_442),
.B(n_461),
.Y(n_533)
);

XNOR2x1_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_448),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_453),
.C(n_460),
.Y(n_478)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx6_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_447),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_453),
.B1(n_454),
.B2(n_460),
.Y(n_448)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_449),
.Y(n_460)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_459),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_462),
.A2(n_475),
.B1(n_476),
.B2(n_529),
.Y(n_528)
);

INVxp33_ASAP7_75t_SL g529 ( 
.A(n_462),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_473),
.C(n_474),
.Y(n_462)
);

XNOR2x2_ASAP7_75t_L g534 ( 
.A(n_463),
.B(n_535),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_467),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_465),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_465),
.A2(n_466),
.B1(n_495),
.B2(n_500),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_466),
.B(n_489),
.C(n_495),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_471),
.Y(n_516)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_471),
.Y(n_557)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_473),
.B(n_474),
.Y(n_535)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_486),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_477),
.B(n_487),
.C(n_488),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_478),
.B(n_480),
.C(n_483),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_483),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

XOR2x2_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_494),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_495),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_495),
.A2(n_500),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_495),
.B(n_509),
.C(n_512),
.Y(n_553)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_524),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_504),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_503),
.B(n_504),
.C(n_524),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_506),
.B1(n_517),
.B2(n_518),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_505),
.B(n_519),
.C(n_523),
.Y(n_563)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_512),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_508),
.A2(n_509),
.B1(n_556),
.B2(n_558),
.Y(n_555)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_519),
.B(n_523),
.Y(n_518)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

AOI21x1_ASAP7_75t_L g545 ( 
.A1(n_526),
.A2(n_546),
.B(n_547),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_530),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_SL g547 ( 
.A(n_527),
.B(n_530),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_534),
.C(n_536),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_531),
.A2(n_532),
.B1(n_534),
.B2(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_534),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_536),
.B(n_542),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_541),
.Y(n_539)
);

NOR2x1_ASAP7_75t_L g546 ( 
.A(n_540),
.B(n_541),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_565),
.Y(n_549)
);

NAND2x1_ASAP7_75t_SL g550 ( 
.A(n_551),
.B(n_564),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_551),
.B(n_564),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_563),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_554),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_559),
.Y(n_554)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_556),
.Y(n_558)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx8_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);


endmodule