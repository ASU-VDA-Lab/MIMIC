module fake_jpeg_8957_n_174 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_29),
.B1(n_27),
.B2(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_16),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_39),
.B(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_36),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_30),
.B1(n_29),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_34),
.B1(n_31),
.B2(n_18),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_19),
.Y(n_58)
);

CKINVDCx10_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

HAxp5_ASAP7_75t_SL g88 ( 
.A(n_56),
.B(n_72),
.CON(n_88),
.SN(n_88)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_22),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_37),
.C(n_36),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_48),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_22),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_18),
.Y(n_86)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_80),
.B(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_82),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_93),
.Y(n_107)
);

XOR2x1_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_58),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_97),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_64),
.B(n_62),
.CI(n_68),
.CON(n_96),
.SN(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_69),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_31),
.B(n_34),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_75),
.B(n_18),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_110),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_87),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_77),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_115),
.C(n_117),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_62),
.B1(n_44),
.B2(n_43),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_108),
.B1(n_114),
.B2(n_94),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_100),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_44),
.B1(n_74),
.B2(n_66),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_76),
.B1(n_66),
.B2(n_75),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_11),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_26),
.Y(n_116)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_1),
.Y(n_117)
);

NAND2x1_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_88),
.Y(n_120)
);

AOI21x1_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_127),
.B(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_114),
.A2(n_87),
.B1(n_96),
.B2(n_97),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_132),
.B1(n_92),
.B2(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_80),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_84),
.B1(n_89),
.B2(n_91),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_89),
.C(n_83),
.Y(n_134)
);

OAI221xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_91),
.B1(n_83),
.B2(n_24),
.C(n_105),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_118),
.C(n_103),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_138),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_113),
.B(n_86),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_117),
.C(n_84),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_144),
.Y(n_153)
);

AOI321xp33_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_145),
.A3(n_28),
.B1(n_21),
.B2(n_17),
.C(n_19),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_1),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_92),
.C(n_108),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_120),
.B1(n_122),
.B2(n_129),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_126),
.B1(n_123),
.B2(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_121),
.B1(n_125),
.B2(n_124),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_128),
.B1(n_20),
.B2(n_19),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_152),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_139),
.Y(n_157)
);

NOR2xp67_ASAP7_75t_R g159 ( 
.A(n_151),
.B(n_28),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_10),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_21),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_17),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_159),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_9),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_12),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_166),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_155),
.C(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_155),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_162),
.A3(n_150),
.B1(n_159),
.B2(n_153),
.C1(n_156),
.C2(n_20),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_170),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_165),
.A3(n_166),
.B1(n_153),
.B2(n_14),
.C1(n_12),
.C2(n_2),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_3),
.B(n_4),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_8),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_171),
.Y(n_174)
);


endmodule