module fake_jpeg_26311_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_21),
.B1(n_28),
.B2(n_24),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_16),
.B1(n_17),
.B2(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_30),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_32),
.C(n_20),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_55),
.Y(n_74)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_30),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_31),
.B(n_27),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_28),
.B1(n_21),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_23),
.B1(n_21),
.B2(n_28),
.Y(n_63)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_32),
.C(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_23),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_21),
.B1(n_28),
.B2(n_23),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_60),
.A2(n_53),
.B(n_45),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_68),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_24),
.B(n_25),
.C(n_27),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_81),
.B1(n_55),
.B2(n_44),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_79),
.B1(n_46),
.B2(n_59),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_23),
.B1(n_20),
.B2(n_32),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_80),
.B1(n_59),
.B2(n_53),
.Y(n_94)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_71),
.Y(n_92)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_83),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_26),
.A3(n_17),
.B1(n_31),
.B2(n_18),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_38),
.B1(n_26),
.B2(n_31),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_42),
.A2(n_32),
.B1(n_20),
.B2(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_18),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_51),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_51),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_59),
.B1(n_53),
.B2(n_46),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_97),
.B1(n_60),
.B2(n_81),
.Y(n_118)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_104),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_109),
.Y(n_131)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_108),
.Y(n_117)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_29),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_72),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_75),
.B(n_84),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_111),
.A2(n_124),
.B(n_3),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_128),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_78),
.B1(n_80),
.B2(n_63),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_123),
.B1(n_126),
.B2(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_122),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_79),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_71),
.B1(n_67),
.B2(n_77),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_97),
.A2(n_62),
.B1(n_73),
.B2(n_45),
.Y(n_126)
);

AO21x2_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_73),
.B(n_54),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_22),
.B(n_1),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_85),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_29),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_29),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_51),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_134),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_51),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_98),
.Y(n_154)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_120),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_133),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_125),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_127),
.B(n_96),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_115),
.B(n_121),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_143),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_148),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_96),
.B1(n_102),
.B2(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_109),
.C(n_104),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_155),
.C(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_103),
.C(n_54),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_22),
.C(n_1),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_0),
.C(n_1),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_111),
.C(n_123),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_160),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_127),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_2),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_119),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_158),
.C(n_157),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_117),
.B(n_115),
.C(n_126),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_175),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_132),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_181),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_183),
.C(n_146),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_156),
.B(n_147),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_184),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_118),
.C(n_134),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_5),
.C(n_6),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

OA21x2_ASAP7_75t_SL g197 ( 
.A1(n_180),
.A2(n_139),
.B(n_138),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_136),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_112),
.Y(n_182)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

XOR2x2_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_112),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

OAI322xp33_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_161),
.A3(n_162),
.B1(n_151),
.B2(n_153),
.C1(n_154),
.C2(n_143),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_197),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_142),
.B1(n_148),
.B2(n_150),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_186),
.A2(n_169),
.B1(n_173),
.B2(n_171),
.Y(n_204)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_201),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_160),
.B1(n_145),
.B2(n_140),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_191),
.A2(n_194),
.B1(n_196),
.B2(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

NAND2x1_ASAP7_75t_SL g194 ( 
.A(n_183),
.B(n_176),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_153),
.B1(n_159),
.B2(n_156),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_146),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_178),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_164),
.B1(n_166),
.B2(n_176),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_208),
.B1(n_190),
.B2(n_189),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_212),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_186),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_210),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_169),
.B1(n_166),
.B2(n_175),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_172),
.B1(n_167),
.B2(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_201),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_168),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_216),
.A2(n_224),
.B1(n_194),
.B2(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_198),
.C(n_188),
.Y(n_218)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_6),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_199),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_223),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_188),
.C(n_181),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_203),
.B(n_187),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_215),
.C(n_200),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_227),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_215),
.C(n_167),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_192),
.B(n_187),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_223),
.B(n_8),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_7),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_232),
.A2(n_216),
.B(n_220),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_234),
.A2(n_238),
.B(n_231),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_224),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_237),
.C(n_12),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_7),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_242),
.B(n_235),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_243),
.B(n_244),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_15),
.C(n_12),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_13),
.B(n_15),
.Y(n_247)
);


endmodule