module fake_jpeg_18830_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_29),
.B1(n_27),
.B2(n_25),
.Y(n_47)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_27),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_29),
.B1(n_33),
.B2(n_31),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_50),
.B1(n_36),
.B2(n_29),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_55),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_29),
.B1(n_31),
.B2(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_20),
.B1(n_21),
.B2(n_30),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_16),
.B1(n_19),
.B2(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_85),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_79),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_40),
.B1(n_36),
.B2(n_38),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_88),
.B1(n_59),
.B2(n_38),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_66),
.B(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_86),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_87),
.B1(n_59),
.B2(n_48),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_39),
.B(n_36),
.C(n_20),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_55),
.B(n_37),
.C(n_41),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_27),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_80),
.B1(n_83),
.B2(n_89),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_39),
.C(n_41),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_76),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_23),
.B1(n_21),
.B2(n_30),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_22),
.B(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_27),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_16),
.B1(n_19),
.B2(n_32),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_35),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_35),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_41),
.B1(n_38),
.B2(n_35),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_21),
.B(n_23),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_31),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_25),
.B(n_22),
.Y(n_135)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_110),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_111),
.B1(n_119),
.B2(n_45),
.Y(n_136)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_108),
.Y(n_142)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_114),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_38),
.B1(n_41),
.B2(n_45),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_73),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_37),
.B(n_54),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_17),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_17),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_117),
.B(n_77),
.Y(n_125)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_110),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_62),
.A2(n_41),
.B1(n_45),
.B2(n_23),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_68),
.C(n_74),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_129),
.C(n_111),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_123),
.B(n_25),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_125),
.B(n_24),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_63),
.B1(n_77),
.B2(n_76),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_127),
.B1(n_133),
.B2(n_102),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_75),
.B1(n_83),
.B2(n_80),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_73),
.C(n_80),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_119),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_83),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_25),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_87),
.B1(n_85),
.B2(n_78),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_137),
.B(n_92),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_143),
.B1(n_114),
.B2(n_98),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_0),
.B(n_1),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_140),
.B(n_144),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_41),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_87),
.B1(n_67),
.B2(n_30),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_94),
.A2(n_60),
.B1(n_32),
.B2(n_28),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_148),
.B1(n_24),
.B2(n_28),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_18),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_147),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_93),
.A2(n_60),
.B1(n_28),
.B2(n_24),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_145),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_149),
.B(n_150),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_155),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_93),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_153),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_91),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_97),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_163),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_114),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_161),
.B(n_168),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_147),
.C(n_140),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_113),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_166),
.B1(n_140),
.B2(n_122),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_99),
.B1(n_100),
.B2(n_96),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_137),
.B1(n_143),
.B2(n_122),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_17),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_170),
.B(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_17),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_173),
.B(n_179),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_101),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_176),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_25),
.B(n_101),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_178),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_18),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_109),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_135),
.Y(n_191)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_188),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_172),
.C(n_173),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_147),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_162),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_197),
.B1(n_204),
.B2(n_205),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_168),
.B1(n_174),
.B2(n_160),
.Y(n_215)
);

BUFx12_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_128),
.Y(n_201)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_138),
.B1(n_135),
.B2(n_98),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_166),
.A2(n_178),
.B1(n_163),
.B2(n_157),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_104),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_209),
.A2(n_169),
.B(n_152),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_216),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_213),
.B(n_224),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_192),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_218),
.C(n_221),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_227),
.Y(n_240)
);

FAx1_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_165),
.CI(n_174),
.CON(n_216),
.SN(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_167),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_203),
.B1(n_209),
.B2(n_187),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_226),
.B1(n_206),
.B2(n_184),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_169),
.B(n_176),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_223),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_155),
.B1(n_154),
.B2(n_104),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_25),
.B(n_7),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_37),
.C(n_70),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_229),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_198),
.B(n_11),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_196),
.B(n_11),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_232),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_37),
.C(n_26),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_247),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_243),
.Y(n_253)
);

OAI322xp33_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_189),
.A3(n_194),
.B1(n_200),
.B2(n_210),
.C1(n_207),
.C2(n_199),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_197),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_212),
.B(n_211),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_188),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_188),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_214),
.C(n_221),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_256),
.C(n_258),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_228),
.C(n_224),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_240),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_232),
.C(n_210),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_223),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_216),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_202),
.C(n_195),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_248),
.C(n_242),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_199),
.B(n_182),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_241),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_264),
.A2(n_245),
.B1(n_237),
.B2(n_234),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_274),
.B1(n_5),
.B2(n_15),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_271),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_233),
.B(n_245),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_272),
.A2(n_6),
.B(n_15),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_235),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_277),
.Y(n_284)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_18),
.B(n_6),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_L g281 ( 
.A1(n_276),
.A2(n_14),
.B(n_15),
.Y(n_281)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_8),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_262),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_274),
.B1(n_8),
.B2(n_2),
.Y(n_291)
);

OAI321xp33_ASAP7_75t_L g282 ( 
.A1(n_279),
.A2(n_255),
.A3(n_266),
.B1(n_254),
.B2(n_256),
.C(n_26),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_286),
.B(n_289),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_252),
.C(n_26),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_267),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_6),
.B(n_13),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_18),
.B(n_4),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_291),
.B(n_292),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_268),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_37),
.A3(n_2),
.B1(n_3),
.B2(n_8),
.C1(n_12),
.C2(n_1),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_4),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_3),
.B(n_12),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_37),
.C(n_2),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_0),
.B(n_1),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g299 ( 
.A1(n_297),
.A2(n_287),
.B(n_284),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.C(n_302),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_290),
.C(n_294),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_297),
.B(n_12),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_303),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_305),
.Y(n_308)
);


endmodule