module fake_ariane_1227_n_1441 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_155, n_127, n_1441);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_155;
input n_127;

output n_1441;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1432;
wire n_1108;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_1015;
wire n_545;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_368;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_1063;
wire n_537;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_329),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_124),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_343),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_326),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_184),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_339),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_43),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_299),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_312),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_131),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_3),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_230),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_277),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_157),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_345),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_247),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_170),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_274),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_186),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_328),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_34),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_325),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_117),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_324),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_259),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_177),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_76),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_102),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_129),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_135),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_207),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_327),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_19),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_218),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_165),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_262),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_111),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_78),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_32),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_59),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_65),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_348),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_140),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_163),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_61),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_69),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_166),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_293),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_346),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_87),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_313),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_56),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_106),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_179),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_161),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_14),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_244),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_290),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_104),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_148),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_110),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_96),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_307),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_279),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_266),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_126),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_227),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_205),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

BUFx10_ASAP7_75t_L g432 ( 
.A(n_203),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_62),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_337),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_99),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_209),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_27),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_316),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_159),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_318),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_50),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_206),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_67),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_267),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_347),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_304),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_134),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_238),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_25),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_211),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_340),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_197),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_26),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_281),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_223),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_229),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_19),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_202),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_14),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_248),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_17),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_322),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_228),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_225),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_94),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_200),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_79),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_198),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_46),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_193),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_66),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_239),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_146),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_214),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_39),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_317),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_344),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_25),
.Y(n_478)
);

BUFx5_ASAP7_75t_L g479 ( 
.A(n_201),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_112),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_119),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_30),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_75),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_168),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_70),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_199),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_53),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_137),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_74),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_153),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_176),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_152),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_255),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_121),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_265),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_351),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_92),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_204),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_257),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_303),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_308),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_349),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_50),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_174),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_41),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_63),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_242),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_354),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_296),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_149),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_28),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g512 ( 
.A(n_355),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_8),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_332),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_331),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_93),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_132),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_1),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_272),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_20),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_158),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_68),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_192),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_12),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_309),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_323),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_150),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_40),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_160),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_71),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_182),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_188),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_352),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_320),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_213),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_103),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_342),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_85),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_273),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_212),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_275),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_295),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_123),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_36),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_73),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_284),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_233),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_172),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_130),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_151),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_84),
.Y(n_551)
);

BUFx10_ASAP7_75t_L g552 ( 
.A(n_38),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_54),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_95),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_1),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_53),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_311),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_16),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_217),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_401),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_414),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_418),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_461),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_461),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_478),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_367),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_372),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_373),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_379),
.B(n_413),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_412),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_449),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_459),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_396),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_528),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_427),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_555),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_497),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_526),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_369),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_395),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_380),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_416),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_423),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_439),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_374),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_527),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_529),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_374),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_432),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_372),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_437),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_432),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_512),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_450),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_441),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_453),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_512),
.Y(n_597)
);

INVxp33_ASAP7_75t_SL g598 ( 
.A(n_457),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_359),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_450),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_470),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_475),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_487),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_503),
.Y(n_604)
);

CKINVDCx16_ASAP7_75t_R g605 ( 
.A(n_394),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_470),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_442),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_417),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_552),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_508),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_552),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_508),
.Y(n_612)
);

INVxp33_ASAP7_75t_SL g613 ( 
.A(n_505),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_511),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_513),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_546),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_518),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_546),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_362),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_364),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_365),
.B(n_0),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_370),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_520),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_396),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_375),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_524),
.Y(n_626)
);

NOR2xp67_ASAP7_75t_L g627 ( 
.A(n_544),
.B(n_0),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_426),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_382),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_553),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_384),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_556),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_558),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_361),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_387),
.B(n_2),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_389),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_363),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_391),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_366),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_426),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_410),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_411),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_523),
.Y(n_643)
);

BUFx2_ASAP7_75t_SL g644 ( 
.A(n_523),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_531),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_531),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_429),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_383),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_469),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_482),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_431),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_438),
.B(n_443),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_446),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_425),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_368),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_371),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_377),
.Y(n_657)
);

INVxp33_ASAP7_75t_SL g658 ( 
.A(n_378),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_381),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_385),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_392),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_565),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_645),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_645),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_585),
.B(n_417),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_568),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_654),
.B(n_448),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_560),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_561),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_577),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_649),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_648),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_608),
.B(n_455),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_562),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_585),
.B(n_360),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_573),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_591),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_571),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_573),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_644),
.B(n_462),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_572),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_569),
.B(n_376),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_634),
.B(n_376),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_619),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_574),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_576),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_620),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_622),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_578),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_625),
.Y(n_690)
);

INVxp67_ASAP7_75t_SL g691 ( 
.A(n_652),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_629),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_605),
.B(n_398),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_631),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_636),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_565),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_638),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_641),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_642),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_647),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_651),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_586),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_653),
.B(n_386),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_566),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_621),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_635),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_579),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_581),
.A2(n_476),
.B(n_464),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_563),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_587),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_582),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_583),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_570),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_575),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_R g715 ( 
.A(n_637),
.B(n_639),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_580),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_633),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_655),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_588),
.Y(n_719)
);

NOR2xp67_ASAP7_75t_L g720 ( 
.A(n_609),
.B(n_390),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_617),
.B(n_458),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_657),
.B(n_661),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_584),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_589),
.Y(n_724)
);

INVx5_ASAP7_75t_L g725 ( 
.A(n_658),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_592),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_594),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_595),
.B(n_509),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_600),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_601),
.Y(n_730)
);

OA21x2_ASAP7_75t_L g731 ( 
.A1(n_627),
.A2(n_483),
.B(n_481),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_596),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_606),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_610),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_612),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_616),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_656),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_618),
.B(n_485),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_624),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_628),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_602),
.B(n_488),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_640),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_643),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_656),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_659),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_646),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_603),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_676),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_668),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_669),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_674),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_663),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_676),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_676),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_691),
.B(n_598),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_676),
.Y(n_756)
);

BUFx4f_ASAP7_75t_L g757 ( 
.A(n_729),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_662),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_679),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_678),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_747),
.B(n_613),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_663),
.Y(n_762)
);

AO21x2_ASAP7_75t_L g763 ( 
.A1(n_708),
.A2(n_496),
.B(n_495),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_675),
.B(n_563),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_711),
.B(n_564),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_711),
.B(n_564),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_672),
.B(n_693),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_681),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_664),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_662),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_SL g771 ( 
.A(n_715),
.B(n_659),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_SL g772 ( 
.A1(n_683),
.A2(n_515),
.B1(n_519),
.B2(n_506),
.Y(n_772)
);

INVx3_ASAP7_75t_R g773 ( 
.A(n_742),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_682),
.A2(n_597),
.B1(n_593),
.B2(n_660),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_672),
.B(n_604),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_712),
.B(n_660),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_685),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_705),
.B(n_665),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_664),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_686),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_705),
.B(n_522),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_682),
.A2(n_388),
.B1(n_404),
.B2(n_386),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_704),
.B(n_614),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_679),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_684),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_728),
.B(n_615),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_684),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_721),
.B(n_623),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_679),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_671),
.B(n_626),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_706),
.B(n_525),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_699),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_699),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_718),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_679),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_700),
.Y(n_796)
);

AND2x6_ASAP7_75t_L g797 ( 
.A(n_747),
.B(n_388),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_666),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_700),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_688),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_716),
.B(n_630),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_670),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_690),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_692),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_682),
.B(n_532),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_713),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_682),
.B(n_550),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_682),
.B(n_404),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_696),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_739),
.B(n_567),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_689),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_695),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_687),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_702),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_722),
.B(n_632),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_687),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_683),
.A2(n_607),
.B1(n_599),
.B2(n_650),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_715),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_694),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_694),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_729),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_732),
.B(n_393),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_SL g823 ( 
.A(n_741),
.B(n_530),
.C(n_521),
.Y(n_823)
);

AND2x6_ASAP7_75t_L g824 ( 
.A(n_703),
.B(n_408),
.Y(n_824)
);

BUFx10_ASAP7_75t_L g825 ( 
.A(n_710),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_697),
.Y(n_826)
);

INVx5_ASAP7_75t_L g827 ( 
.A(n_729),
.Y(n_827)
);

BUFx10_ASAP7_75t_L g828 ( 
.A(n_745),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_667),
.B(n_567),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_698),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_701),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_714),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_725),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_732),
.B(n_397),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_719),
.B(n_590),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_725),
.B(n_399),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_729),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_730),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_833),
.B(n_725),
.Y(n_839)
);

AND2x6_ASAP7_75t_SL g840 ( 
.A(n_810),
.B(n_717),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_L g841 ( 
.A(n_818),
.B(n_725),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_815),
.B(n_673),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_778),
.B(n_719),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_778),
.B(n_731),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_752),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_748),
.Y(n_846)
);

O2A1O1Ixp5_ASAP7_75t_L g847 ( 
.A1(n_781),
.A2(n_727),
.B(n_733),
.C(n_726),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_749),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_788),
.B(n_677),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_791),
.A2(n_724),
.B1(n_738),
.B2(n_677),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_767),
.B(n_742),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_755),
.A2(n_724),
.B1(n_730),
.B2(n_734),
.Y(n_852)
);

NAND2x1_ASAP7_75t_L g853 ( 
.A(n_795),
.B(n_731),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_816),
.B(n_680),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_782),
.A2(n_731),
.B1(n_712),
.B2(n_723),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_761),
.B(n_730),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_829),
.B(n_740),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_SL g858 ( 
.A(n_794),
.B(n_737),
.Y(n_858)
);

NOR3xp33_ASAP7_75t_L g859 ( 
.A(n_783),
.B(n_744),
.C(n_737),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_L g860 ( 
.A(n_835),
.B(n_730),
.C(n_738),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_816),
.B(n_735),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_791),
.B(n_736),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_781),
.B(n_703),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_762),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_775),
.B(n_743),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_750),
.B(n_751),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_760),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_801),
.B(n_720),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_768),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_777),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_782),
.A2(n_772),
.B1(n_823),
.B2(n_824),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_832),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_780),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_L g874 ( 
.A(n_771),
.B(n_744),
.C(n_746),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_800),
.B(n_703),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_776),
.B(n_723),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_803),
.B(n_707),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_757),
.B(n_707),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_804),
.B(n_543),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_SL g880 ( 
.A(n_802),
.B(n_590),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_757),
.B(n_611),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_821),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_812),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_826),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_786),
.B(n_611),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_830),
.B(n_400),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_831),
.B(n_402),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_790),
.B(n_709),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_772),
.A2(n_823),
.B1(n_824),
.B2(n_807),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_822),
.A2(n_516),
.B(n_424),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_813),
.B(n_403),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_819),
.B(n_405),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_824),
.A2(n_421),
.B1(n_467),
.B2(n_408),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_834),
.A2(n_789),
.B(n_820),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_L g895 ( 
.A(n_811),
.B(n_406),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_764),
.B(n_709),
.Y(n_896)
);

BUFx12f_ASAP7_75t_L g897 ( 
.A(n_825),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_764),
.B(n_696),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_758),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_748),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_824),
.A2(n_409),
.B1(n_415),
.B2(n_407),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_773),
.B(n_419),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_776),
.B(n_420),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_785),
.B(n_422),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_787),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_792),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_765),
.B(n_428),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_805),
.A2(n_467),
.B(n_421),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_765),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_805),
.A2(n_504),
.B(n_474),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_793),
.B(n_430),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_796),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_807),
.A2(n_474),
.B1(n_510),
.B2(n_504),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_814),
.B(n_433),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_799),
.B(n_434),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_766),
.B(n_435),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_748),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_836),
.A2(n_510),
.B(n_4),
.C(n_2),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_766),
.B(n_436),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_769),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_779),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_SL g922 ( 
.A(n_798),
.B(n_440),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_808),
.A2(n_445),
.B(n_444),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_808),
.B(n_447),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_797),
.B(n_479),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_806),
.B(n_774),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_825),
.B(n_451),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_817),
.A2(n_454),
.B1(n_456),
.B2(n_452),
.Y(n_928)
);

NOR2x1p5_ASAP7_75t_L g929 ( 
.A(n_828),
.B(n_460),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_797),
.B(n_821),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_837),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_753),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_838),
.Y(n_933)
);

BUFx8_ASAP7_75t_L g934 ( 
.A(n_770),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_806),
.B(n_463),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_882),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_842),
.B(n_809),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_843),
.A2(n_763),
.B(n_754),
.Y(n_938)
);

NAND2xp33_ASAP7_75t_SL g939 ( 
.A(n_862),
.B(n_821),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_845),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_934),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_872),
.B(n_839),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_844),
.B(n_797),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_899),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_864),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_848),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_867),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_920),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_851),
.B(n_828),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_863),
.B(n_797),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_934),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_900),
.Y(n_952)
);

AND2x4_ASAP7_75t_SL g953 ( 
.A(n_839),
.B(n_810),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_882),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_869),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_921),
.Y(n_956)
);

INVx3_ASAP7_75t_SL g957 ( 
.A(n_849),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_844),
.B(n_827),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_876),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_909),
.B(n_827),
.Y(n_960)
);

INVxp67_ASAP7_75t_SL g961 ( 
.A(n_900),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_897),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_857),
.B(n_810),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_870),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_900),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_874),
.B(n_827),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_873),
.B(n_754),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_858),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_883),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_898),
.B(n_795),
.Y(n_970)
);

BUFx12f_ASAP7_75t_L g971 ( 
.A(n_840),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_905),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_846),
.Y(n_973)
);

NAND2xp33_ASAP7_75t_R g974 ( 
.A(n_888),
.B(n_784),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_865),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_871),
.A2(n_784),
.B1(n_756),
.B2(n_759),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_906),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_846),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_884),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_926),
.B(n_753),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_912),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_896),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_917),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_866),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_885),
.B(n_753),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_850),
.B(n_756),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_R g987 ( 
.A(n_841),
.B(n_756),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_877),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_850),
.A2(n_763),
.B1(n_759),
.B2(n_465),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_852),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_875),
.Y(n_991)
);

BUFx10_ASAP7_75t_L g992 ( 
.A(n_935),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_929),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_855),
.B(n_759),
.Y(n_994)
);

NAND2xp33_ASAP7_75t_SL g995 ( 
.A(n_927),
.B(n_559),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_854),
.B(n_466),
.Y(n_996)
);

BUFx4f_ASAP7_75t_L g997 ( 
.A(n_917),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_931),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_879),
.B(n_468),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_889),
.A2(n_860),
.B1(n_923),
.B2(n_922),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_932),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_R g1002 ( 
.A(n_880),
.B(n_471),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_933),
.Y(n_1003)
);

INVxp67_ASAP7_75t_SL g1004 ( 
.A(n_853),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_881),
.B(n_557),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_938),
.A2(n_847),
.B(n_923),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_958),
.A2(n_894),
.B(n_856),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_944),
.Y(n_1008)
);

BUFx2_ASAP7_75t_R g1009 ( 
.A(n_962),
.Y(n_1009)
);

O2A1O1Ixp5_ASAP7_75t_L g1010 ( 
.A1(n_986),
.A2(n_890),
.B(n_878),
.C(n_914),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_958),
.A2(n_930),
.B(n_910),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_975),
.B(n_903),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_984),
.B(n_908),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_937),
.B(n_907),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_943),
.A2(n_910),
.B(n_908),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_SL g1016 ( 
.A1(n_967),
.A2(n_918),
.B(n_861),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_959),
.B(n_916),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_946),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_942),
.B(n_859),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_947),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_942),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_982),
.B(n_919),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_1004),
.A2(n_924),
.B(n_887),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_996),
.A2(n_886),
.B(n_868),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_959),
.B(n_895),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_1000),
.A2(n_904),
.B(n_915),
.C(n_911),
.Y(n_1026)
);

BUFx4_ASAP7_75t_SL g1027 ( 
.A(n_941),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_955),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_991),
.B(n_963),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_943),
.A2(n_925),
.B(n_892),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_970),
.B(n_902),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_972),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_949),
.B(n_928),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_988),
.B(n_928),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_992),
.B(n_893),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_952),
.Y(n_1036)
);

OA21x2_ASAP7_75t_L g1037 ( 
.A1(n_994),
.A2(n_925),
.B(n_913),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_967),
.A2(n_891),
.B(n_901),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_SL g1039 ( 
.A1(n_966),
.A2(n_3),
.B(n_4),
.Y(n_1039)
);

OA21x2_ASAP7_75t_L g1040 ( 
.A1(n_994),
.A2(n_473),
.B(n_472),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_950),
.A2(n_479),
.B(n_64),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_990),
.B(n_964),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_969),
.B(n_479),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_980),
.A2(n_479),
.A3(n_498),
.B(n_425),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_979),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_977),
.Y(n_1046)
);

NOR2x1_ASAP7_75t_SL g1047 ( 
.A(n_970),
.B(n_425),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_976),
.A2(n_479),
.B(n_72),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_992),
.B(n_5),
.Y(n_1049)
);

INVx6_ASAP7_75t_L g1050 ( 
.A(n_971),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_951),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_952),
.Y(n_1052)
);

OA21x2_ASAP7_75t_L g1053 ( 
.A1(n_989),
.A2(n_480),
.B(n_477),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_952),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_981),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_1002),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_948),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_1003),
.A2(n_479),
.A3(n_498),
.B(n_425),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_953),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_985),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_968),
.B(n_484),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_968),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_999),
.B(n_5),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_973),
.A2(n_77),
.B(n_60),
.Y(n_1064)
);

O2A1O1Ixp5_ASAP7_75t_L g1065 ( 
.A1(n_939),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_997),
.B(n_498),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_965),
.Y(n_1067)
);

OA21x2_ASAP7_75t_L g1068 ( 
.A1(n_1006),
.A2(n_989),
.B(n_1000),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_1027),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1033),
.A2(n_956),
.B1(n_998),
.B2(n_1005),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1014),
.A2(n_974),
.B1(n_957),
.B2(n_970),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1032),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1046),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1023),
.A2(n_997),
.B(n_961),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1018),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1030),
.A2(n_983),
.B(n_973),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1055),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_SL g1078 ( 
.A1(n_1053),
.A2(n_993),
.B1(n_960),
.B2(n_966),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1020),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1028),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_1042),
.B(n_940),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1045),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1042),
.Y(n_1083)
);

OA21x2_ASAP7_75t_L g1084 ( 
.A1(n_1006),
.A2(n_945),
.B(n_960),
.Y(n_1084)
);

AO21x2_ASAP7_75t_L g1085 ( 
.A1(n_1007),
.A2(n_987),
.B(n_1001),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_1015),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_1021),
.B(n_936),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_1021),
.B(n_936),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1029),
.B(n_965),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1012),
.B(n_983),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_SL g1091 ( 
.A1(n_1016),
.A2(n_995),
.B(n_978),
.Y(n_1091)
);

OAI221xp5_ASAP7_75t_SL g1092 ( 
.A1(n_1022),
.A2(n_954),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1048),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1057),
.Y(n_1094)
);

AO31x2_ASAP7_75t_L g1095 ( 
.A1(n_1026),
.A2(n_1001),
.A3(n_978),
.B(n_965),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1043),
.Y(n_1096)
);

OA21x2_ASAP7_75t_L g1097 ( 
.A1(n_1038),
.A2(n_489),
.B(n_486),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1034),
.A2(n_954),
.B(n_978),
.C(n_1001),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1053),
.A2(n_498),
.B1(n_491),
.B2(n_492),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_1052),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1058),
.Y(n_1101)
);

AO21x1_ASAP7_75t_L g1102 ( 
.A1(n_1013),
.A2(n_6),
.B(n_9),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1052),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1064),
.A2(n_1010),
.B(n_1043),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1060),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_1008),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_1052),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1024),
.A2(n_493),
.B(n_490),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1063),
.A2(n_499),
.B(n_494),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_1067),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1013),
.A2(n_501),
.B(n_502),
.C(n_500),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1019),
.A2(n_514),
.B1(n_517),
.B2(n_507),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1058),
.Y(n_1113)
);

AO21x2_ASAP7_75t_L g1114 ( 
.A1(n_1047),
.A2(n_534),
.B(n_533),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1060),
.B(n_10),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_1067),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1039),
.A2(n_81),
.B(n_80),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_1056),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1062),
.B(n_11),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1017),
.A2(n_536),
.B1(n_537),
.B2(n_535),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1025),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1040),
.A2(n_83),
.B(n_82),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1067),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1031),
.A2(n_539),
.B(n_538),
.Y(n_1124)
);

OR2x6_ASAP7_75t_L g1125 ( 
.A(n_1098),
.B(n_1031),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1083),
.B(n_1062),
.Y(n_1126)
);

OR2x2_ASAP7_75t_L g1127 ( 
.A(n_1105),
.B(n_1049),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1106),
.B(n_1019),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1075),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1079),
.Y(n_1130)
);

OAI211xp5_ASAP7_75t_SL g1131 ( 
.A1(n_1090),
.A2(n_1065),
.B(n_1061),
.C(n_1035),
.Y(n_1131)
);

BUFx12f_ASAP7_75t_L g1132 ( 
.A(n_1069),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_1069),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1070),
.B(n_1051),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1118),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1072),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_1081),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1092),
.A2(n_1070),
.B1(n_1120),
.B2(n_1109),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1121),
.B(n_1059),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1072),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1115),
.B(n_1036),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1100),
.B(n_1116),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1071),
.A2(n_1050),
.B1(n_1066),
.B2(n_1054),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1100),
.Y(n_1144)
);

CKINVDCx11_ASAP7_75t_R g1145 ( 
.A(n_1116),
.Y(n_1145)
);

INVx4_ASAP7_75t_SL g1146 ( 
.A(n_1123),
.Y(n_1146)
);

AOI22x1_ASAP7_75t_L g1147 ( 
.A1(n_1091),
.A2(n_1036),
.B1(n_1054),
.B2(n_1009),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1099),
.A2(n_1040),
.B1(n_1037),
.B2(n_1050),
.Y(n_1148)
);

OAI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1119),
.A2(n_1037),
.B1(n_541),
.B2(n_542),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1123),
.Y(n_1150)
);

OAI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1112),
.A2(n_540),
.B1(n_545),
.B2(n_547),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1080),
.B(n_11),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_1087),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1082),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1098),
.B(n_548),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1073),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1073),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1068),
.A2(n_549),
.B1(n_551),
.B2(n_554),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1099),
.A2(n_1044),
.B1(n_1058),
.B2(n_15),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1077),
.B(n_1044),
.Y(n_1160)
);

AOI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_1097),
.A2(n_1044),
.B(n_12),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1108),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1078),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_1103),
.Y(n_1164)
);

CKINVDCx11_ASAP7_75t_R g1165 ( 
.A(n_1087),
.Y(n_1165)
);

NOR2x1_ASAP7_75t_SL g1166 ( 
.A(n_1089),
.B(n_18),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1103),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1074),
.A2(n_20),
.B(n_21),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1068),
.A2(n_21),
.B(n_22),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1068),
.A2(n_1097),
.B1(n_1120),
.B2(n_1102),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1096),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_1171)
);

AOI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1097),
.A2(n_88),
.B(n_86),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1111),
.A2(n_1089),
.B(n_1124),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_1087),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1077),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1094),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1084),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1107),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1084),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1101),
.A2(n_1113),
.A3(n_1111),
.B(n_1084),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1095),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1088),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1088),
.B(n_27),
.Y(n_1183)
);

AO21x2_ASAP7_75t_L g1184 ( 
.A1(n_1101),
.A2(n_90),
.B(n_89),
.Y(n_1184)
);

OAI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1138),
.A2(n_1107),
.B1(n_1110),
.B2(n_1088),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1150),
.Y(n_1186)
);

OAI211xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1128),
.A2(n_1086),
.B(n_1110),
.C(n_30),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1134),
.A2(n_1114),
.B1(n_1113),
.B2(n_1085),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1129),
.Y(n_1189)
);

OAI211xp5_ASAP7_75t_SL g1190 ( 
.A1(n_1133),
.A2(n_1086),
.B(n_29),
.C(n_31),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1158),
.A2(n_1114),
.B1(n_1085),
.B2(n_1122),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1162),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1158),
.A2(n_1117),
.B1(n_1076),
.B2(n_1104),
.Y(n_1193)
);

OA21x2_ASAP7_75t_L g1194 ( 
.A1(n_1161),
.A2(n_1093),
.B(n_1076),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1170),
.A2(n_1095),
.B1(n_33),
.B2(n_34),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1141),
.B(n_1095),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1130),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1170),
.A2(n_1095),
.B1(n_33),
.B2(n_35),
.Y(n_1198)
);

OAI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1143),
.A2(n_1125),
.B1(n_1182),
.B2(n_1127),
.Y(n_1199)
);

NAND2x1_ASAP7_75t_L g1200 ( 
.A(n_1125),
.B(n_32),
.Y(n_1200)
);

AO21x2_ASAP7_75t_L g1201 ( 
.A1(n_1160),
.A2(n_97),
.B(n_91),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1156),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1157),
.Y(n_1203)
);

OAI211xp5_ASAP7_75t_SL g1204 ( 
.A1(n_1171),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_1204)
);

AO21x2_ASAP7_75t_L g1205 ( 
.A1(n_1149),
.A2(n_100),
.B(n_98),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1154),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1126),
.B(n_37),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1137),
.B(n_38),
.Y(n_1208)
);

AOI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1169),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.C(n_42),
.Y(n_1209)
);

OAI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1143),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1176),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1163),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1175),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1136),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1125),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1164),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1137),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1131),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1173),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_1219)
);

OAI221xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1168),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.C(n_55),
.Y(n_1220)
);

INVx6_ASAP7_75t_L g1221 ( 
.A(n_1132),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1181),
.A2(n_235),
.A3(n_357),
.B(n_353),
.Y(n_1222)
);

AOI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1151),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.C(n_58),
.Y(n_1223)
);

INVx5_ASAP7_75t_SL g1224 ( 
.A(n_1142),
.Y(n_1224)
);

AOI221xp5_ASAP7_75t_L g1225 ( 
.A1(n_1152),
.A2(n_57),
.B1(n_58),
.B2(n_101),
.C(n_105),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1142),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1140),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1150),
.B(n_107),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1139),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1148),
.A2(n_1155),
.B1(n_1183),
.B2(n_1159),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1183),
.A2(n_108),
.B1(n_109),
.B2(n_113),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1177),
.Y(n_1232)
);

BUFx4f_ASAP7_75t_SL g1233 ( 
.A(n_1174),
.Y(n_1233)
);

AOI222xp33_ASAP7_75t_L g1234 ( 
.A1(n_1166),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.C1(n_118),
.C2(n_120),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1146),
.B(n_1144),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1145),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1179),
.Y(n_1237)
);

OAI211xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1165),
.A2(n_128),
.B(n_133),
.C(n_136),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_1224),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1200),
.A2(n_1172),
.B(n_1228),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1217),
.B(n_1180),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1189),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1235),
.Y(n_1243)
);

AND2x4_ASAP7_75t_SL g1244 ( 
.A(n_1235),
.B(n_1153),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1192),
.A2(n_1184),
.B1(n_1147),
.B2(n_1178),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1196),
.B(n_1180),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1237),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1197),
.B(n_1180),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1206),
.B(n_1167),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1211),
.B(n_1153),
.Y(n_1250)
);

OAI222xp33_ASAP7_75t_L g1251 ( 
.A1(n_1195),
.A2(n_1135),
.B1(n_1184),
.B2(n_1146),
.C1(n_142),
.C2(n_143),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1213),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1216),
.B(n_138),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1202),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1216),
.B(n_139),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1232),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1229),
.B(n_1203),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1214),
.Y(n_1258)
);

NAND2x1_ASAP7_75t_L g1259 ( 
.A(n_1186),
.B(n_1226),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1227),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1186),
.Y(n_1261)
);

INVx2_ASAP7_75t_R g1262 ( 
.A(n_1224),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1194),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1219),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_1264)
);

INVxp67_ASAP7_75t_SL g1265 ( 
.A(n_1199),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1194),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1224),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1207),
.B(n_147),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1208),
.B(n_154),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1198),
.B(n_155),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1188),
.B(n_156),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1201),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1222),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1228),
.B(n_162),
.Y(n_1274)
);

AND2x4_ASAP7_75t_SL g1275 ( 
.A(n_1230),
.B(n_164),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1201),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1193),
.B(n_167),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1185),
.B(n_358),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1220),
.A2(n_169),
.B1(n_171),
.B2(n_173),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1222),
.B(n_175),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1222),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1215),
.B(n_1210),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1191),
.B(n_178),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1258),
.Y(n_1284)
);

OAI211xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1282),
.A2(n_1223),
.B(n_1218),
.C(n_1209),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1257),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1265),
.A2(n_1192),
.B1(n_1212),
.B2(n_1231),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1257),
.Y(n_1288)
);

AOI31xp33_ASAP7_75t_L g1289 ( 
.A1(n_1253),
.A2(n_1234),
.A3(n_1231),
.B(n_1225),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1242),
.B(n_1252),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1261),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1279),
.A2(n_1190),
.B1(n_1204),
.B2(n_1187),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1254),
.Y(n_1293)
);

OAI221xp5_ASAP7_75t_L g1294 ( 
.A1(n_1245),
.A2(n_1269),
.B1(n_1234),
.B2(n_1270),
.C(n_1280),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1248),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1253),
.B(n_1238),
.C(n_1236),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1248),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1243),
.B(n_1205),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1249),
.B(n_1205),
.Y(n_1299)
);

AOI211xp5_ASAP7_75t_L g1300 ( 
.A1(n_1251),
.A2(n_1233),
.B(n_1221),
.C(n_183),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1243),
.B(n_1221),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1270),
.A2(n_180),
.B1(n_181),
.B2(n_185),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1277),
.A2(n_1275),
.B(n_1267),
.Y(n_1303)
);

AOI211xp5_ASAP7_75t_L g1304 ( 
.A1(n_1277),
.A2(n_1255),
.B(n_1264),
.C(n_1268),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1243),
.B(n_187),
.Y(n_1305)
);

AOI221xp5_ASAP7_75t_L g1306 ( 
.A1(n_1273),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.C(n_194),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1243),
.B(n_195),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1258),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1275),
.A2(n_196),
.B1(n_208),
.B2(n_210),
.Y(n_1309)
);

OAI211xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1263),
.A2(n_215),
.B(n_216),
.C(n_219),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1284),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1291),
.B(n_1249),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1290),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1286),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1295),
.B(n_1263),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1308),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1297),
.B(n_1266),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1288),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1293),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1299),
.B(n_1250),
.Y(n_1320)
);

AOI221x1_ASAP7_75t_L g1321 ( 
.A1(n_1287),
.A2(n_1278),
.B1(n_1255),
.B2(n_1260),
.C(n_1276),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1301),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1301),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1298),
.B(n_1241),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1298),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1294),
.B(n_1241),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1304),
.B(n_1266),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1303),
.B(n_1250),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1305),
.B(n_1267),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1322),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1324),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1328),
.B(n_1289),
.Y(n_1332)
);

NAND2x1_ASAP7_75t_L g1333 ( 
.A(n_1323),
.B(n_1267),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1324),
.Y(n_1334)
);

AOI21xp33_ASAP7_75t_L g1335 ( 
.A1(n_1326),
.A2(n_1300),
.B(n_1285),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1323),
.B(n_1322),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1319),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1323),
.B(n_1244),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1322),
.B(n_1320),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1327),
.B(n_1256),
.Y(n_1340)
);

NAND4xp25_ASAP7_75t_L g1341 ( 
.A(n_1332),
.B(n_1292),
.C(n_1321),
.D(n_1312),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1332),
.B(n_1327),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1337),
.B(n_1313),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1336),
.B(n_1329),
.Y(n_1344)
);

OR2x6_ASAP7_75t_L g1345 ( 
.A(n_1338),
.B(n_1268),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1335),
.A2(n_1326),
.B(n_1296),
.Y(n_1346)
);

NAND4xp25_ASAP7_75t_L g1347 ( 
.A(n_1335),
.B(n_1292),
.C(n_1302),
.D(n_1269),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1338),
.B(n_1329),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1331),
.B(n_1314),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1334),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1340),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1339),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1340),
.B(n_1318),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1346),
.A2(n_1333),
.B(n_1330),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1341),
.B(n_1315),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1343),
.Y(n_1356)
);

OAI32xp33_ASAP7_75t_L g1357 ( 
.A1(n_1342),
.A2(n_1325),
.A3(n_1274),
.B1(n_1318),
.B2(n_1280),
.Y(n_1357)
);

NOR3xp33_ASAP7_75t_L g1358 ( 
.A(n_1347),
.B(n_1310),
.C(n_1306),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1345),
.Y(n_1359)
);

OAI332xp33_ASAP7_75t_L g1360 ( 
.A1(n_1351),
.A2(n_1271),
.A3(n_1276),
.B1(n_1272),
.B2(n_1281),
.B3(n_1311),
.C1(n_1316),
.C2(n_1256),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1348),
.B(n_1329),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1345),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1356),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1355),
.B(n_1349),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1362),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1359),
.Y(n_1366)
);

NAND3xp33_ASAP7_75t_SL g1367 ( 
.A(n_1358),
.B(n_1352),
.C(n_1350),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1361),
.Y(n_1368)
);

OAI31xp33_ASAP7_75t_L g1369 ( 
.A1(n_1354),
.A2(n_1283),
.A3(n_1353),
.B(n_1271),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1368),
.B(n_1344),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1365),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1363),
.B(n_1357),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1366),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1364),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1367),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1369),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1375),
.B(n_1371),
.C(n_1373),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1371),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1374),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1370),
.Y(n_1380)
);

AND3x1_ASAP7_75t_L g1381 ( 
.A(n_1372),
.B(n_1369),
.C(n_1307),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1376),
.B(n_1315),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1371),
.B(n_1360),
.Y(n_1383)
);

NAND4xp25_ASAP7_75t_L g1384 ( 
.A(n_1374),
.B(n_1309),
.C(n_1305),
.D(n_1283),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1376),
.A2(n_1360),
.B(n_1281),
.C(n_1317),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1383),
.A2(n_1317),
.B1(n_1272),
.B2(n_1244),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1380),
.B(n_1259),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1379),
.B(n_1239),
.Y(n_1388)
);

XNOR2xp5_ASAP7_75t_L g1389 ( 
.A(n_1381),
.B(n_1240),
.Y(n_1389)
);

AOI222xp33_ASAP7_75t_L g1390 ( 
.A1(n_1377),
.A2(n_1385),
.B1(n_1378),
.B2(n_1382),
.C1(n_1384),
.C2(n_1246),
.Y(n_1390)
);

AOI221xp5_ASAP7_75t_L g1391 ( 
.A1(n_1383),
.A2(n_1316),
.B1(n_1311),
.B2(n_1246),
.C(n_1247),
.Y(n_1391)
);

NAND3xp33_ASAP7_75t_L g1392 ( 
.A(n_1377),
.B(n_1239),
.C(n_1247),
.Y(n_1392)
);

AOI211xp5_ASAP7_75t_L g1393 ( 
.A1(n_1377),
.A2(n_1262),
.B(n_1239),
.C(n_222),
.Y(n_1393)
);

AOI221xp5_ASAP7_75t_L g1394 ( 
.A1(n_1389),
.A2(n_1239),
.B1(n_1262),
.B2(n_224),
.C(n_226),
.Y(n_1394)
);

AOI221xp5_ASAP7_75t_L g1395 ( 
.A1(n_1391),
.A2(n_1239),
.B1(n_221),
.B2(n_231),
.C(n_232),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1387),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1388),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_R g1398 ( 
.A(n_1393),
.B(n_220),
.Y(n_1398)
);

INVx5_ASAP7_75t_L g1399 ( 
.A(n_1392),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1390),
.B(n_234),
.Y(n_1400)
);

BUFx12f_ASAP7_75t_L g1401 ( 
.A(n_1386),
.Y(n_1401)
);

AOI21xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1388),
.A2(n_236),
.B(n_237),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1396),
.B(n_240),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1397),
.B(n_241),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1399),
.B(n_243),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1399),
.B(n_245),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1400),
.B(n_246),
.C(n_249),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1401),
.B(n_250),
.Y(n_1408)
);

NOR2x1_ASAP7_75t_L g1409 ( 
.A(n_1398),
.B(n_251),
.Y(n_1409)
);

NAND4xp25_ASAP7_75t_L g1410 ( 
.A(n_1394),
.B(n_252),
.C(n_253),
.D(n_254),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1402),
.B(n_256),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_SL g1412 ( 
.A(n_1406),
.B(n_1395),
.C(n_260),
.Y(n_1412)
);

NAND3xp33_ASAP7_75t_L g1413 ( 
.A(n_1407),
.B(n_258),
.C(n_261),
.Y(n_1413)
);

OAI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_1405),
.A2(n_263),
.B1(n_264),
.B2(n_268),
.C(n_269),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1403),
.A2(n_270),
.B(n_271),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1404),
.B(n_276),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1409),
.A2(n_278),
.B1(n_280),
.B2(n_283),
.Y(n_1417)
);

OAI322xp33_ASAP7_75t_L g1418 ( 
.A1(n_1408),
.A2(n_285),
.A3(n_286),
.B1(n_287),
.B2(n_288),
.C1(n_289),
.C2(n_291),
.Y(n_1418)
);

NOR3xp33_ASAP7_75t_L g1419 ( 
.A(n_1410),
.B(n_292),
.C(n_294),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1411),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1420),
.B(n_1412),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1416),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1417),
.Y(n_1423)
);

OAI211xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1415),
.A2(n_297),
.B(n_298),
.C(n_300),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1413),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1421),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1422),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1423),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1425),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1426),
.B(n_1419),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1429),
.B(n_1428),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1431),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1430),
.B(n_1427),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1432),
.A2(n_1414),
.B(n_1424),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1433),
.A2(n_1418),
.B1(n_302),
.B2(n_305),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1434),
.Y(n_1436)
);

OR2x6_ASAP7_75t_L g1437 ( 
.A(n_1435),
.B(n_301),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1434),
.A2(n_306),
.B1(n_310),
.B2(n_314),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1436),
.A2(n_315),
.B1(n_321),
.B2(n_330),
.Y(n_1439)
);

OAI221xp5_ASAP7_75t_R g1440 ( 
.A1(n_1439),
.A2(n_1437),
.B1(n_1438),
.B2(n_335),
.C(n_336),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1440),
.A2(n_333),
.B1(n_334),
.B2(n_338),
.Y(n_1441)
);


endmodule