module fake_netlist_6_297_n_271 (n_41, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_49, n_7, n_30, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_31, n_25, n_40, n_44, n_271);

input n_41;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_49;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_31;
input n_25;
input n_40;
input n_44;

output n_271;

wire n_52;
wire n_119;
wire n_91;
wire n_163;
wire n_146;
wire n_235;
wire n_256;
wire n_193;
wire n_147;
wire n_269;
wire n_258;
wire n_154;
wire n_191;
wire n_88;
wire n_209;
wire n_98;
wire n_260;
wire n_265;
wire n_113;
wire n_63;
wire n_223;
wire n_270;
wire n_73;
wire n_148;
wire n_226;
wire n_138;
wire n_161;
wire n_208;
wire n_199;
wire n_68;
wire n_228;
wire n_252;
wire n_266;
wire n_166;
wire n_184;
wire n_212;
wire n_268;
wire n_50;
wire n_158;
wire n_216;
wire n_217;
wire n_83;
wire n_206;
wire n_210;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_227;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_204;
wire n_245;
wire n_87;
wire n_195;
wire n_261;
wire n_189;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_213;
wire n_164;
wire n_257;
wire n_100;
wire n_129;
wire n_121;
wire n_197;
wire n_137;
wire n_203;
wire n_254;
wire n_142;
wire n_143;
wire n_207;
wire n_242;
wire n_180;
wire n_62;
wire n_155;
wire n_219;
wire n_75;
wire n_109;
wire n_150;
wire n_233;
wire n_263;
wire n_122;
wire n_264;
wire n_255;
wire n_205;
wire n_140;
wire n_218;
wire n_70;
wire n_120;
wire n_234;
wire n_251;
wire n_214;
wire n_67;
wire n_82;
wire n_236;
wire n_246;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_237;
wire n_81;
wire n_59;
wire n_244;
wire n_181;
wire n_76;
wire n_182;
wire n_124;
wire n_238;
wire n_243;
wire n_55;
wire n_126;
wire n_202;
wire n_97;
wire n_108;
wire n_94;
wire n_239;
wire n_267;
wire n_58;
wire n_116;
wire n_211;
wire n_64;
wire n_220;
wire n_117;
wire n_118;
wire n_175;
wire n_224;
wire n_231;
wire n_65;
wire n_230;
wire n_93;
wire n_80;
wire n_141;
wire n_240;
wire n_135;
wire n_196;
wire n_200;
wire n_165;
wire n_139;
wire n_134;
wire n_259;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_95;
wire n_179;
wire n_248;
wire n_107;
wire n_71;
wire n_74;
wire n_229;
wire n_253;
wire n_190;
wire n_123;
wire n_262;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_249;
wire n_173;
wire n_201;
wire n_250;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_183;
wire n_232;
wire n_115;
wire n_69;
wire n_128;
wire n_241;
wire n_79;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_56;
wire n_221;

INVxp33_ASAP7_75t_SL g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_30),
.Y(n_51)
);

INVxp33_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_4),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_23),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_73),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_50),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_0),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_1),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_52),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_105),
.B(n_50),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_105),
.B(n_77),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_56),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_77),
.Y(n_115)
);

O2A1O1Ixp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_97),
.B(n_103),
.C(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_81),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_69),
.B1(n_58),
.B2(n_53),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_69),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_58),
.B1(n_53),
.B2(n_3),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_1),
.Y(n_123)
);

AOI221xp5_ASAP7_75t_L g124 ( 
.A1(n_82),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.C(n_7),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_125)
);

BUFx8_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_104),
.B(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2x1p5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_95),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_93),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

AND2x4_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_119),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_87),
.B(n_97),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_140),
.A2(n_111),
.B1(n_115),
.B2(n_109),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_109),
.Y(n_147)
);

AOI21x1_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_87),
.B(n_110),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_141),
.B(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_115),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_110),
.B(n_122),
.C(n_96),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_98),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

CKINVDCx8_ASAP7_75t_R g156 ( 
.A(n_140),
.Y(n_156)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

AND2x4_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_83),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_124),
.B1(n_125),
.B2(n_101),
.Y(n_159)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_83),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_91),
.B1(n_98),
.B2(n_126),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_152),
.A2(n_132),
.B(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

AOI21x1_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_128),
.B(n_136),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

OR2x6_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_132),
.Y(n_170)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_136),
.B(n_127),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_98),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_91),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_145),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_152),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_153),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_156),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_160),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_162),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

NOR4xp25_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_161),
.C(n_173),
.D(n_146),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_172),
.B(n_154),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_182),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_188),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_170),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_170),
.B1(n_167),
.B2(n_171),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_171),
.B1(n_126),
.B2(n_169),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_169),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_175),
.C(n_168),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_195),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

NAND2x1p5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_197),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_197),
.B1(n_189),
.B2(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_181),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_207),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_215),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_207),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_206),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_226),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_221),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_201),
.B1(n_187),
.B2(n_190),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_199),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_209),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_229),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_SL g245 ( 
.A1(n_240),
.A2(n_8),
.B(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_235),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_240),
.Y(n_251)
);

NAND4xp25_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_241),
.C(n_238),
.D(n_234),
.Y(n_252)
);

NAND4xp25_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_246),
.C(n_249),
.D(n_248),
.Y(n_253)
);

AOI211xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_239),
.B(n_233),
.C(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_235),
.Y(n_255)
);

AOI221xp5_ASAP7_75t_L g256 ( 
.A1(n_252),
.A2(n_253),
.B1(n_251),
.B2(n_254),
.C(n_255),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_259),
.A2(n_250),
.B1(n_236),
.B2(n_237),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

AOI211xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_212),
.B(n_12),
.C(n_13),
.Y(n_263)
);

OR4x1_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_10),
.C(n_15),
.D(n_16),
.Y(n_264)
);

OAI22x1_ASAP7_75t_L g265 ( 
.A1(n_263),
.A2(n_200),
.B1(n_198),
.B2(n_211),
.Y(n_265)
);

OAI322xp33_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_17),
.A3(n_19),
.B1(n_21),
.B2(n_22),
.C1(n_27),
.C2(n_29),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_32),
.B(n_33),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_35),
.B(n_37),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_171),
.B1(n_175),
.B2(n_41),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_270),
.A2(n_269),
.B1(n_268),
.B2(n_45),
.Y(n_271)
);


endmodule