module real_jpeg_18701_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_556),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_0),
.B(n_557),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_1),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_1),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_1),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_1),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_1),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_1),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_1),
.B(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_1),
.A2(n_6),
.B1(n_268),
.B2(n_272),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_1),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_2),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_2),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_2),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_2),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_2),
.B(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_2),
.B(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_2),
.B(n_494),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_3),
.Y(n_96)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_3),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_3),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_4),
.Y(n_98)
);

NAND2x1_ASAP7_75t_L g103 ( 
.A(n_4),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_4),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_4),
.B(n_156),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_4),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_4),
.B(n_42),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_4),
.B(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_4),
.B(n_229),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g375 ( 
.A(n_5),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_6),
.B(n_74),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_6),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_6),
.B(n_339),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_6),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_6),
.B(n_219),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_6),
.B(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_6),
.B(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_6),
.B(n_94),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_7),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_7),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_7),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_7),
.B(n_219),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_7),
.B(n_290),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_7),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_7),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_8),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_8),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_8),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_8),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_8),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_8),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_8),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_8),
.B(n_550),
.Y(n_549)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_9),
.Y(n_235)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_9),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_9),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_10),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_11),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_11),
.B(n_57),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_11),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_11),
.B(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_11),
.B(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_11),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g333 ( 
.A(n_11),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_12),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_12),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_12),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_12),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_12),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_12),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_12),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_12),
.B(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_13),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_14),
.Y(n_40)
);

AND2x4_ASAP7_75t_SL g93 ( 
.A(n_14),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_14),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_14),
.B(n_58),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_14),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_15),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_16),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_16),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_16),
.Y(n_220)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_16),
.Y(n_286)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_16),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_18),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_539),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_257),
.B(n_534),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_171),
.C(n_251),
.Y(n_23)
);

OAI21x1_ASAP7_75t_SL g534 ( 
.A1(n_24),
.A2(n_535),
.B(n_538),
.Y(n_534)
);

NOR2x1_ASAP7_75t_R g24 ( 
.A(n_25),
.B(n_147),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_25),
.B(n_147),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_110),
.C(n_125),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_26),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_72),
.C(n_90),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_28),
.B(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_48),
.C(n_61),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_29),
.B(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_37),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_30),
.B(n_39),
.C(n_43),
.Y(n_123)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_36),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_36),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_36),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_38),
.A2(n_39),
.B1(n_113),
.B2(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_SL g128 ( 
.A(n_39),
.B(n_113),
.C(n_118),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_40),
.B(n_547),
.Y(n_546)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_43),
.A2(n_44),
.B1(n_93),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_44),
.B(n_93),
.C(n_97),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_46),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_47),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_48),
.B(n_61),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.C(n_56),
.Y(n_48)
);

XNOR2x1_ASAP7_75t_L g196 ( 
.A(n_49),
.B(n_56),
.Y(n_196)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2x1_ASAP7_75t_L g195 ( 
.A(n_53),
.B(n_196),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g464 ( 
.A(n_55),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_59),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_67),
.C(n_71),
.Y(n_124)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_65),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_70),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_72),
.B(n_90),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_73),
.B(n_84),
.C(n_89),
.Y(n_146)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_85),
.B2(n_89),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_83),
.Y(n_274)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_101),
.C(n_107),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_91),
.A2(n_92),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_93),
.B(n_198),
.C(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_93),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_93),
.A2(n_199),
.B1(n_206),
.B2(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_96),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_97),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_97),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_97),
.A2(n_203),
.B1(n_278),
.B2(n_326),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_101),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_103),
.B(n_107),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_103),
.B(n_228),
.C(n_231),
.Y(n_227)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_105),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_107),
.A2(n_190),
.B1(n_193),
.B2(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_110),
.A2(n_125),
.B1(n_126),
.B2(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_110),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_123),
.C(n_124),
.Y(n_110)
);

XNOR2x2_ASAP7_75t_L g245 ( 
.A(n_111),
.B(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_118),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_117),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_130),
.C(n_134),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_122),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_123),
.B(n_124),
.Y(n_246)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_136),
.C(n_170),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_134),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_135),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_134),
.B(n_155),
.C(n_157),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_146),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_141),
.C(n_146),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_169),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_149),
.B(n_150),
.C(n_169),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_164),
.B2(n_165),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_151),
.B(n_166),
.C(n_168),
.Y(n_553)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_154),
.A2(n_155),
.B1(n_546),
.B2(n_548),
.Y(n_545)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_241),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g536 ( 
.A(n_172),
.B(n_241),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_207),
.C(n_209),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_173),
.B(n_207),
.Y(n_355)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_194),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_175),
.B(n_178),
.C(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_190),
.C(n_193),
.Y(n_178)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_179),
.B(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.C(n_188),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_188),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_182),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_192),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_194),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.C(n_202),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_195),
.B(n_197),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_200),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_201),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_202),
.B(n_306),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_203),
.B(n_276),
.C(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_209),
.B(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_226),
.C(n_238),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_210),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.C(n_224),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_211),
.B(n_214),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.C(n_221),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_215),
.A2(n_221),
.B1(n_222),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_215),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_218),
.B(n_351),
.Y(n_350)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_221),
.B(n_399),
.C(n_402),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_221),
.A2(n_222),
.B1(n_399),
.B2(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_224),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_226),
.B(n_238),
.Y(n_308)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_234),
.C(n_236),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_SL g301 ( 
.A(n_227),
.B(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_233),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_234),
.Y(n_303)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_235),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_236),
.A2(n_237),
.B1(n_371),
.B2(n_372),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_237),
.B(n_364),
.C(n_371),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_245),
.C(n_249),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_245),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AOI21x1_ASAP7_75t_L g535 ( 
.A1(n_252),
.A2(n_536),
.B(n_537),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_253),
.B(n_256),
.Y(n_537)
);

AO21x2_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_358),
.B(n_531),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_353),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_311),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_260),
.B(n_311),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_304),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_261),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_281),
.C(n_300),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_263),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.C(n_275),
.Y(n_263)
);

XNOR2x2_ASAP7_75t_L g410 ( 
.A(n_264),
.B(n_411),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_266),
.A2(n_267),
.B1(n_275),
.B2(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_267),
.A2(n_378),
.B(n_384),
.Y(n_377)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_271),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_275),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_281),
.A2(n_300),
.B1(n_301),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_293),
.C(n_297),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.C(n_289),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_283),
.B(n_287),
.C(n_289),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_283),
.B(n_289),
.Y(n_390)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_283),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_286),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_287),
.B(n_390),
.Y(n_389)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_292),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_293),
.A2(n_294),
.B1(n_297),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_297),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_299),
.Y(n_401)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_304)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_305),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_310),
.C(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.C(n_320),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_313),
.A2(n_314),
.B1(n_317),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_317),
.Y(n_419)
);

XOR2x2_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_321),
.B(n_418),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_346),
.C(n_350),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_322),
.B(n_414),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_327),
.C(n_337),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_L g405 ( 
.A(n_324),
.B(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_327),
.B(n_337),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_333),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_328),
.B(n_333),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_335),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.C(n_342),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_338),
.A2(n_341),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_338),
.Y(n_395)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_341),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_341),
.A2(n_396),
.B1(n_471),
.B2(n_472),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_341),
.B(n_471),
.C(n_477),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_342),
.B(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_346),
.B(n_350),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_353),
.A2(n_532),
.B(n_533),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_354),
.B(n_356),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_527),
.Y(n_358)
);

NAND3xp33_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_415),
.C(n_420),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_407),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_SL g530 ( 
.A(n_361),
.B(n_407),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_391),
.C(n_405),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_362),
.B(n_525),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_376),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_377),
.C(n_389),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_364),
.B(n_516),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_365),
.B(n_368),
.Y(n_461)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_365),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_365),
.A2(n_480),
.B1(n_481),
.B2(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_370),
.Y(n_388)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_389),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_392),
.B(n_405),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_397),
.C(n_403),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_393),
.B(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_398),
.B(n_404),
.Y(n_511)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_399),
.Y(n_457)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_413),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_410),
.C(n_413),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_416),
.Y(n_529)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_417),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_421),
.A2(n_522),
.B(n_526),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_507),
.B(n_521),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_423),
.A2(n_465),
.B(n_506),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_452),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_424),
.B(n_452),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_439),
.C(n_446),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_426),
.B(n_502),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_428),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_430),
.C(n_434),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_434),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_439),
.A2(n_440),
.B1(n_446),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_441),
.B(n_443),
.Y(n_478)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_446),
.Y(n_503)
);

AO22x1_ASAP7_75t_SL g446 ( 
.A1(n_447),
.A2(n_449),
.B1(n_450),
.B2(n_451),
.Y(n_446)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_447),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_449),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_450),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_451),
.B(n_493),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_458),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_454),
.B(n_458),
.C(n_520),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_455),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

MAJx2_ASAP7_75t_L g518 ( 
.A(n_459),
.B(n_461),
.C(n_462),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_466),
.A2(n_500),
.B(n_505),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_467),
.A2(n_482),
.B(n_499),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_479),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_468),
.B(n_479),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_469),
.A2(n_470),
.B1(n_477),
.B2(n_478),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_481),
.Y(n_491)
);

AOI21x1_ASAP7_75t_SL g482 ( 
.A1(n_483),
.A2(n_492),
.B(n_498),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_490),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_490),
.Y(n_498)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_504),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_501),
.B(n_504),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_508),
.B(n_519),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_519),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_509),
.A2(n_510),
.B1(n_512),
.B2(n_513),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_509),
.B(n_514),
.C(n_518),
.Y(n_523)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_514),
.A2(n_515),
.B1(n_517),
.B2(n_518),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_524),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_524),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.C(n_530),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_555),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_554),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_541),
.B(n_554),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_553),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_544),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_549),
.Y(n_544)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_546),
.Y(n_548)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx6_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);


endmodule