module fake_ariane_1753_n_666 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_666);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_666;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_244;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_663;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_665;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_661;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_306;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_10),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_37),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_51),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_47),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_8),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_57),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_106),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_110),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_7),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_71),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_114),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_61),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_91),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_64),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_24),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_86),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_55),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_12),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_13),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_90),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_66),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_39),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_45),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_78),
.Y(n_180)
);

BUFx8_ASAP7_75t_SL g181 ( 
.A(n_46),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_65),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_30),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_28),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_25),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_136),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_63),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_119),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_124),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_72),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_100),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_40),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_6),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_49),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_50),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_12),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_52),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_17),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_69),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_0),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_94),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_29),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_54),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_9),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_97),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_139),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_59),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_156),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_181),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_146),
.B(n_166),
.Y(n_216)
);

INVxp33_ASAP7_75t_SL g217 ( 
.A(n_151),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_R g218 ( 
.A(n_155),
.B(n_18),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_144),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_181),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_159),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_158),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_156),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_173),
.Y(n_226)
);

BUFx6f_ASAP7_75t_SL g227 ( 
.A(n_163),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_0),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_173),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_175),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_197),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_202),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_204),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_177),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_145),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_195),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_148),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_153),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_154),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_160),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_147),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_161),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_149),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_150),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_152),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_157),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_165),
.B(n_1),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_167),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_162),
.B(n_1),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_172),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_179),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_171),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_219),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_205),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_214),
.A2(n_162),
.B1(n_169),
.B2(n_176),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

OA21x2_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_182),
.B(n_190),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_229),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_238),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_255),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_214),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_220),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_259),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_231),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_228),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_217),
.A2(n_216),
.B1(n_241),
.B2(n_259),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g294 ( 
.A(n_222),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_243),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_244),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_225),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_247),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_249),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_227),
.B(n_169),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_178),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_226),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_235),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_236),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_218),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_239),
.B(n_183),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_225),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_232),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_237),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_237),
.B1(n_192),
.B2(n_189),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_180),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_270),
.B(n_185),
.Y(n_315)
);

BUFx8_ASAP7_75t_SL g316 ( 
.A(n_294),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_279),
.B(n_196),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_261),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_203),
.C(n_207),
.Y(n_321)
);

AND2x6_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_170),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_262),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_281),
.B(n_210),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_271),
.A2(n_170),
.B1(n_176),
.B2(n_186),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_291),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_265),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_272),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_283),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_186),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_283),
.B(n_187),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_278),
.B(n_188),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_273),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_261),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_268),
.Y(n_339)
);

AND2x6_ASAP7_75t_L g340 ( 
.A(n_290),
.B(n_186),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_268),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_191),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_263),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_278),
.B(n_193),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_304),
.B(n_260),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_304),
.B(n_194),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_269),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_269),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_305),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_307),
.B(n_186),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_307),
.B(n_198),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_277),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_287),
.Y(n_356)
);

BUFx10_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_264),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_295),
.B(n_199),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_295),
.B(n_296),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_305),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_274),
.B(n_201),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_277),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_305),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_286),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_277),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_276),
.B(n_206),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_308),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_296),
.B(n_212),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_304),
.B(n_208),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_289),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_303),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_303),
.B(n_306),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_312),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_282),
.B(n_211),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_299),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_306),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g380 ( 
.A(n_299),
.B(n_19),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_282),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_338),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_320),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_360),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_282),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_300),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_300),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_352),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_339),
.A2(n_300),
.B(n_263),
.Y(n_390)
);

O2A1O1Ixp5_ASAP7_75t_L g391 ( 
.A1(n_344),
.A2(n_300),
.B(n_311),
.C(n_310),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_356),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_325),
.A2(n_300),
.B1(n_310),
.B2(n_267),
.Y(n_393)
);

NAND3xp33_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_288),
.C(n_280),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_267),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_2),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_347),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_314),
.A2(n_288),
.B1(n_284),
.B2(n_280),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_2),
.Y(n_400)
);

A2O1A1Ixp33_ASAP7_75t_L g401 ( 
.A1(n_317),
.A2(n_284),
.B(n_302),
.C(n_309),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_323),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_366),
.A2(n_294),
.B1(n_309),
.B2(n_5),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_371),
.B(n_3),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_357),
.B(n_285),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_371),
.B(n_3),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_375),
.B(n_285),
.Y(n_407)
);

AND3x1_ASAP7_75t_L g408 ( 
.A(n_346),
.B(n_297),
.C(n_5),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_4),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_366),
.B(n_297),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_338),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_348),
.B(n_4),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_6),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_375),
.B(n_7),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_368),
.Y(n_415)
);

NOR3xp33_ASAP7_75t_L g416 ( 
.A(n_313),
.B(n_8),
.C(n_9),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_319),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_363),
.B(n_10),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_325),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_315),
.B(n_11),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_338),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_313),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_333),
.B(n_15),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_333),
.B(n_345),
.Y(n_426)
);

OAI221xp5_ASAP7_75t_L g427 ( 
.A1(n_373),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.C(n_21),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_326),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_367),
.Y(n_429)
);

INVxp33_ASAP7_75t_L g430 ( 
.A(n_343),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_330),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_351),
.B(n_22),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_351),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_337),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_362),
.B(n_23),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_376),
.B(n_26),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_328),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_345),
.B(n_143),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_362),
.B(n_27),
.Y(n_439)
);

NAND3xp33_ASAP7_75t_SL g440 ( 
.A(n_332),
.B(n_31),
.C(n_32),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_317),
.B(n_324),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_376),
.B(n_142),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_347),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_347),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_361),
.B(n_33),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_349),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_445),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_384),
.B(n_369),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

AO21x1_ASAP7_75t_L g451 ( 
.A1(n_426),
.A2(n_353),
.B(n_331),
.Y(n_451)
);

AO22x1_ASAP7_75t_L g452 ( 
.A1(n_416),
.A2(n_380),
.B1(n_322),
.B2(n_316),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_384),
.B(n_364),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_402),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_437),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_423),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_434),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_329),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_417),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_324),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_422),
.B(n_429),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_334),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_415),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_397),
.B(n_347),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_383),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_395),
.B(n_350),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_SL g469 ( 
.A(n_397),
.B(n_377),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_400),
.B(n_335),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_336),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_392),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_441),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_399),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_400),
.B(n_321),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_445),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_409),
.B(n_322),
.Y(n_477)
);

OAI221xp5_ASAP7_75t_L g478 ( 
.A1(n_424),
.A2(n_354),
.B1(n_342),
.B2(n_353),
.C(n_331),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_447),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_446),
.B(n_365),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_430),
.Y(n_482)
);

AND2x6_ASAP7_75t_SL g483 ( 
.A(n_409),
.B(n_380),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_382),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_446),
.B(n_365),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_407),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_R g488 ( 
.A(n_440),
.B(n_322),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_396),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

AOI21xp33_ASAP7_75t_L g492 ( 
.A1(n_449),
.A2(n_393),
.B(n_404),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_456),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_451),
.A2(n_438),
.B(n_425),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_450),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_454),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_460),
.B(n_424),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_449),
.B(n_432),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g500 ( 
.A1(n_487),
.A2(n_490),
.B(n_406),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_477),
.A2(n_391),
.B(n_355),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_489),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_453),
.A2(n_381),
.B(n_388),
.Y(n_503)
);

OAI21x1_ASAP7_75t_SL g504 ( 
.A1(n_470),
.A2(n_412),
.B(n_413),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_SL g505 ( 
.A(n_474),
.B(n_416),
.C(n_401),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_453),
.B(n_465),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_472),
.Y(n_507)
);

AOI221x1_ASAP7_75t_L g508 ( 
.A1(n_475),
.A2(n_419),
.B1(n_432),
.B2(n_420),
.C(n_403),
.Y(n_508)
);

NOR3xp33_ASAP7_75t_L g509 ( 
.A(n_481),
.B(n_394),
.C(n_427),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_465),
.B(n_393),
.Y(n_510)
);

AOI221x1_ASAP7_75t_L g511 ( 
.A1(n_468),
.A2(n_469),
.B1(n_390),
.B2(n_387),
.C(n_479),
.Y(n_511)
);

AO31x2_ASAP7_75t_L g512 ( 
.A1(n_468),
.A2(n_385),
.A3(n_411),
.B(n_421),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_480),
.A2(n_410),
.B1(n_405),
.B2(n_414),
.Y(n_513)
);

BUFx6f_ASAP7_75t_SL g514 ( 
.A(n_480),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_461),
.B(n_386),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_480),
.B(n_414),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_485),
.A2(n_444),
.B(n_439),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_407),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_485),
.A2(n_415),
.B(n_435),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_491),
.B(n_443),
.Y(n_520)
);

AOI21xp33_ASAP7_75t_L g521 ( 
.A1(n_486),
.A2(n_418),
.B(n_355),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_463),
.B(n_436),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_506),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_495),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_498),
.A2(n_486),
.B1(n_457),
.B2(n_480),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_512),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_512),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_502),
.B(n_491),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_512),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_505),
.B(n_482),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_511),
.A2(n_478),
.B(n_484),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_495),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_501),
.A2(n_466),
.B(n_448),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_501),
.A2(n_473),
.B(n_462),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_498),
.B(n_459),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_499),
.A2(n_492),
.B1(n_510),
.B2(n_522),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_514),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_519),
.A2(n_448),
.B(n_458),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_514),
.Y(n_539)
);

NAND2x1_ASAP7_75t_L g540 ( 
.A(n_504),
.B(n_476),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_512),
.Y(n_541)
);

O2A1O1Ixp33_ASAP7_75t_SL g542 ( 
.A1(n_499),
.A2(n_464),
.B(n_459),
.C(n_483),
.Y(n_542)
);

OA21x2_ASAP7_75t_L g543 ( 
.A1(n_503),
.A2(n_471),
.B(n_380),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_512),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_506),
.A2(n_452),
.B(n_491),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_504),
.A2(n_380),
.B(n_464),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_515),
.A2(n_471),
.B(n_491),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_494),
.A2(n_380),
.B(n_488),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_510),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_530),
.A2(n_514),
.B1(n_522),
.B2(n_518),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_532),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_535),
.A2(n_509),
.B1(n_493),
.B2(n_513),
.Y(n_552)
);

AO21x2_ASAP7_75t_L g553 ( 
.A1(n_526),
.A2(n_517),
.B(n_516),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_523),
.A2(n_496),
.B1(n_497),
.B2(n_507),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_525),
.A2(n_467),
.B1(n_322),
.B2(n_500),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_SL g556 ( 
.A1(n_547),
.A2(n_508),
.B1(n_537),
.B2(n_523),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_524),
.B(n_502),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_536),
.A2(n_322),
.B1(n_500),
.B2(n_476),
.Y(n_558)
);

AOI221xp5_ASAP7_75t_L g559 ( 
.A1(n_542),
.A2(n_521),
.B1(n_488),
.B2(n_493),
.C(n_489),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_R g560 ( 
.A(n_539),
.B(n_500),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_SL g561 ( 
.A(n_540),
.B(n_489),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_534),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_540),
.A2(n_494),
.B(n_520),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_549),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_545),
.A2(n_494),
.B(n_520),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_537),
.B(n_502),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_549),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_537),
.B(n_489),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_537),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_548),
.A2(n_327),
.B(n_340),
.C(n_36),
.Y(n_570)
);

CKINVDCx6p67_ASAP7_75t_R g571 ( 
.A(n_526),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_538),
.B(n_34),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_534),
.B(n_340),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_534),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_528),
.B(n_534),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_541),
.A2(n_340),
.B1(n_327),
.B2(n_41),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_528),
.B(n_35),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_528),
.B(n_340),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_541),
.A2(n_340),
.B1(n_327),
.B2(n_43),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_531),
.Y(n_580)
);

AOI221xp5_ASAP7_75t_L g581 ( 
.A1(n_554),
.A2(n_544),
.B1(n_529),
.B2(n_527),
.C(n_531),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_574),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_564),
.A2(n_544),
.B1(n_529),
.B2(n_527),
.Y(n_583)
);

AOI222xp33_ASAP7_75t_L g584 ( 
.A1(n_552),
.A2(n_527),
.B1(n_529),
.B2(n_548),
.C1(n_546),
.C2(n_538),
.Y(n_584)
);

AOI221xp5_ASAP7_75t_L g585 ( 
.A1(n_554),
.A2(n_531),
.B1(n_543),
.B2(n_546),
.C(n_533),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_550),
.A2(n_543),
.B1(n_531),
.B2(n_533),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_567),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_551),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_556),
.A2(n_543),
.B1(n_327),
.B2(n_44),
.Y(n_589)
);

AOI221xp5_ASAP7_75t_L g590 ( 
.A1(n_580),
.A2(n_543),
.B1(n_42),
.B2(n_48),
.C(n_53),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_557),
.B(n_38),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_555),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_558),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_593)
);

AOI211xp5_ASAP7_75t_L g594 ( 
.A1(n_577),
.A2(n_75),
.B(n_77),
.C(n_79),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_580),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_595)
);

OAI21xp33_ASAP7_75t_L g596 ( 
.A1(n_572),
.A2(n_83),
.B(n_84),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_563),
.A2(n_85),
.B(n_87),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_571),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_SL g599 ( 
.A1(n_572),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_579),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_569),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_566),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_553),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_582),
.B(n_575),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_588),
.B(n_566),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_553),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_598),
.B(n_568),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_582),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_601),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_603),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_602),
.B(n_601),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_597),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_602),
.Y(n_613)
);

OAI221xp5_ASAP7_75t_L g614 ( 
.A1(n_596),
.A2(n_560),
.B1(n_565),
.B2(n_559),
.C(n_570),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_583),
.B(n_565),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_583),
.B(n_562),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_581),
.B(n_573),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_586),
.B(n_573),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_604),
.B(n_605),
.Y(n_619)
);

AOI221xp5_ASAP7_75t_L g620 ( 
.A1(n_615),
.A2(n_614),
.B1(n_617),
.B2(n_589),
.C(n_607),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_609),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_L g622 ( 
.A(n_607),
.B(n_594),
.C(n_590),
.Y(n_622)
);

INVxp67_ASAP7_75t_R g623 ( 
.A(n_604),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_R g624 ( 
.A(n_613),
.B(n_561),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_606),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_615),
.A2(n_592),
.B1(n_593),
.B2(n_595),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_625),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_619),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_621),
.B(n_608),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_624),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_623),
.B(n_611),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_620),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_620),
.B(n_611),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_627),
.B(n_626),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_628),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_629),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_628),
.B(n_613),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_611),
.Y(n_638)
);

NOR4xp25_ASAP7_75t_SL g639 ( 
.A(n_636),
.B(n_630),
.C(n_632),
.D(n_634),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_635),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_634),
.A2(n_622),
.B1(n_633),
.B2(n_629),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_637),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_638),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_640),
.Y(n_644)
);

OAI21xp33_ASAP7_75t_L g645 ( 
.A1(n_641),
.A2(n_615),
.B(n_595),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_639),
.A2(n_599),
.B(n_592),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_644),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_645),
.B(n_643),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_647),
.Y(n_649)
);

NOR3x1_ASAP7_75t_L g650 ( 
.A(n_649),
.B(n_646),
.C(n_642),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_650),
.A2(n_648),
.B(n_640),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_651),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_652),
.Y(n_653)
);

OAI211xp5_ASAP7_75t_SL g654 ( 
.A1(n_653),
.A2(n_593),
.B(n_591),
.C(n_600),
.Y(n_654)
);

O2A1O1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_654),
.A2(n_612),
.B(n_576),
.C(n_578),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_655),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_656),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_657),
.Y(n_658)
);

OAI222xp33_ASAP7_75t_L g659 ( 
.A1(n_658),
.A2(n_612),
.B1(n_616),
.B2(n_618),
.C1(n_610),
.C2(n_585),
.Y(n_659)
);

AOI21xp33_ASAP7_75t_L g660 ( 
.A1(n_658),
.A2(n_101),
.B(n_102),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_660),
.B(n_103),
.Y(n_661)
);

OAI321xp33_ASAP7_75t_L g662 ( 
.A1(n_659),
.A2(n_104),
.A3(n_105),
.B1(n_107),
.B2(n_109),
.C(n_111),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_661),
.A2(n_584),
.B1(n_115),
.B2(n_116),
.Y(n_663)
);

AOI322xp5_ASAP7_75t_L g664 ( 
.A1(n_662),
.A2(n_112),
.A3(n_118),
.B1(n_121),
.B2(n_123),
.C1(n_129),
.C2(n_131),
.Y(n_664)
);

OAI221xp5_ASAP7_75t_L g665 ( 
.A1(n_663),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.C(n_137),
.Y(n_665)
);

AOI211xp5_ASAP7_75t_L g666 ( 
.A1(n_665),
.A2(n_664),
.B(n_140),
.C(n_141),
.Y(n_666)
);


endmodule