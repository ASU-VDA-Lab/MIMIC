module fake_jpeg_18475_n_162 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_162);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR3xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_10),
.C(n_1),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_12),
.B1(n_21),
.B2(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_29),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_28),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_41),
.Y(n_52)
);

AND2x6_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_32),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_16),
.B1(n_19),
.B2(n_18),
.Y(n_49)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_57),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_20),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx24_ASAP7_75t_SL g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx24_ASAP7_75t_SL g70 ( 
.A(n_62),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_67),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_47),
.B1(n_48),
.B2(n_42),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_33),
.B1(n_44),
.B2(n_36),
.Y(n_86)
);

AOI31xp33_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_19),
.A3(n_16),
.B(n_18),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_74),
.B1(n_54),
.B2(n_22),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_26),
.B1(n_36),
.B2(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_61),
.B(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_80),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_59),
.B(n_57),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_82),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_14),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_52),
.C(n_63),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_63),
.C(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_72),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_94),
.C(n_31),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_46),
.C(n_43),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_21),
.Y(n_107)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_100),
.B1(n_33),
.B2(n_37),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_20),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_14),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_112),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_26),
.B1(n_37),
.B2(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_17),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_101),
.B(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_111),
.B(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_33),
.B1(n_29),
.B2(n_25),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_37),
.B1(n_25),
.B2(n_29),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_94),
.B1(n_89),
.B2(n_93),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_124),
.B1(n_114),
.B2(n_110),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_R g123 ( 
.A1(n_112),
.A2(n_17),
.B(n_15),
.Y(n_123)
);

NOR2x1_ASAP7_75t_R g131 ( 
.A(n_123),
.B(n_108),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_17),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_126),
.B(n_0),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_113),
.B1(n_109),
.B2(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_123),
.B1(n_122),
.B2(n_116),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_132),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_29),
.B1(n_24),
.B2(n_31),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_134),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_31),
.B(n_17),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_139),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_121),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_141),
.C(n_135),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_116),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_144),
.C(n_15),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_130),
.C(n_15),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_2),
.B(n_3),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_2),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_4),
.B(n_5),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_3),
.B(n_4),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_4),
.B(n_6),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_147),
.A2(n_142),
.B1(n_24),
.B2(n_6),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_6),
.B(n_7),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_7),
.B(n_8),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_10),
.B(n_8),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_156),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_SL g159 ( 
.A(n_157),
.B(n_152),
.C(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_155),
.B1(n_158),
.B2(n_9),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_9),
.Y(n_162)
);


endmodule