module fake_jpeg_23781_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx2_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_12),
.Y(n_34)
);

CKINVDCx12_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_10),
.B1(n_23),
.B2(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_31),
.B1(n_10),
.B2(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_39),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_27),
.A2(n_22),
.B(n_13),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_13),
.B(n_11),
.Y(n_51)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_14),
.Y(n_48)
);

AND2x4_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_22),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_45),
.B(n_29),
.C(n_24),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_15),
.B(n_18),
.C(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_0),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_11),
.C(n_37),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_5),
.Y(n_74)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_66),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_50),
.B(n_28),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_54),
.B1(n_51),
.B2(n_52),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_20),
.B1(n_39),
.B2(n_10),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_49),
.C(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_72),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_61),
.B1(n_59),
.B2(n_65),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_74),
.B(n_76),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_75),
.Y(n_78)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_61),
.B1(n_66),
.B2(n_64),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_83),
.B1(n_71),
.B2(n_73),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_60),
.C(n_58),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_84),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_87),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_70),
.B(n_1),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_88)
);

AO21x1_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_84),
.B(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_79),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_17),
.C(n_3),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_81),
.C(n_17),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_93),
.C(n_0),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_85),
.B(n_89),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_0),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_96),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_100),
.B(n_4),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_100),
.C(n_4),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g108 ( 
.A(n_107),
.Y(n_108)
);


endmodule