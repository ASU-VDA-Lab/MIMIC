module fake_jpeg_2551_n_229 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_229);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_83),
.Y(n_95)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_49),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_57),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_98),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_70),
.B1(n_61),
.B2(n_64),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_96),
.B1(n_84),
.B2(n_60),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_85),
.A2(n_70),
.B1(n_61),
.B2(n_74),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_68),
.B(n_74),
.C(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_53),
.B1(n_64),
.B2(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_53),
.B1(n_72),
.B2(n_55),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_101),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_97),
.Y(n_103)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_115),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_65),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_66),
.C(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_117),
.Y(n_118)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_78),
.B1(n_81),
.B2(n_98),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_78),
.Y(n_117)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_67),
.A3(n_56),
.B1(n_75),
.B2(n_73),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_123),
.Y(n_154)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_30),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_135),
.Y(n_153)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_132),
.B1(n_111),
.B2(n_58),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_62),
.B1(n_55),
.B2(n_54),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_54),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_136),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_99),
.B(n_0),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_1),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_1),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_5),
.Y(n_161)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_141),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_114),
.B1(n_58),
.B2(n_71),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_143),
.B1(n_39),
.B2(n_38),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_139),
.A2(n_114),
.B1(n_58),
.B2(n_63),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_23),
.B(n_48),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_158),
.B(n_32),
.Y(n_172)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_148),
.Y(n_171)
);

NAND2x1_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_63),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_9),
.B(n_10),
.Y(n_178)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_47),
.C(n_46),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_155),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_2),
.B(n_3),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_44),
.C(n_43),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_161),
.B(n_11),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_42),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_122),
.Y(n_164)
);

OAI22x1_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_123),
.B1(n_138),
.B2(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_170),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_167),
.A2(n_176),
.B1(n_12),
.B2(n_13),
.Y(n_197)
);

OAI22x1_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_149),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_178),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_31),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_159),
.C(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_180),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_28),
.B(n_27),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_183),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_25),
.B(n_22),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_171),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_150),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_196),
.C(n_14),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_140),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_193),
.Y(n_205)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_11),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_208)
);

AOI221xp5_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_165),
.B1(n_163),
.B2(n_176),
.C(n_167),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_199),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_172),
.B(n_168),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_166),
.B1(n_175),
.B2(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_182),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_202),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_189),
.A2(n_184),
.B1(n_185),
.B2(n_192),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_12),
.Y(n_203)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_203),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

AOI221xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_194),
.B1(n_197),
.B2(n_195),
.C(n_193),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_206),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_206),
.B1(n_201),
.B2(n_205),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_203),
.Y(n_219)
);

AOI31xp67_ASAP7_75t_SL g222 ( 
.A1(n_221),
.A2(n_214),
.A3(n_204),
.B(n_216),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_215),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_213),
.A3(n_212),
.B1(n_19),
.B2(n_20),
.C1(n_21),
.C2(n_18),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_226),
.A2(n_19),
.B(n_16),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_18),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_228),
.Y(n_229)
);


endmodule