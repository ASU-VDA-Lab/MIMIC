module real_jpeg_27504_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_281, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_281;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g61 ( 
.A(n_0),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_3),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_3),
.A2(n_41),
.B1(n_43),
.B2(n_183),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_183),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_183),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_5),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_5),
.A2(n_41),
.B1(n_43),
.B2(n_96),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_96),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_96),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_80),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_8),
.A2(n_11),
.B(n_60),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_9),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_9),
.A2(n_27),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_9),
.A2(n_27),
.B1(n_41),
.B2(n_43),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_SL g56 ( 
.A1(n_11),
.A2(n_31),
.B(n_33),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_11),
.A2(n_36),
.B1(n_59),
.B2(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_11),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_11),
.B(n_32),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_11),
.A2(n_41),
.B(n_45),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_11),
.B(n_40),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_272),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_263),
.B(n_271),
.Y(n_13)
);

OAI321xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_232),
.A3(n_256),
.B1(n_261),
.B2(n_262),
.C(n_281),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_213),
.B(n_231),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_194),
.B(n_212),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_113),
.B(n_175),
.C(n_193),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_101),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_19),
.B(n_101),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_67),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_20),
.B(n_68),
.C(n_86),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_53),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_37),
.B1(n_51),
.B2(n_52),
.Y(n_21)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_22),
.B(n_52),
.C(n_53),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_22),
.A2(n_51),
.B1(n_70),
.B2(n_104),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_22),
.B(n_104),
.C(n_200),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_22),
.A2(n_51),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_22),
.B(n_242),
.C(n_253),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_24),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_26),
.A2(n_30),
.B(n_36),
.C(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_28),
.B(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_28),
.B(n_32),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_28),
.A2(n_32),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_34),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_33),
.A2(n_36),
.B(n_46),
.C(n_120),
.Y(n_119)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_35),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_36),
.A2(n_41),
.B(n_80),
.C(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_36),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_36),
.B(n_81),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_37),
.B(n_110),
.C(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_37),
.A2(n_52),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_37),
.A2(n_219),
.B(n_221),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_37),
.B(n_219),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_39),
.B(n_40),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_39),
.A2(n_40),
.B1(n_239),
.B2(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_40),
.A2(n_239),
.B(n_240),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_43),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_50),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_48),
.B(n_190),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_57),
.A2(n_108),
.B1(n_144),
.B2(n_147),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_57),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_57),
.B(n_159),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_57),
.B(n_134),
.C(n_146),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_58),
.A2(n_66),
.B(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_59),
.B(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_62),
.B(n_63),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_62),
.A2(n_66),
.B1(n_95),
.B2(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_85),
.B2(n_86),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.C(n_82),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_70),
.A2(n_87),
.B1(n_88),
.B2(n_104),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_71),
.Y(n_240)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_77),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_75),
.A2(n_77),
.B1(n_81),
.B2(n_90),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_76),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_77),
.A2(n_81),
.B1(n_205),
.B2(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_81),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_82),
.A2(n_105),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_82),
.A2(n_105),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_82),
.A2(n_105),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_82),
.B(n_238),
.C(n_241),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_82),
.B(n_248),
.C(n_255),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_83),
.A2(n_84),
.B(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_87),
.A2(n_88),
.B1(n_141),
.B2(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_87),
.B(n_94),
.Y(n_186)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_104),
.C(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_88),
.B(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B(n_92),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_92),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_97),
.B(n_98),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.C(n_109),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_102),
.B(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_105),
.B(n_186),
.C(n_188),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_109),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_110),
.B(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_174),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_169),
.B(n_173),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_137),
.B(n_168),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_125),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_125),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_124),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_134),
.C(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_128),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_129),
.B(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_136),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_134),
.A2(n_136),
.B1(n_181),
.B2(n_184),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_134),
.B(n_181),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_163),
.B(n_167),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_148),
.B(n_162),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_143),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_144),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_152),
.B(n_161),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_158),
.B(n_160),
.Y(n_152)
);

INVx5_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_177),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_191),
.B2(n_192),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_185),
.C(n_192),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_181),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_191),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_196),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_211),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_203),
.C(n_211),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_208),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_207),
.A2(n_208),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_208),
.A2(n_223),
.B(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_215),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_229),
.B2(n_230),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_222),
.C(n_230),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_234),
.C(n_244),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_234),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_229),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_246),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_242),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_245),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_265),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_265),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_268),
.CI(n_270),
.CON(n_265),
.SN(n_265)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_277),
.Y(n_279)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);


endmodule