module real_aes_16576_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g114 ( .A(n_0), .B(n_115), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_1), .A2(n_4), .B1(n_284), .B2(n_285), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_2), .A2(n_43), .B1(n_185), .B2(n_233), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_3), .A2(n_24), .B1(n_233), .B2(n_267), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_5), .A2(n_16), .B1(n_534), .B2(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_6), .A2(n_62), .B1(n_170), .B2(n_171), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_7), .A2(n_17), .B1(n_185), .B2(n_186), .Y(n_184) );
INVx1_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_9), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_10), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_11), .A2(n_18), .B1(n_535), .B2(n_579), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_12), .A2(n_66), .B1(n_143), .B2(n_144), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
BUFx2_ASAP7_75t_L g108 ( .A(n_13), .Y(n_108) );
OR2x2_ASAP7_75t_L g132 ( .A(n_13), .B(n_38), .Y(n_132) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_14), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_15), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_19), .A2(n_99), .B1(n_285), .B2(n_534), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_20), .A2(n_39), .B1(n_163), .B2(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_21), .B(n_161), .Y(n_595) );
OAI21x1_ASAP7_75t_L g175 ( .A1(n_22), .A2(n_60), .B(n_176), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_23), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_25), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_26), .B(n_158), .Y(n_225) );
INVx4_ASAP7_75t_R g209 ( .A(n_27), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_28), .A2(n_47), .B1(n_189), .B2(n_282), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_29), .A2(n_55), .B1(n_189), .B2(n_534), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_30), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_31), .B(n_559), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_32), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_33), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g289 ( .A(n_34), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_SL g264 ( .A1(n_35), .A2(n_157), .B(n_185), .C(n_265), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_36), .A2(n_56), .B1(n_185), .B2(n_189), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g812 ( .A(n_37), .Y(n_812) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_38), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_40), .A2(n_87), .B1(n_185), .B2(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_SL g830 ( .A1(n_41), .A2(n_54), .B1(n_831), .B2(n_832), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_41), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_42), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_44), .A2(n_46), .B1(n_185), .B2(n_186), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_45), .A2(n_61), .B1(n_534), .B2(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g229 ( .A(n_48), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_49), .B(n_185), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_50), .Y(n_243) );
INVx2_ASAP7_75t_L g137 ( .A(n_51), .Y(n_137) );
INVx1_ASAP7_75t_L g117 ( .A(n_52), .Y(n_117) );
BUFx3_ASAP7_75t_L g140 ( .A(n_52), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_53), .Y(n_834) );
INVx1_ASAP7_75t_L g831 ( .A(n_54), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_57), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_58), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_59), .A2(n_88), .B1(n_185), .B2(n_189), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_63), .A2(n_76), .B1(n_282), .B2(n_551), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_64), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_65), .A2(n_79), .B1(n_185), .B2(n_186), .Y(n_536) );
INVx1_ASAP7_75t_L g144 ( .A(n_66), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_67), .A2(n_98), .B1(n_534), .B2(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g176 ( .A(n_68), .Y(n_176) );
AND2x4_ASAP7_75t_L g179 ( .A(n_69), .B(n_180), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_70), .A2(n_90), .B1(n_189), .B2(n_282), .Y(n_281) );
AO22x1_ASAP7_75t_L g159 ( .A1(n_71), .A2(n_77), .B1(n_160), .B2(n_163), .Y(n_159) );
INVx1_ASAP7_75t_L g180 ( .A(n_72), .Y(n_180) );
AND2x2_ASAP7_75t_L g268 ( .A(n_73), .B(n_221), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_74), .B(n_170), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_75), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_78), .B(n_233), .Y(n_244) );
INVx2_ASAP7_75t_L g158 ( .A(n_80), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_81), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_82), .B(n_221), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_83), .A2(n_97), .B1(n_170), .B2(n_189), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_84), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_85), .B(n_174), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_86), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_89), .B(n_221), .Y(n_600) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_91), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_92), .B(n_221), .Y(n_240) );
INVx1_ASAP7_75t_L g119 ( .A(n_93), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_93), .B(n_130), .Y(n_129) );
NAND2xp33_ASAP7_75t_L g598 ( .A(n_94), .B(n_161), .Y(n_598) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_95), .A2(n_170), .B(n_191), .C(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g214 ( .A(n_96), .B(n_215), .Y(n_214) );
NAND2xp33_ASAP7_75t_L g248 ( .A(n_100), .B(n_210), .Y(n_248) );
AOI21xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_120), .B(n_833), .Y(n_101) );
INVx6_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx6_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx8_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_111), .Y(n_105) );
OR2x6_ASAP7_75t_L g836 ( .A(n_106), .B(n_111), .Y(n_836) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .C(n_118), .Y(n_112) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g130 ( .A(n_117), .Y(n_130) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g506 ( .A(n_119), .Y(n_506) );
NAND2x1p5_ASAP7_75t_L g120 ( .A(n_121), .B(n_819), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_133), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_123), .A2(n_825), .B(n_827), .Y(n_824) );
NOR2x1_ASAP7_75t_R g123 ( .A(n_124), .B(n_125), .Y(n_123) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx3_ASAP7_75t_L g826 ( .A(n_126), .Y(n_826) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
CKINVDCx8_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
AND2x6_ASAP7_75t_SL g128 ( .A(n_129), .B(n_131), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_131), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2x1_ASAP7_75t_L g818 ( .A(n_132), .B(n_140), .Y(n_818) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_141), .B(n_811), .Y(n_133) );
BUFx12f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x6_ASAP7_75t_SL g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_137), .B(n_816), .Y(n_815) );
INVx3_ASAP7_75t_L g823 ( .A(n_137), .Y(n_823) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI22xp33_ASAP7_75t_SL g141 ( .A1(n_142), .A2(n_145), .B1(n_146), .B2(n_810), .Y(n_141) );
INVx1_ASAP7_75t_L g810 ( .A(n_142), .Y(n_810) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OAI22x1_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_504), .B1(n_507), .B2(n_809), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_414), .Y(n_148) );
NOR3xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_343), .C(n_385), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_317), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_216), .B1(n_292), .B2(n_303), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OR2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_197), .Y(n_153) );
AOI21xp33_ASAP7_75t_L g336 ( .A1(n_154), .A2(n_337), .B(n_339), .Y(n_336) );
AOI21xp33_ASAP7_75t_L g409 ( .A1(n_154), .A2(n_410), .B(n_411), .Y(n_409) );
OR2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_181), .Y(n_154) );
INVx2_ASAP7_75t_L g329 ( .A(n_155), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_155), .B(n_182), .Y(n_359) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_165), .C(n_177), .Y(n_156) );
INVx6_ASAP7_75t_L g187 ( .A(n_157), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_157), .A2(n_248), .B(n_249), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_157), .B(n_159), .Y(n_301) );
O2A1O1Ixp5_ASAP7_75t_L g593 ( .A1(n_157), .A2(n_186), .B(n_594), .C(n_595), .Y(n_593) );
BUFx8_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g168 ( .A(n_158), .Y(n_168) );
INVx1_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
INVx1_ASAP7_75t_L g228 ( .A(n_158), .Y(n_228) );
INVxp67_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g534 ( .A(n_161), .Y(n_534) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g164 ( .A(n_162), .Y(n_164) );
INVx1_ASAP7_75t_L g170 ( .A(n_162), .Y(n_170) );
INVx1_ASAP7_75t_L g172 ( .A(n_162), .Y(n_172) );
INVx3_ASAP7_75t_L g185 ( .A(n_162), .Y(n_185) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_162), .Y(n_211) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_162), .Y(n_233) );
INVx1_ASAP7_75t_L g261 ( .A(n_162), .Y(n_261) );
INVx2_ASAP7_75t_L g267 ( .A(n_162), .Y(n_267) );
OAI21xp33_ASAP7_75t_SL g224 ( .A1(n_163), .A2(n_225), .B(n_226), .Y(n_224) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g300 ( .A(n_165), .Y(n_300) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_173), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_166), .A2(n_231), .B(n_232), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_166), .A2(n_187), .B1(n_272), .B2(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g517 ( .A(n_167), .Y(n_517) );
BUFx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g246 ( .A(n_168), .Y(n_246) );
INVx1_ASAP7_75t_L g579 ( .A(n_171), .Y(n_579) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_172), .B(n_206), .Y(n_205) );
OAI21xp33_ASAP7_75t_L g177 ( .A1(n_173), .A2(n_174), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g192 ( .A(n_174), .Y(n_192) );
INVx2_ASAP7_75t_L g196 ( .A(n_174), .Y(n_196) );
INVx2_ASAP7_75t_L g202 ( .A(n_174), .Y(n_202) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_175), .Y(n_222) );
INVx1_ASAP7_75t_L g302 ( .A(n_177), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_178), .A2(n_257), .B(n_264), .Y(n_256) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
BUFx10_ASAP7_75t_L g193 ( .A(n_179), .Y(n_193) );
BUFx10_ASAP7_75t_L g235 ( .A(n_179), .Y(n_235) );
INVx1_ASAP7_75t_L g287 ( .A(n_179), .Y(n_287) );
AND2x2_ASAP7_75t_L g399 ( .A(n_181), .B(n_238), .Y(n_399) );
INVx1_ASAP7_75t_L g432 ( .A(n_181), .Y(n_432) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g294 ( .A(n_182), .B(n_239), .Y(n_294) );
AND2x2_ASAP7_75t_L g325 ( .A(n_182), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g334 ( .A(n_182), .Y(n_334) );
OR2x2_ASAP7_75t_L g353 ( .A(n_182), .B(n_199), .Y(n_353) );
AND2x2_ASAP7_75t_L g368 ( .A(n_182), .B(n_199), .Y(n_368) );
AO31x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_192), .A3(n_193), .B(n_194), .Y(n_182) );
OAI22x1_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_187), .B1(n_188), .B2(n_190), .Y(n_183) );
INVx4_ASAP7_75t_L g186 ( .A(n_185), .Y(n_186) );
INVx1_ASAP7_75t_L g535 ( .A(n_185), .Y(n_535) );
INVx1_ASAP7_75t_L g551 ( .A(n_185), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_186), .A2(n_243), .B(n_244), .C(n_245), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_187), .A2(n_190), .B1(n_281), .B2(n_283), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_187), .A2(n_516), .B1(n_517), .B2(n_518), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_187), .A2(n_190), .B1(n_525), .B2(n_527), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_187), .A2(n_533), .B1(n_536), .B2(n_537), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_187), .A2(n_517), .B1(n_549), .B2(n_550), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_187), .A2(n_517), .B1(n_558), .B2(n_560), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_187), .A2(n_517), .B1(n_568), .B2(n_569), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_187), .A2(n_537), .B1(n_578), .B2(n_580), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_187), .A2(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_189), .B(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g284 ( .A(n_189), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_190), .B(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_SL g537 ( .A(n_191), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_192), .B(n_553), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_192), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g213 ( .A(n_193), .Y(n_213) );
AO31x2_ASAP7_75t_L g514 ( .A1(n_193), .A2(n_274), .A3(n_515), .B(n_519), .Y(n_514) );
AO31x2_ASAP7_75t_L g556 ( .A1(n_193), .A2(n_523), .A3(n_557), .B(n_562), .Y(n_556) );
AO31x2_ASAP7_75t_L g576 ( .A1(n_193), .A2(n_255), .A3(n_577), .B(n_581), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx2_ASAP7_75t_L g215 ( .A(n_196), .Y(n_215) );
BUFx2_ASAP7_75t_L g255 ( .A(n_196), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_196), .B(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_196), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_198), .B(n_367), .Y(n_410) );
OR2x2_ASAP7_75t_L g498 ( .A(n_198), .B(n_359), .Y(n_498) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g326 ( .A(n_199), .Y(n_326) );
AND2x2_ASAP7_75t_L g335 ( .A(n_199), .B(n_298), .Y(n_335) );
AND2x2_ASAP7_75t_L g338 ( .A(n_199), .B(n_239), .Y(n_338) );
AND2x2_ASAP7_75t_L g357 ( .A(n_199), .B(n_238), .Y(n_357) );
AND2x4_ASAP7_75t_L g376 ( .A(n_199), .B(n_299), .Y(n_376) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_203), .B(n_214), .Y(n_199) );
AO31x2_ASAP7_75t_L g547 ( .A1(n_200), .A2(n_538), .A3(n_548), .B(n_552), .Y(n_547) );
AO31x2_ASAP7_75t_L g566 ( .A1(n_200), .A2(n_286), .A3(n_567), .B(n_570), .Y(n_566) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_202), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_SL g581 ( .A(n_202), .B(n_582), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_207), .B(n_213), .Y(n_203) );
OAI22xp33_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B1(n_211), .B2(n_212), .Y(n_208) );
INVx2_ASAP7_75t_L g282 ( .A(n_210), .Y(n_282) );
INVx1_ASAP7_75t_L g559 ( .A(n_210), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_211), .Y(n_561) );
INVx1_ASAP7_75t_L g538 ( .A(n_213), .Y(n_538) );
OAI21xp33_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_236), .B(n_277), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_217), .B(n_371), .Y(n_474) );
CKINVDCx14_ASAP7_75t_R g217 ( .A(n_218), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_219), .B(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g307 ( .A(n_219), .Y(n_307) );
OR2x2_ASAP7_75t_L g315 ( .A(n_219), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_219), .B(n_308), .Y(n_340) );
AND2x2_ASAP7_75t_L g365 ( .A(n_219), .B(n_279), .Y(n_365) );
AND2x2_ASAP7_75t_L g383 ( .A(n_219), .B(n_313), .Y(n_383) );
INVx1_ASAP7_75t_L g422 ( .A(n_219), .Y(n_422) );
AND2x2_ASAP7_75t_L g424 ( .A(n_219), .B(n_425), .Y(n_424) );
NAND2x1p5_ASAP7_75t_SL g443 ( .A(n_219), .B(n_364), .Y(n_443) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_223), .Y(n_219) );
NOR2x1_ASAP7_75t_L g250 ( .A(n_221), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g274 ( .A(n_221), .Y(n_274) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g234 ( .A(n_222), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_222), .B(n_520), .Y(n_519) );
BUFx3_ASAP7_75t_L g523 ( .A(n_222), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_222), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_222), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_SL g591 ( .A(n_222), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_230), .B(n_234), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
BUFx4f_ASAP7_75t_L g263 ( .A(n_228), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_233), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g251 ( .A(n_235), .Y(n_251) );
AO31x2_ASAP7_75t_L g270 ( .A1(n_235), .A2(n_271), .A3(n_274), .B(n_275), .Y(n_270) );
OAI32xp33_ASAP7_75t_L g327 ( .A1(n_236), .A2(n_319), .A3(n_328), .B1(n_330), .B2(n_332), .Y(n_327) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_252), .Y(n_236) );
INVx1_ASAP7_75t_L g367 ( .A(n_237), .Y(n_367) );
AND2x2_ASAP7_75t_L g375 ( .A(n_237), .B(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g374 ( .A(n_238), .B(n_298), .Y(n_374) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
BUFx3_ASAP7_75t_L g324 ( .A(n_239), .Y(n_324) );
AND2x2_ASAP7_75t_L g333 ( .A(n_239), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g439 ( .A(n_239), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_247), .B(n_250), .Y(n_241) );
INVx2_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g309 ( .A(n_252), .Y(n_309) );
OR2x2_ASAP7_75t_L g319 ( .A(n_252), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g441 ( .A(n_252), .Y(n_441) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_269), .Y(n_252) );
AND2x2_ASAP7_75t_L g342 ( .A(n_253), .B(n_270), .Y(n_342) );
INVx2_ASAP7_75t_L g364 ( .A(n_253), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_253), .B(n_279), .Y(n_384) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g291 ( .A(n_254), .Y(n_291) );
AOI21x1_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_268), .Y(n_254) );
AO31x2_ASAP7_75t_L g279 ( .A1(n_255), .A2(n_280), .A3(n_286), .B(n_288), .Y(n_279) );
AO31x2_ASAP7_75t_L g531 ( .A1(n_255), .A2(n_532), .A3(n_538), .B(n_539), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_260), .B(n_263), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g285 ( .A(n_261), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_SL g526 ( .A(n_267), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_269), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g373 ( .A(n_269), .Y(n_373) );
INVx2_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
BUFx2_ASAP7_75t_L g313 ( .A(n_270), .Y(n_313) );
OR2x2_ASAP7_75t_L g379 ( .A(n_270), .B(n_279), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_270), .B(n_279), .Y(n_412) );
INVx2_ASAP7_75t_L g360 ( .A(n_277), .Y(n_360) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_290), .Y(n_277) );
OR2x2_ASAP7_75t_L g347 ( .A(n_278), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g425 ( .A(n_278), .Y(n_425) );
INVx1_ASAP7_75t_L g308 ( .A(n_279), .Y(n_308) );
INVx1_ASAP7_75t_L g316 ( .A(n_279), .Y(n_316) );
INVx1_ASAP7_75t_L g331 ( .A(n_279), .Y(n_331) );
AO31x2_ASAP7_75t_L g522 ( .A1(n_286), .A2(n_523), .A3(n_524), .B(n_528), .Y(n_522) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_SL g599 ( .A(n_287), .Y(n_599) );
OR2x2_ASAP7_75t_L g435 ( .A(n_290), .B(n_412), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_291), .B(n_307), .Y(n_348) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_291), .Y(n_350) );
OR2x2_ASAP7_75t_L g449 ( .A(n_291), .B(n_373), .Y(n_449) );
INVxp67_ASAP7_75t_L g473 ( .A(n_291), .Y(n_473) );
INVx2_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
NAND2x1_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_294), .B(n_335), .Y(n_402) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g351 ( .A(n_296), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g464 ( .A(n_297), .Y(n_464) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g493 ( .A(n_298), .B(n_326), .Y(n_493) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g419 ( .A(n_299), .B(n_326), .Y(n_419) );
AOI21x1_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B(n_302), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_310), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_306), .B(n_342), .Y(n_456) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx2_ASAP7_75t_L g320 ( .A(n_307), .Y(n_320) );
AND2x2_ASAP7_75t_L g370 ( .A(n_307), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_307), .B(n_364), .Y(n_413) );
OR2x2_ASAP7_75t_L g485 ( .A(n_307), .B(n_372), .Y(n_485) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g405 ( .A(n_311), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx2_ASAP7_75t_L g396 ( .A(n_312), .Y(n_396) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g386 ( .A(n_315), .B(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_315), .Y(n_397) );
OR2x2_ASAP7_75t_L g448 ( .A(n_315), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g503 ( .A(n_315), .Y(n_503) );
AOI211xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B(n_327), .C(n_336), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g392 ( .A(n_320), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_320), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g465 ( .A(n_320), .B(n_342), .Y(n_465) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_323), .B(n_368), .Y(n_390) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_323), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g475 ( .A(n_323), .B(n_476), .Y(n_475) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx2_ASAP7_75t_L g418 ( .A(n_324), .Y(n_418) );
AND2x2_ASAP7_75t_L g446 ( .A(n_325), .B(n_374), .Y(n_446) );
INVx2_ASAP7_75t_L g469 ( .A(n_325), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_325), .B(n_367), .Y(n_501) );
AND2x4_ASAP7_75t_SL g455 ( .A(n_328), .B(n_333), .Y(n_455) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g408 ( .A(n_329), .B(n_334), .Y(n_408) );
OR2x2_ASAP7_75t_L g460 ( .A(n_329), .B(n_353), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_330), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_330), .B(n_342), .Y(n_496) );
BUFx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g444 ( .A(n_331), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g427 ( .A(n_333), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_333), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g477 ( .A(n_334), .Y(n_477) );
BUFx2_ASAP7_75t_L g345 ( .A(n_335), .Y(n_345) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g463 ( .A(n_338), .B(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g387 ( .A(n_342), .Y(n_387) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_342), .Y(n_404) );
NAND3xp33_ASAP7_75t_SL g343 ( .A(n_344), .B(n_354), .C(n_369), .Y(n_343) );
AOI22xp33_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_346), .B1(n_349), .B2(n_351), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_351), .A2(n_377), .B1(n_458), .B2(n_461), .C1(n_463), .C2(n_465), .Y(n_457) );
AND2x2_ASAP7_75t_L g489 ( .A(n_352), .B(n_438), .Y(n_489) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g437 ( .A(n_353), .B(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_360), .B1(n_361), .B2(n_366), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx2_ASAP7_75t_SL g433 ( .A(n_357), .Y(n_433) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_365), .Y(n_361) );
AND2x2_ASAP7_75t_L g420 ( .A(n_362), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g378 ( .A(n_363), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g372 ( .A(n_364), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g487 ( .A(n_365), .Y(n_487) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_368), .B(n_464), .Y(n_483) );
INVx1_ASAP7_75t_L g500 ( .A(n_368), .Y(n_500) );
AOI222xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_374), .B1(n_375), .B2(n_377), .C1(n_380), .C2(n_381), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_376), .Y(n_380) );
AND2x2_ASAP7_75t_L g398 ( .A(n_376), .B(n_399), .Y(n_398) );
INVx3_ASAP7_75t_L g429 ( .A(n_376), .Y(n_429) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g393 ( .A(n_379), .Y(n_393) );
OR2x2_ASAP7_75t_L g462 ( .A(n_379), .B(n_443), .Y(n_462) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_391), .C(n_400), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI21xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_398), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_392), .A2(n_430), .B1(n_479), .B2(n_482), .C(n_484), .Y(n_478) );
AND2x4_ASAP7_75t_L g421 ( .A(n_393), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g452 ( .A(n_399), .Y(n_452) );
AOI211x1_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B(n_405), .C(n_409), .Y(n_400) );
INVxp67_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g470 ( .A(n_408), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_411), .B(n_459), .C(n_460), .Y(n_458) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g494 ( .A(n_412), .Y(n_494) );
NOR2x1_ASAP7_75t_L g414 ( .A(n_415), .B(n_466), .Y(n_414) );
NAND4xp25_ASAP7_75t_L g415 ( .A(n_416), .B(n_423), .C(n_445), .D(n_457), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
AND2x2_ASAP7_75t_L g476 ( .A(n_419), .B(n_477), .Y(n_476) );
AOI221x1_ASAP7_75t_L g445 ( .A1(n_421), .A2(n_446), .B1(n_447), .B2(n_450), .C(n_453), .Y(n_445) );
AND2x2_ASAP7_75t_L g471 ( .A(n_421), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g481 ( .A(n_422), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_430), .B2(n_434), .C(n_436), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_428), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_433), .A2(n_437), .B1(n_440), .B2(n_442), .Y(n_436) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_437), .A2(n_454), .B(n_456), .Y(n_453) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g459 ( .A(n_439), .Y(n_459) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_L g480 ( .A(n_449), .Y(n_480) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g499 ( .A1(n_462), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_478), .C(n_490), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_471), .B1(n_474), .B2(n_475), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g486 ( .A(n_473), .B(n_487), .Y(n_486) );
NAND2x1_ASAP7_75t_L g502 ( .A(n_473), .B(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_488), .Y(n_484) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_494), .B1(n_495), .B2(n_497), .C(n_499), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx3_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
INVx4_ASAP7_75t_L g809 ( .A(n_504), .Y(n_809) );
BUFx12f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g817 ( .A(n_506), .B(n_818), .Y(n_817) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_507), .B(n_830), .Y(n_829) );
NOR2x1p5_ASAP7_75t_L g507 ( .A(n_508), .B(n_719), .Y(n_507) );
NAND4xp75_ASAP7_75t_L g508 ( .A(n_509), .B(n_664), .C(n_684), .D(n_700), .Y(n_508) );
NOR2x1p5_ASAP7_75t_SL g509 ( .A(n_510), .B(n_634), .Y(n_509) );
NAND4xp75_ASAP7_75t_L g510 ( .A(n_511), .B(n_572), .C(n_611), .D(n_620), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_541), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_521), .Y(n_512) );
AND2x4_ASAP7_75t_L g744 ( .A(n_513), .B(n_671), .Y(n_744) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_514), .Y(n_587) );
INVx2_ASAP7_75t_L g605 ( .A(n_514), .Y(n_605) );
AND2x2_ASAP7_75t_L g628 ( .A(n_514), .B(n_590), .Y(n_628) );
OR2x2_ASAP7_75t_L g683 ( .A(n_514), .B(n_522), .Y(n_683) );
AND2x2_ASAP7_75t_L g601 ( .A(n_521), .B(n_602), .Y(n_601) );
AND2x4_ASAP7_75t_L g751 ( .A(n_521), .B(n_628), .Y(n_751) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_530), .Y(n_521) );
OR2x2_ASAP7_75t_L g588 ( .A(n_522), .B(n_589), .Y(n_588) );
BUFx2_ASAP7_75t_L g619 ( .A(n_522), .Y(n_619) );
AND2x2_ASAP7_75t_L g625 ( .A(n_522), .B(n_531), .Y(n_625) );
INVx1_ASAP7_75t_L g643 ( .A(n_522), .Y(n_643) );
INVx2_ASAP7_75t_L g672 ( .A(n_522), .Y(n_672) );
INVx3_ASAP7_75t_L g648 ( .A(n_530), .Y(n_648) );
INVx2_ASAP7_75t_L g653 ( .A(n_530), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_530), .B(n_604), .Y(n_658) );
AND2x2_ASAP7_75t_L g681 ( .A(n_530), .B(n_660), .Y(n_681) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_530), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_530), .B(n_736), .Y(n_735) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g670 ( .A(n_531), .Y(n_670) );
AND2x2_ASAP7_75t_L g718 ( .A(n_531), .B(n_672), .Y(n_718) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_554), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_543), .B(n_662), .Y(n_709) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2x1p5_ASAP7_75t_L g706 ( .A(n_544), .B(n_662), .Y(n_706) );
INVx1_ASAP7_75t_L g807 ( .A(n_544), .Y(n_807) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g757 ( .A(n_545), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g610 ( .A(n_546), .Y(n_610) );
OR2x2_ASAP7_75t_L g691 ( .A(n_546), .B(n_565), .Y(n_691) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g633 ( .A(n_547), .Y(n_633) );
AND2x4_ASAP7_75t_L g639 ( .A(n_547), .B(n_640), .Y(n_639) );
AOI32xp33_ASAP7_75t_L g777 ( .A1(n_554), .A2(n_680), .A3(n_778), .B1(n_780), .B2(n_781), .Y(n_777) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g726 ( .A(n_555), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_564), .Y(n_555) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_556), .Y(n_574) );
OR2x2_ASAP7_75t_L g608 ( .A(n_556), .B(n_566), .Y(n_608) );
INVx1_ASAP7_75t_L g623 ( .A(n_556), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_556), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g638 ( .A(n_556), .Y(n_638) );
INVx2_ASAP7_75t_L g663 ( .A(n_556), .Y(n_663) );
AND2x2_ASAP7_75t_L g782 ( .A(n_556), .B(n_576), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_564), .B(n_615), .Y(n_702) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g575 ( .A(n_566), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g631 ( .A(n_566), .Y(n_631) );
INVx2_ASAP7_75t_L g640 ( .A(n_566), .Y(n_640) );
AND2x4_ASAP7_75t_L g662 ( .A(n_566), .B(n_663), .Y(n_662) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_566), .Y(n_754) );
AOI22x1_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_583), .B1(n_601), .B2(n_606), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NAND4xp25_ASAP7_75t_L g731 ( .A(n_575), .B(n_732), .C(n_733), .D(n_734), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_575), .B(n_632), .Y(n_762) );
INVx4_ASAP7_75t_SL g615 ( .A(n_576), .Y(n_615) );
BUFx2_ASAP7_75t_L g678 ( .A(n_576), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_576), .B(n_623), .Y(n_741) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g703 ( .A(n_585), .B(n_652), .Y(n_703) );
NOR2x1_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_L g626 ( .A(n_589), .B(n_604), .Y(n_626) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_590), .B(n_605), .Y(n_650) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B(n_600), .Y(n_590) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_591), .A2(n_592), .B(n_600), .Y(n_645) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_596), .B(n_599), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_602), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g668 ( .A(n_602), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g707 ( .A(n_603), .B(n_625), .Y(n_707) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g750 ( .A(n_605), .B(n_660), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_606), .A2(n_723), .B1(n_725), .B2(n_728), .C(n_730), .Y(n_722) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx2_ASAP7_75t_L g616 ( .A(n_608), .Y(n_616) );
OR2x2_ASAP7_75t_L g716 ( .A(n_608), .B(n_655), .Y(n_716) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_617), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_612), .A2(n_738), .B1(n_742), .B2(n_745), .Y(n_737) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_616), .Y(n_612) );
AND2x4_ASAP7_75t_L g661 ( .A(n_613), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g773 ( .A(n_613), .B(n_691), .Y(n_773) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x4_ASAP7_75t_L g621 ( .A(n_615), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g637 ( .A(n_615), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g696 ( .A(n_615), .B(n_633), .Y(n_696) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_615), .Y(n_713) );
INVx1_ASAP7_75t_L g727 ( .A(n_615), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_615), .B(n_640), .Y(n_770) );
AND2x4_ASAP7_75t_L g677 ( .A(n_616), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g675 ( .A(n_618), .Y(n_675) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_619), .B(n_660), .Y(n_659) );
NAND2x1_ASAP7_75t_L g779 ( .A(n_619), .B(n_681), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_624), .B1(n_627), .B2(n_629), .Y(n_620) );
AND2x2_ASAP7_75t_L g646 ( .A(n_621), .B(n_639), .Y(n_646) );
INVx1_ASAP7_75t_L g687 ( .A(n_621), .Y(n_687) );
AND2x2_ASAP7_75t_L g794 ( .A(n_621), .B(n_655), .Y(n_794) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x4_ASAP7_75t_SL g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AND2x2_ASAP7_75t_L g627 ( .A(n_625), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g767 ( .A(n_625), .Y(n_767) );
AND2x2_ASAP7_75t_L g784 ( .A(n_625), .B(n_644), .Y(n_784) );
AND2x2_ASAP7_75t_L g800 ( .A(n_625), .B(n_750), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_626), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g723 ( .A(n_626), .B(n_724), .Y(n_723) );
OAI22xp33_ASAP7_75t_L g730 ( .A1(n_626), .A2(n_716), .B1(n_731), .B2(n_735), .Y(n_730) );
INVx1_ASAP7_75t_L g686 ( .A(n_628), .Y(n_686) );
AND2x2_ASAP7_75t_L g717 ( .A(n_628), .B(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_628), .B(n_724), .Y(n_746) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g752 ( .A(n_632), .B(n_753), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_632), .A2(n_656), .B1(n_761), .B2(n_763), .Y(n_760) );
INVx3_ASAP7_75t_L g655 ( .A(n_633), .Y(n_655) );
AND2x2_ASAP7_75t_L g787 ( .A(n_633), .B(n_640), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_651), .Y(n_634) );
AOI32xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_641), .A3(n_644), .B1(n_646), .B2(n_647), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_638), .Y(n_733) );
INVx1_ASAP7_75t_L g758 ( .A(n_638), .Y(n_758) );
INVx3_ASAP7_75t_L g714 ( .A(n_639), .Y(n_714) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g789 ( .A1(n_642), .A2(n_790), .B1(n_791), .B2(n_792), .C(n_793), .Y(n_789) );
BUFx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g766 ( .A(n_644), .B(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_L g802 ( .A(n_644), .B(n_763), .Y(n_802) );
BUFx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g660 ( .A(n_645), .Y(n_660) );
NAND2x1p5_ASAP7_75t_L g674 ( .A(n_647), .B(n_675), .Y(n_674) );
AO22x1_ASAP7_75t_L g704 ( .A1(n_647), .A2(n_705), .B1(n_707), .B2(n_708), .Y(n_704) );
NAND2x1p5_ASAP7_75t_L g808 ( .A(n_647), .B(n_675), .Y(n_808) );
AND2x4_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx2_ASAP7_75t_L g724 ( .A(n_648), .Y(n_724) );
INVx1_ASAP7_75t_L g734 ( .A(n_648), .Y(n_734) );
AND2x2_ASAP7_75t_L g654 ( .A(n_649), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVxp67_ASAP7_75t_SL g736 ( .A(n_650), .Y(n_736) );
INVx1_ASAP7_75t_L g776 ( .A(n_650), .Y(n_776) );
A2O1A1Ixp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B(n_656), .C(n_661), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2x1p5_ASAP7_75t_L g763 ( .A(n_653), .B(n_683), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_654), .B(n_713), .Y(n_790) );
AOI31xp33_ASAP7_75t_L g673 ( .A1(n_655), .A2(n_674), .A3(n_676), .B(n_679), .Y(n_673) );
INVx4_ASAP7_75t_L g732 ( .A(n_655), .Y(n_732) );
OR2x2_ASAP7_75t_L g769 ( .A(n_655), .B(n_770), .Y(n_769) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
AND2x4_ASAP7_75t_L g671 ( .A(n_660), .B(n_672), .Y(n_671) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_662), .Y(n_667) );
AND2x2_ASAP7_75t_L g698 ( .A(n_662), .B(n_696), .Y(n_698) );
NOR2xp67_ASAP7_75t_L g664 ( .A(n_665), .B(n_673), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g791 ( .A(n_668), .Y(n_791) );
INVx1_ASAP7_75t_L g699 ( .A(n_669), .Y(n_699) );
AND2x4_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g729 ( .A(n_670), .Y(n_729) );
AND2x2_ASAP7_75t_L g728 ( .A(n_671), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI322xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .A3(n_688), .B1(n_692), .B2(n_695), .C1(n_697), .C2(n_699), .Y(n_685) );
INVxp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI211x1_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B(n_704), .C(n_710), .Y(n_700) );
INVx1_ASAP7_75t_L g805 ( .A(n_701), .Y(n_805) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g759 ( .A(n_703), .Y(n_759) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OA21x2_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_715), .B(n_717), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx2_ASAP7_75t_L g780 ( .A(n_714), .Y(n_780) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp33_ASAP7_75t_L g775 ( .A(n_718), .B(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_788), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_755), .C(n_771), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_737), .C(n_747), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_724), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI21xp33_ASAP7_75t_L g783 ( .A1(n_728), .A2(n_784), .B(n_785), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_732), .B(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_732), .B(n_782), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_733), .B(n_807), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_734), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OAI21xp5_ASAP7_75t_L g793 ( .A1(n_744), .A2(n_794), .B(n_795), .Y(n_793) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_751), .B(n_752), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OAI211xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_759), .B(n_760), .C(n_764), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_765), .B(n_768), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_SL g774 ( .A(n_766), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_770), .Y(n_792) );
OAI211xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_774), .B(n_777), .C(n_783), .Y(n_771) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_782), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g803 ( .A(n_782), .Y(n_803) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g799 ( .A(n_787), .Y(n_799) );
NOR3xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_797), .C(n_804), .Y(n_788) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AOI21xp33_ASAP7_75t_SL g797 ( .A1(n_798), .A2(n_801), .B(n_803), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AOI21xp33_ASAP7_75t_R g804 ( .A1(n_805), .A2(n_806), .B(n_808), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
INVx6_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
BUFx10_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
OR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_824), .Y(n_819) );
INVxp67_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
BUFx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
INVx8_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
endmodule