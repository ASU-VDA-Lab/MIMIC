module real_aes_7869_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_723, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_723;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_686;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g448 ( .A1(n_0), .A2(n_186), .B(n_449), .C(n_452), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_1), .B(n_443), .Y(n_453) );
INVx1_ASAP7_75t_L g684 ( .A(n_2), .Y(n_684) );
INVx1_ASAP7_75t_L g221 ( .A(n_3), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_4), .B(n_138), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_5), .A2(n_438), .B(n_526), .Y(n_525) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_6), .A2(n_161), .B(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_7), .A2(n_37), .B1(n_131), .B2(n_155), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_8), .B(n_161), .Y(n_233) );
AND2x6_ASAP7_75t_L g146 ( .A(n_9), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_10), .A2(n_146), .B(n_429), .C(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_11), .B(n_38), .Y(n_685) );
INVx1_ASAP7_75t_L g127 ( .A(n_12), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_13), .B(n_136), .Y(n_169) );
INVx1_ASAP7_75t_L g213 ( .A(n_14), .Y(n_213) );
AOI222xp33_ASAP7_75t_L g101 ( .A1(n_15), .A2(n_102), .B1(n_689), .B2(n_698), .C1(n_714), .C2(n_720), .Y(n_101) );
OAI22xp33_ASAP7_75t_SL g700 ( .A1(n_15), .A2(n_701), .B1(n_706), .B2(n_707), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_15), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_16), .B(n_138), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_17), .B(n_162), .Y(n_200) );
AO32x2_ASAP7_75t_L g183 ( .A1(n_18), .A2(n_160), .A3(n_161), .B1(n_184), .B2(n_188), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_19), .B(n_131), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_20), .B(n_162), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_21), .A2(n_53), .B1(n_131), .B2(n_155), .Y(n_187) );
AOI22xp33_ASAP7_75t_SL g158 ( .A1(n_22), .A2(n_80), .B1(n_131), .B2(n_136), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_23), .B(n_131), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_24), .A2(n_160), .B(n_429), .C(n_476), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_25), .A2(n_160), .B(n_429), .C(n_491), .Y(n_490) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_26), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_27), .B(n_123), .Y(n_242) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_28), .A2(n_89), .B1(n_107), .B2(n_108), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_28), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_29), .A2(n_438), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_30), .B(n_123), .Y(n_148) );
INVx2_ASAP7_75t_L g133 ( .A(n_31), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_32), .A2(n_435), .B(n_461), .C(n_462), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_33), .B(n_131), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_34), .B(n_123), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g704 ( .A1(n_35), .A2(n_42), .B1(n_419), .B2(n_705), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_35), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_36), .B(n_171), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_39), .B(n_474), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_40), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_41), .B(n_138), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g113 ( .A1(n_42), .A2(n_114), .B1(n_419), .B2(n_420), .Y(n_113) );
INVx1_ASAP7_75t_L g419 ( .A(n_42), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_43), .B(n_438), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_44), .A2(n_435), .B(n_461), .C(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_45), .B(n_131), .Y(n_228) );
INVx1_ASAP7_75t_L g450 ( .A(n_46), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_47), .A2(n_88), .B1(n_155), .B2(n_156), .Y(n_154) );
INVx1_ASAP7_75t_L g513 ( .A(n_48), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_49), .B(n_131), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_50), .B(n_131), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_51), .B(n_438), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_52), .B(n_219), .Y(n_232) );
AOI22xp33_ASAP7_75t_SL g204 ( .A1(n_54), .A2(n_58), .B1(n_131), .B2(n_136), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_55), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_56), .B(n_131), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_57), .B(n_131), .Y(n_241) );
INVx1_ASAP7_75t_L g147 ( .A(n_59), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_60), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_61), .B(n_443), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_62), .A2(n_216), .B(n_219), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_63), .B(n_131), .Y(n_222) );
INVx1_ASAP7_75t_L g126 ( .A(n_64), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_65), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_66), .B(n_138), .Y(n_466) );
AO32x2_ASAP7_75t_L g152 ( .A1(n_67), .A2(n_153), .A3(n_159), .B1(n_160), .B2(n_161), .Y(n_152) );
AOI22xp5_ASAP7_75t_SL g103 ( .A1(n_68), .A2(n_104), .B1(n_682), .B2(n_686), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_69), .B(n_139), .Y(n_503) );
INVx1_ASAP7_75t_L g240 ( .A(n_70), .Y(n_240) );
INVx1_ASAP7_75t_L g134 ( .A(n_71), .Y(n_134) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_72), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_73), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_74), .B(n_465), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g428 ( .A1(n_75), .A2(n_429), .B(n_431), .C(n_435), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_76), .B(n_136), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g527 ( .A(n_77), .Y(n_527) );
INVx1_ASAP7_75t_L g693 ( .A(n_78), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_79), .B(n_464), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_81), .B(n_155), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_82), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_83), .B(n_136), .Y(n_143) );
INVx2_ASAP7_75t_L g124 ( .A(n_84), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_85), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_86), .B(n_157), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_87), .B(n_136), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_89), .Y(n_107) );
INVx2_ASAP7_75t_L g112 ( .A(n_90), .Y(n_112) );
OR2x2_ASAP7_75t_L g697 ( .A(n_90), .B(n_682), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_91), .A2(n_100), .B1(n_136), .B2(n_137), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_92), .B(n_438), .Y(n_459) );
INVx1_ASAP7_75t_L g463 ( .A(n_93), .Y(n_463) );
INVxp67_ASAP7_75t_L g530 ( .A(n_94), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_95), .B(n_136), .Y(n_238) );
INVx1_ASAP7_75t_L g432 ( .A(n_96), .Y(n_432) );
INVx1_ASAP7_75t_L g499 ( .A(n_97), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_98), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g515 ( .A(n_99), .B(n_123), .Y(n_515) );
INVxp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_106), .B1(n_109), .B2(n_681), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g681 ( .A(n_111), .Y(n_681) );
AO22x2_ASAP7_75t_SL g111 ( .A1(n_112), .A2(n_113), .B1(n_421), .B2(n_680), .Y(n_111) );
INVx1_ASAP7_75t_L g680 ( .A(n_112), .Y(n_680) );
NOR2x2_ASAP7_75t_L g688 ( .A(n_112), .B(n_682), .Y(n_688) );
INVx1_ASAP7_75t_L g420 ( .A(n_114), .Y(n_420) );
OAI22xp5_ASAP7_75t_SL g702 ( .A1(n_114), .A2(n_420), .B1(n_703), .B2(n_704), .Y(n_702) );
OR2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_340), .Y(n_114) );
NAND3xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_289), .C(n_331), .Y(n_115) );
AOI211xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_194), .B(n_243), .C(n_265), .Y(n_116) );
OAI211xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_149), .B(n_177), .C(n_189), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_119), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g352 ( .A(n_119), .B(n_269), .Y(n_352) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g254 ( .A(n_120), .B(n_180), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_120), .B(n_165), .Y(n_371) );
INVx1_ASAP7_75t_L g389 ( .A(n_120), .Y(n_389) );
AND2x2_ASAP7_75t_L g398 ( .A(n_120), .B(n_286), .Y(n_398) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g281 ( .A(n_121), .B(n_165), .Y(n_281) );
AND2x2_ASAP7_75t_L g339 ( .A(n_121), .B(n_286), .Y(n_339) );
INVx1_ASAP7_75t_L g383 ( .A(n_121), .Y(n_383) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g260 ( .A(n_122), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g268 ( .A(n_122), .Y(n_268) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_122), .Y(n_308) );
OA21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_128), .B(n_148), .Y(n_122) );
INVx2_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_123), .A2(n_166), .B(n_176), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_123), .A2(n_459), .B(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g482 ( .A(n_123), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_123), .A2(n_510), .B(n_511), .Y(n_509) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x2_ASAP7_75t_L g162 ( .A(n_124), .B(n_125), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_141), .B(n_146), .Y(n_128) );
O2A1O1Ixp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_134), .B(n_135), .C(n_138), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_131), .Y(n_434) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_132), .Y(n_156) );
AND2x6_ASAP7_75t_L g429 ( .A(n_132), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g137 ( .A(n_133), .Y(n_137) );
INVx1_ASAP7_75t_L g220 ( .A(n_133), .Y(n_220) );
INVx2_ASAP7_75t_L g214 ( .A(n_136), .Y(n_214) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_138), .A2(n_228), .B(n_229), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_138), .A2(n_237), .B(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_138), .B(n_530), .Y(n_529) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OAI22xp5_ASAP7_75t_SL g153 ( .A1(n_139), .A2(n_154), .B1(n_157), .B2(n_158), .Y(n_153) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_140), .Y(n_145) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
INVx1_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
INVx1_ASAP7_75t_L g430 ( .A(n_140), .Y(n_430) );
AND2x2_ASAP7_75t_L g439 ( .A(n_140), .B(n_220), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g216 ( .A(n_144), .Y(n_216) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g465 ( .A(n_145), .Y(n_465) );
BUFx3_ASAP7_75t_L g160 ( .A(n_146), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g166 ( .A1(n_146), .A2(n_167), .B(n_172), .Y(n_166) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_146), .A2(n_212), .B(n_217), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_146), .A2(n_227), .B(n_230), .Y(n_226) );
INVx4_ASAP7_75t_SL g436 ( .A(n_146), .Y(n_436) );
AND2x4_ASAP7_75t_L g438 ( .A(n_146), .B(n_439), .Y(n_438) );
NAND2x1p5_ASAP7_75t_L g500 ( .A(n_146), .B(n_439), .Y(n_500) );
INVxp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_163), .Y(n_150) );
AND2x2_ASAP7_75t_L g247 ( .A(n_151), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g280 ( .A(n_151), .Y(n_280) );
OR2x2_ASAP7_75t_L g406 ( .A(n_151), .B(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_151), .B(n_165), .Y(n_410) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
INVx1_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
AND2x2_ASAP7_75t_L g269 ( .A(n_152), .B(n_182), .Y(n_269) );
AND2x2_ASAP7_75t_L g309 ( .A(n_152), .B(n_183), .Y(n_309) );
INVx2_ASAP7_75t_L g452 ( .A(n_156), .Y(n_452) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_156), .Y(n_467) );
INVx2_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_157), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_157), .A2(n_186), .B1(n_203), .B2(n_204), .Y(n_202) );
INVx4_ASAP7_75t_L g451 ( .A(n_157), .Y(n_451) );
INVx1_ASAP7_75t_L g479 ( .A(n_159), .Y(n_479) );
NAND3xp33_ASAP7_75t_L g201 ( .A(n_160), .B(n_202), .C(n_205), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_160), .A2(n_236), .B(n_239), .Y(n_235) );
INVx4_ASAP7_75t_L g205 ( .A(n_161), .Y(n_205) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_161), .A2(n_226), .B(n_233), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_161), .A2(n_489), .B(n_490), .Y(n_488) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_161), .Y(n_524) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
INVxp67_ASAP7_75t_L g351 ( .A(n_163), .Y(n_351) );
AND2x4_ASAP7_75t_L g376 ( .A(n_163), .B(n_269), .Y(n_376) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_164), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g181 ( .A(n_165), .B(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g255 ( .A(n_165), .B(n_183), .Y(n_255) );
INVx1_ASAP7_75t_L g261 ( .A(n_165), .Y(n_261) );
INVx2_ASAP7_75t_L g287 ( .A(n_165), .Y(n_287) );
AND2x2_ASAP7_75t_L g303 ( .A(n_165), .B(n_304), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_170), .Y(n_167) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .Y(n_172) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_175), .A2(n_218), .B(n_240), .C(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_178), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_181), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx2_ASAP7_75t_L g258 ( .A(n_180), .Y(n_258) );
AND2x2_ASAP7_75t_L g366 ( .A(n_180), .B(n_182), .Y(n_366) );
AND2x2_ASAP7_75t_L g283 ( .A(n_181), .B(n_268), .Y(n_283) );
AND2x2_ASAP7_75t_L g382 ( .A(n_181), .B(n_383), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g304 ( .A(n_182), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g407 ( .A(n_182), .B(n_268), .Y(n_407) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx2_ASAP7_75t_L g193 ( .A(n_183), .Y(n_193) );
AND2x2_ASAP7_75t_L g286 ( .A(n_183), .B(n_287), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_186), .A2(n_218), .B(n_221), .C(n_222), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_186), .A2(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g210 ( .A(n_188), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_188), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_193), .Y(n_190) );
AND2x2_ASAP7_75t_L g332 ( .A(n_191), .B(n_267), .Y(n_332) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_192), .B(n_268), .Y(n_317) );
INVx2_ASAP7_75t_L g316 ( .A(n_193), .Y(n_316) );
OAI222xp33_ASAP7_75t_L g320 ( .A1(n_193), .A2(n_260), .B1(n_321), .B2(n_323), .C1(n_324), .C2(n_327), .Y(n_320) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_206), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g245 ( .A(n_198), .Y(n_245) );
OR2x2_ASAP7_75t_L g356 ( .A(n_198), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx3_ASAP7_75t_L g278 ( .A(n_199), .Y(n_278) );
NOR2x1_ASAP7_75t_L g329 ( .A(n_199), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g335 ( .A(n_199), .B(n_249), .Y(n_335) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g296 ( .A(n_200), .Y(n_296) );
AO21x1_ASAP7_75t_L g295 ( .A1(n_202), .A2(n_205), .B(n_296), .Y(n_295) );
AO21x2_ASAP7_75t_L g426 ( .A1(n_205), .A2(n_427), .B(n_440), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_205), .B(n_441), .Y(n_440) );
INVx3_ASAP7_75t_L g443 ( .A(n_205), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_205), .B(n_469), .Y(n_468) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_205), .A2(n_498), .B(n_505), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_206), .A2(n_299), .B1(n_338), .B2(n_339), .Y(n_337) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_224), .Y(n_206) );
INVx3_ASAP7_75t_L g271 ( .A(n_207), .Y(n_271) );
OR2x2_ASAP7_75t_L g404 ( .A(n_207), .B(n_280), .Y(n_404) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g277 ( .A(n_208), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g293 ( .A(n_208), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g301 ( .A(n_208), .B(n_249), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_208), .B(n_225), .Y(n_357) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g248 ( .A(n_209), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g252 ( .A(n_209), .B(n_225), .Y(n_252) );
AND2x2_ASAP7_75t_L g328 ( .A(n_209), .B(n_275), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_209), .B(n_234), .Y(n_368) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_223), .Y(n_209) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_210), .A2(n_235), .B(n_242), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .C(n_216), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_214), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_214), .A2(n_503), .B(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g431 ( .A1(n_216), .A2(n_432), .B(n_433), .C(n_434), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_218), .A2(n_477), .B(n_478), .Y(n_476) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_224), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g284 ( .A(n_224), .B(n_245), .Y(n_284) );
AND2x2_ASAP7_75t_L g288 ( .A(n_224), .B(n_278), .Y(n_288) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_234), .Y(n_224) );
INVx3_ASAP7_75t_L g249 ( .A(n_225), .Y(n_249) );
AND2x2_ASAP7_75t_L g274 ( .A(n_225), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g409 ( .A(n_225), .B(n_392), .Y(n_409) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
INVx2_ASAP7_75t_L g275 ( .A(n_234), .Y(n_275) );
AND2x2_ASAP7_75t_L g319 ( .A(n_234), .B(n_295), .Y(n_319) );
INVx1_ASAP7_75t_L g362 ( .A(n_234), .Y(n_362) );
OR2x2_ASAP7_75t_L g393 ( .A(n_234), .B(n_295), .Y(n_393) );
AND2x2_ASAP7_75t_L g413 ( .A(n_234), .B(n_249), .Y(n_413) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_246), .B(n_250), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g251 ( .A(n_245), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_245), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g370 ( .A(n_247), .Y(n_370) );
INVx2_ASAP7_75t_SL g264 ( .A(n_248), .Y(n_264) );
AND2x2_ASAP7_75t_L g384 ( .A(n_248), .B(n_278), .Y(n_384) );
INVx2_ASAP7_75t_L g330 ( .A(n_249), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_249), .B(n_362), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_253), .B1(n_256), .B2(n_262), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_252), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g418 ( .A(n_252), .Y(n_418) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g343 ( .A(n_254), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_254), .B(n_286), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_255), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g359 ( .A(n_255), .B(n_308), .Y(n_359) );
INVx2_ASAP7_75t_L g415 ( .A(n_255), .Y(n_415) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g285 ( .A(n_258), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_258), .B(n_303), .Y(n_336) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_260), .B(n_280), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g397 ( .A(n_263), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_SL g347 ( .A1(n_264), .A2(n_348), .B(n_350), .C(n_353), .Y(n_347) );
OR2x2_ASAP7_75t_L g374 ( .A(n_264), .B(n_278), .Y(n_374) );
OAI221xp5_ASAP7_75t_SL g265 ( .A1(n_266), .A2(n_270), .B1(n_272), .B2(n_279), .C(n_282), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_267), .B(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_267), .B(n_316), .Y(n_323) );
AND2x2_ASAP7_75t_L g365 ( .A(n_267), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g401 ( .A(n_267), .Y(n_401) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
INVx1_ASAP7_75t_L g305 ( .A(n_268), .Y(n_305) );
NOR2xp67_ASAP7_75t_L g325 ( .A(n_271), .B(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_L g379 ( .A(n_271), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_271), .B(n_319), .Y(n_395) );
INVx2_ASAP7_75t_L g381 ( .A(n_272), .Y(n_381) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g322 ( .A(n_274), .B(n_293), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_274), .A2(n_290), .B(n_332), .C(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g300 ( .A(n_275), .B(n_295), .Y(n_300) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_279), .B(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
OR2x2_ASAP7_75t_L g348 ( .A(n_280), .B(n_349), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_285), .B2(n_288), .Y(n_282) );
INVx1_ASAP7_75t_L g402 ( .A(n_284), .Y(n_402) );
INVx1_ASAP7_75t_L g349 ( .A(n_286), .Y(n_349) );
INVx1_ASAP7_75t_L g400 ( .A(n_288), .Y(n_400) );
AOI211xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_293), .B(n_297), .C(n_320), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g312 ( .A(n_292), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g363 ( .A(n_293), .Y(n_363) );
AND2x2_ASAP7_75t_L g412 ( .A(n_293), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI21xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_302), .B(n_310), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g326 ( .A(n_300), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_300), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g318 ( .A(n_301), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g394 ( .A(n_301), .Y(n_394) );
OAI32xp33_ASAP7_75t_L g405 ( .A1(n_301), .A2(n_353), .A3(n_360), .B1(n_401), .B2(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_SL g302 ( .A(n_303), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_SL g373 ( .A(n_303), .Y(n_373) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g313 ( .A(n_309), .Y(n_313) );
OAI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B(n_318), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g385 ( .A1(n_312), .A2(n_360), .B1(n_386), .B2(n_388), .Y(n_385) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_316), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g353 ( .A(n_319), .Y(n_353) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g346 ( .A(n_330), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B(n_337), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_339), .A2(n_381), .B1(n_382), .B2(n_384), .C(n_385), .Y(n_380) );
NAND5xp2_ASAP7_75t_L g340 ( .A(n_341), .B(n_364), .C(n_380), .D(n_390), .E(n_408), .Y(n_340) );
AOI211xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_344), .B(n_347), .C(n_354), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g411 ( .A(n_348), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_358), .B2(n_360), .Y(n_354) );
INVx1_ASAP7_75t_SL g387 ( .A(n_357), .Y(n_387) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI322xp33_ASAP7_75t_L g369 ( .A1(n_360), .A2(n_370), .A3(n_371), .B1(n_372), .B2(n_373), .C1(n_374), .C2(n_375), .Y(n_369) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g372 ( .A(n_362), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_362), .B(n_387), .Y(n_386) );
AOI211xp5_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_367), .B(n_369), .C(n_377), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_373), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_399) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_398), .B1(n_399), .B2(n_403), .C(n_405), .Y(n_390) );
OAI211xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_394), .B(n_395), .C(n_396), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g417 ( .A(n_393), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_411), .B2(n_412), .C(n_414), .Y(n_408) );
AOI21xp33_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B(n_417), .Y(n_414) );
NAND2x1p5_ASAP7_75t_L g421 ( .A(n_422), .B(n_623), .Y(n_421) );
AND4x1_ASAP7_75t_L g422 ( .A(n_423), .B(n_563), .C(n_578), .D(n_603), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g423 ( .A(n_424), .B(n_536), .Y(n_423) );
OAI21xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_454), .B(n_516), .Y(n_424) );
AND2x2_ASAP7_75t_L g566 ( .A(n_425), .B(n_471), .Y(n_566) );
AND2x2_ASAP7_75t_L g579 ( .A(n_425), .B(n_470), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_425), .B(n_455), .Y(n_629) );
INVx1_ASAP7_75t_L g633 ( .A(n_425), .Y(n_633) );
AND2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_442), .Y(n_425) );
INVx2_ASAP7_75t_L g550 ( .A(n_426), .Y(n_550) );
BUFx2_ASAP7_75t_L g577 ( .A(n_426), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_437), .Y(n_427) );
INVx5_ASAP7_75t_L g447 ( .A(n_429), .Y(n_447) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
O2A1O1Ixp33_ASAP7_75t_SL g445 ( .A1(n_436), .A2(n_446), .B(n_447), .C(n_448), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_436), .A2(n_447), .B(n_527), .C(n_528), .Y(n_526) );
BUFx2_ASAP7_75t_L g474 ( .A(n_438), .Y(n_474) );
AND2x2_ASAP7_75t_L g517 ( .A(n_442), .B(n_471), .Y(n_517) );
INVx2_ASAP7_75t_L g533 ( .A(n_442), .Y(n_533) );
AND2x2_ASAP7_75t_L g542 ( .A(n_442), .B(n_470), .Y(n_542) );
AND2x2_ASAP7_75t_L g621 ( .A(n_442), .B(n_550), .Y(n_621) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_453), .Y(n_442) );
INVx2_ASAP7_75t_L g461 ( .A(n_447), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_483), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_455), .B(n_548), .Y(n_586) );
INVx1_ASAP7_75t_L g674 ( .A(n_455), .Y(n_674) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_470), .Y(n_455) );
AND2x2_ASAP7_75t_L g532 ( .A(n_456), .B(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g546 ( .A(n_456), .B(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_456), .Y(n_575) );
OR2x2_ASAP7_75t_L g607 ( .A(n_456), .B(n_549), .Y(n_607) );
AND2x2_ASAP7_75t_L g615 ( .A(n_456), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g648 ( .A(n_456), .B(n_617), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_456), .B(n_517), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_456), .B(n_577), .Y(n_673) );
AND2x2_ASAP7_75t_L g679 ( .A(n_456), .B(n_566), .Y(n_679) );
INVx5_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g539 ( .A(n_457), .Y(n_539) );
AND2x2_ASAP7_75t_L g569 ( .A(n_457), .B(n_549), .Y(n_569) );
AND2x2_ASAP7_75t_L g602 ( .A(n_457), .B(n_562), .Y(n_602) );
AND2x2_ASAP7_75t_L g622 ( .A(n_457), .B(n_471), .Y(n_622) );
AND2x2_ASAP7_75t_L g656 ( .A(n_457), .B(n_522), .Y(n_656) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_468), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B(n_466), .C(n_467), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_464), .A2(n_467), .B(n_513), .C(n_514), .Y(n_512) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g562 ( .A(n_470), .B(n_533), .Y(n_562) );
AND2x2_ASAP7_75t_L g573 ( .A(n_470), .B(n_569), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_470), .B(n_549), .Y(n_612) );
INVx2_ASAP7_75t_L g627 ( .A(n_470), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_470), .B(n_561), .Y(n_650) );
AND2x2_ASAP7_75t_L g669 ( .A(n_470), .B(n_621), .Y(n_669) );
INVx5_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_471), .Y(n_568) );
AND2x2_ASAP7_75t_L g576 ( .A(n_471), .B(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g617 ( .A(n_471), .B(n_533), .Y(n_617) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_480), .Y(n_471) );
AOI21xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_475), .B(n_479), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
AND2x2_ASAP7_75t_L g540 ( .A(n_485), .B(n_523), .Y(n_540) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_486), .B(n_497), .Y(n_520) );
OR2x2_ASAP7_75t_L g553 ( .A(n_486), .B(n_523), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_486), .B(n_523), .Y(n_558) );
AND2x2_ASAP7_75t_L g585 ( .A(n_486), .B(n_522), .Y(n_585) );
AND2x2_ASAP7_75t_L g637 ( .A(n_486), .B(n_496), .Y(n_637) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_487), .B(n_507), .Y(n_545) );
AND2x2_ASAP7_75t_L g581 ( .A(n_487), .B(n_497), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_494), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g571 ( .A(n_495), .B(n_553), .Y(n_571) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_507), .Y(n_495) );
OAI322xp33_ASAP7_75t_L g536 ( .A1(n_496), .A2(n_537), .A3(n_541), .B1(n_543), .B2(n_546), .C1(n_551), .C2(n_559), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_496), .B(n_522), .Y(n_544) );
OR2x2_ASAP7_75t_L g554 ( .A(n_496), .B(n_508), .Y(n_554) );
AND2x2_ASAP7_75t_L g556 ( .A(n_496), .B(n_508), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_496), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_496), .B(n_523), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_496), .B(n_652), .Y(n_651) );
INVx5_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_497), .B(n_540), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B(n_501), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_507), .B(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g534 ( .A(n_507), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_507), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g596 ( .A(n_507), .B(n_523), .Y(n_596) );
AOI211xp5_ASAP7_75t_SL g624 ( .A1(n_507), .A2(n_625), .B(n_628), .C(n_640), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_507), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g662 ( .A(n_507), .B(n_637), .Y(n_662) );
INVx5_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g590 ( .A(n_508), .B(n_523), .Y(n_590) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_508), .Y(n_599) );
AND2x2_ASAP7_75t_L g639 ( .A(n_508), .B(n_637), .Y(n_639) );
AND2x2_ASAP7_75t_SL g670 ( .A(n_508), .B(n_540), .Y(n_670) );
AND2x2_ASAP7_75t_L g677 ( .A(n_508), .B(n_636), .Y(n_677) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_515), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B1(n_532), .B2(n_534), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_517), .B(n_539), .Y(n_587) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g535 ( .A(n_520), .Y(n_535) );
OR2x2_ASAP7_75t_L g595 ( .A(n_520), .B(n_596), .Y(n_595) );
OAI221xp5_ASAP7_75t_SL g643 ( .A1(n_520), .A2(n_644), .B1(n_646), .B2(n_647), .C(n_649), .Y(n_643) );
INVx2_ASAP7_75t_L g582 ( .A(n_521), .Y(n_582) );
AND2x2_ASAP7_75t_L g555 ( .A(n_522), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g645 ( .A(n_522), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_522), .B(n_637), .Y(n_658) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVxp67_ASAP7_75t_L g600 ( .A(n_523), .Y(n_600) );
AND2x2_ASAP7_75t_L g636 ( .A(n_523), .B(n_637), .Y(n_636) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_531), .Y(n_523) );
AND2x2_ASAP7_75t_L g638 ( .A(n_532), .B(n_577), .Y(n_638) );
AND2x2_ASAP7_75t_L g548 ( .A(n_533), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_533), .B(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_SL g619 ( .A(n_535), .B(n_582), .Y(n_619) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g625 ( .A(n_538), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
OR2x2_ASAP7_75t_L g611 ( .A(n_539), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g676 ( .A(n_539), .B(n_621), .Y(n_676) );
INVx2_ASAP7_75t_L g609 ( .A(n_540), .Y(n_609) );
NAND4xp25_ASAP7_75t_SL g672 ( .A(n_541), .B(n_673), .C(n_674), .D(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_542), .B(n_606), .Y(n_641) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_SL g678 ( .A(n_545), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_SL g640 ( .A1(n_546), .A2(n_609), .B(n_613), .C(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g635 ( .A(n_548), .B(n_627), .Y(n_635) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_549), .Y(n_561) );
INVx1_ASAP7_75t_L g616 ( .A(n_549), .Y(n_616) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_550), .Y(n_593) );
AOI211xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_554), .B(n_555), .C(n_557), .Y(n_551) );
AND2x2_ASAP7_75t_L g572 ( .A(n_552), .B(n_556), .Y(n_572) );
OAI322xp33_ASAP7_75t_SL g610 ( .A1(n_552), .A2(n_611), .A3(n_613), .B1(n_614), .B2(n_618), .C1(n_619), .C2(n_620), .Y(n_610) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g632 ( .A(n_554), .B(n_558), .Y(n_632) );
INVx1_ASAP7_75t_L g613 ( .A(n_556), .Y(n_613) );
INVx1_ASAP7_75t_SL g631 ( .A(n_558), .Y(n_631) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AOI222xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_570), .B1(n_572), .B2(n_573), .C1(n_574), .C2(n_723), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_565), .B(n_567), .Y(n_564) );
OAI322xp33_ASAP7_75t_L g653 ( .A1(n_565), .A2(n_627), .A3(n_632), .B1(n_654), .B2(n_655), .C1(n_657), .C2(n_658), .Y(n_653) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_566), .A2(n_580), .B1(n_604), .B2(n_608), .C(n_610), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OAI222xp33_ASAP7_75t_L g583 ( .A1(n_571), .A2(n_584), .B1(n_586), .B2(n_587), .C1(n_588), .C2(n_591), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_573), .A2(n_580), .B1(n_650), .B2(n_651), .Y(n_649) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AOI211xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B(n_583), .C(n_594), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g659 ( .A1(n_580), .A2(n_617), .B(n_660), .C(n_663), .Y(n_659) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g589 ( .A(n_581), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_SL g652 ( .A(n_585), .Y(n_652) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_592), .B(n_617), .Y(n_646) );
BUFx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI21xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B(n_601), .Y(n_594) );
OAI221xp5_ASAP7_75t_SL g663 ( .A1(n_595), .A2(n_664), .B1(n_665), .B2(n_666), .C(n_667), .Y(n_663) );
INVxp33_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_599), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_606), .B(n_617), .Y(n_657) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
AND2x2_ASAP7_75t_L g668 ( .A(n_621), .B(n_627), .Y(n_668) );
AND4x1_ASAP7_75t_L g623 ( .A(n_624), .B(n_642), .C(n_659), .D(n_671), .Y(n_623) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI221xp5_ASAP7_75t_SL g628 ( .A1(n_629), .A2(n_630), .B1(n_632), .B2(n_633), .C(n_634), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B1(n_638), .B2(n_639), .Y(n_634) );
INVx1_ASAP7_75t_L g664 ( .A(n_635), .Y(n_664) );
INVx1_ASAP7_75t_SL g654 ( .A(n_639), .Y(n_654) );
NOR2xp33_ASAP7_75t_SL g642 ( .A(n_643), .B(n_653), .Y(n_642) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_655), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_662), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_671) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx3_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_695), .Y(n_690) );
NOR2xp33_ASAP7_75t_SL g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVx1_ASAP7_75t_SL g719 ( .A(n_692), .Y(n_719) );
INVx1_ASAP7_75t_L g718 ( .A(n_694), .Y(n_718) );
OA21x2_ASAP7_75t_L g721 ( .A1(n_694), .A2(n_709), .B(n_719), .Y(n_721) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g709 ( .A(n_697), .Y(n_709) );
INVx2_ASAP7_75t_L g713 ( .A(n_697), .Y(n_713) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_708), .B(n_710), .Y(n_699) );
INVx1_ASAP7_75t_L g707 ( .A(n_701), .Y(n_707) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
BUFx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_715), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
endmodule