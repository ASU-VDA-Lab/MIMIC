module fake_jpeg_14024_n_645 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_645);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_645;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_61),
.Y(n_197)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_64),
.B(n_72),
.Y(n_143)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_66),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_67),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_73),
.B(n_91),
.Y(n_136)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_78),
.B(n_80),
.Y(n_146)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_79),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_16),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_82),
.Y(n_180)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_83),
.Y(n_181)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_84),
.Y(n_186)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

CKINVDCx9p33_ASAP7_75t_R g151 ( 
.A(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_88),
.Y(n_214)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_89),
.Y(n_217)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_40),
.B(n_16),
.Y(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_94),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_38),
.Y(n_95)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_97),
.B(n_109),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_99),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

CKINVDCx6p67_ASAP7_75t_R g177 ( 
.A(n_100),
.Y(n_177)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_32),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_40),
.B(n_41),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_105),
.B(n_33),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_38),
.B(n_1),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_59),
.C(n_30),
.Y(n_133)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_53),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_25),
.Y(n_110)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_114),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

BUFx2_ASAP7_75t_SL g194 ( 
.A(n_117),
.Y(n_194)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_53),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_124),
.Y(n_166)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_25),
.Y(n_123)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

BUFx16f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_28),
.B(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_126),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_33),
.B(n_16),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_58),
.Y(n_128)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_133),
.B(n_162),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_36),
.B1(n_21),
.B2(n_55),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_135),
.A2(n_31),
.B1(n_30),
.B2(n_44),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_73),
.B(n_55),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_137),
.B(n_171),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_66),
.A2(n_58),
.B1(n_57),
.B2(n_54),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_142),
.A2(n_144),
.B1(n_201),
.B2(n_206),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_61),
.A2(n_57),
.B1(n_54),
.B2(n_52),
.Y(n_144)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_152),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_161),
.B(n_163),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_47),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_125),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_91),
.B(n_47),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_168),
.B(n_175),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_100),
.A2(n_28),
.B(n_50),
.C(n_46),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_170),
.A2(n_211),
.B(n_115),
.C(n_56),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_95),
.B(n_26),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_26),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_174),
.B(n_195),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_63),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_128),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_85),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_67),
.B(n_29),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_67),
.B(n_29),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_196),
.B(n_199),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_122),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_209),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_102),
.B(n_45),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_89),
.A2(n_57),
.B1(n_54),
.B2(n_52),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_102),
.B(n_45),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_212),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_104),
.A2(n_21),
.B1(n_36),
.B2(n_52),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_208),
.A2(n_21),
.B1(n_56),
.B2(n_4),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_117),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_108),
.A2(n_50),
.B(n_46),
.C(n_44),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_108),
.B(n_31),
.Y(n_212)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_60),
.Y(n_216)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_169),
.A2(n_82),
.B1(n_121),
.B2(n_116),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g329 ( 
.A1(n_218),
.A2(n_219),
.B1(n_223),
.B2(n_260),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_162),
.A2(n_81),
.B1(n_68),
.B2(n_112),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_220),
.A2(n_241),
.B1(n_272),
.B2(n_149),
.Y(n_319)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_222),
.Y(n_315)
);

AO22x1_ASAP7_75t_SL g223 ( 
.A1(n_130),
.A2(n_127),
.B1(n_115),
.B2(n_98),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_224),
.A2(n_269),
.B(n_288),
.Y(n_307)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_225),
.Y(n_326)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_227),
.Y(n_333)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_138),
.Y(n_229)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_229),
.Y(n_323)
);

BUFx4f_ASAP7_75t_L g230 ( 
.A(n_151),
.Y(n_230)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_230),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_160),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_231),
.B(n_232),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_166),
.Y(n_232)
);

CKINVDCx9p33_ASAP7_75t_R g234 ( 
.A(n_134),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_234),
.Y(n_301)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_236),
.Y(n_338)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_237),
.Y(n_343)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_239),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_144),
.A2(n_88),
.B1(n_71),
.B2(n_36),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_132),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_243),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_141),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_244),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_245),
.A2(n_250),
.B1(n_263),
.B2(n_281),
.Y(n_310)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_155),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_246),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_146),
.B(n_15),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_247),
.B(n_253),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_141),
.Y(n_249)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_249),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_56),
.B1(n_3),
.B2(n_5),
.Y(n_250)
);

NAND2xp33_ASAP7_75t_SL g251 ( 
.A(n_140),
.B(n_2),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_251),
.A2(n_224),
.B(n_288),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_136),
.B(n_15),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_172),
.B(n_2),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_254),
.B(n_259),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_143),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_273),
.Y(n_303)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_148),
.Y(n_258)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_159),
.B(n_2),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_215),
.A2(n_56),
.B1(n_8),
.B2(n_10),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_261),
.Y(n_318)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_262),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_215),
.A2(n_56),
.B1(n_8),
.B2(n_10),
.Y(n_263)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

INVx5_ASAP7_75t_L g311 ( 
.A(n_264),
.Y(n_311)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_165),
.Y(n_265)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_153),
.Y(n_266)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_267),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_134),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_268),
.B(n_271),
.Y(n_350)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_185),
.Y(n_270)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_158),
.B(n_6),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_201),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_156),
.B(n_6),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_176),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_274),
.Y(n_297)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_157),
.Y(n_275)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_275),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_179),
.B(n_12),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_278),
.Y(n_309)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_152),
.Y(n_278)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_217),
.Y(n_280)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_216),
.A2(n_12),
.B1(n_13),
.B2(n_164),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_149),
.A2(n_12),
.B1(n_13),
.B2(n_164),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_282),
.A2(n_177),
.B1(n_214),
.B2(n_180),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_156),
.B(n_13),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_251),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_147),
.B(n_13),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_285),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_147),
.B(n_192),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_191),
.Y(n_286)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_286),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_157),
.Y(n_287)
);

BUFx8_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_156),
.A2(n_206),
.B1(n_217),
.B2(n_200),
.Y(n_288)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_200),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_202),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_187),
.B(n_207),
.C(n_142),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_140),
.C(n_134),
.Y(n_300)
);

CKINVDCx12_ASAP7_75t_R g292 ( 
.A(n_154),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_292),
.Y(n_302)
);

BUFx12_ASAP7_75t_L g293 ( 
.A(n_154),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_293),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_300),
.A2(n_306),
.B(n_332),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_241),
.A2(n_223),
.B1(n_250),
.B2(n_170),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_308),
.A2(n_319),
.B1(n_322),
.B2(n_325),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_291),
.A2(n_202),
.B(n_187),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_312),
.A2(n_264),
.B(n_289),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_314),
.B(n_320),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_316),
.A2(n_335),
.B1(n_310),
.B2(n_318),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_248),
.B(n_173),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_223),
.A2(n_150),
.B1(n_203),
.B2(n_180),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_269),
.A2(n_150),
.B1(n_203),
.B2(n_214),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_255),
.B(n_173),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_226),
.B(n_167),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_346),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_245),
.A2(n_207),
.B1(n_139),
.B2(n_167),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_345),
.A2(n_348),
.B1(n_349),
.B2(n_177),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_240),
.B(n_177),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_279),
.A2(n_284),
.B1(n_229),
.B2(n_242),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_234),
.A2(n_184),
.B1(n_182),
.B2(n_194),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_228),
.B(n_184),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_352),
.B(n_233),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_354),
.B(n_356),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_279),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_370),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_235),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_222),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_357),
.B(n_358),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_309),
.B(n_221),
.Y(n_358)
);

INVx13_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_359),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_303),
.B(n_277),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_360),
.B(n_365),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_361),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_362),
.A2(n_338),
.B(n_343),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_306),
.A2(n_289),
.B(n_285),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_363),
.A2(n_374),
.B(n_386),
.Y(n_422)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_364),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_270),
.Y(n_365)
);

INVxp67_ASAP7_75t_R g366 ( 
.A(n_352),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_366),
.B(n_368),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_319),
.A2(n_227),
.B1(n_266),
.B2(n_275),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_367),
.A2(n_379),
.B1(n_390),
.B2(n_340),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_280),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_290),
.Y(n_370)
);

INVx13_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_371),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_331),
.B(n_261),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_372),
.B(n_375),
.Y(n_415)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_373),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_307),
.A2(n_225),
.B1(n_256),
.B2(n_267),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_296),
.B(n_256),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_243),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_376),
.B(n_377),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_298),
.B(n_304),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_322),
.A2(n_252),
.B1(n_287),
.B2(n_249),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_315),
.Y(n_380)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_380),
.Y(n_411)
);

AO22x1_ASAP7_75t_SL g382 ( 
.A1(n_329),
.A2(n_193),
.B1(n_145),
.B2(n_131),
.Y(n_382)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

BUFx8_ASAP7_75t_L g383 ( 
.A(n_335),
.Y(n_383)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_331),
.B(n_312),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_387),
.Y(n_403)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_315),
.Y(n_385)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_385),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_310),
.A2(n_213),
.B(n_145),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_351),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_324),
.B(n_262),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_392),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_325),
.A2(n_244),
.B1(n_185),
.B2(n_182),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_391),
.A2(n_394),
.B1(n_297),
.B2(n_323),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_317),
.B(n_213),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_393),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_316),
.A2(n_131),
.B1(n_193),
.B2(n_230),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_323),
.B(n_230),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_398),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_313),
.B(n_293),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_396),
.A2(n_397),
.B(n_344),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_326),
.A2(n_293),
.B1(n_318),
.B2(n_341),
.Y(n_397)
);

AO22x1_ASAP7_75t_L g400 ( 
.A1(n_363),
.A2(n_329),
.B1(n_345),
.B2(n_326),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_400),
.A2(n_424),
.B(n_432),
.Y(n_454)
);

OAI22x1_ASAP7_75t_SL g405 ( 
.A1(n_374),
.A2(n_329),
.B1(n_341),
.B2(n_330),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_405),
.B(n_420),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_384),
.C(n_398),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_406),
.B(n_418),
.C(n_428),
.Y(n_441)
);

AOI22x1_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_329),
.B1(n_332),
.B2(n_297),
.Y(n_407)
);

OA22x2_ASAP7_75t_L g469 ( 
.A1(n_407),
.A2(n_417),
.B1(n_391),
.B2(n_382),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_412),
.A2(n_361),
.B1(n_390),
.B2(n_378),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_387),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_414),
.B(n_423),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_321),
.C(n_347),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_419),
.Y(n_449)
);

OAI32xp33_ASAP7_75t_L g420 ( 
.A1(n_370),
.A2(n_338),
.A3(n_343),
.B1(n_347),
.B2(n_333),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_377),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_362),
.A2(n_363),
.B(n_366),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_375),
.Y(n_426)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_426),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_368),
.B(n_366),
.C(n_354),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_369),
.A2(n_311),
.B1(n_295),
.B2(n_299),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_386),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_355),
.B(n_333),
.C(n_344),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_372),
.C(n_376),
.Y(n_443)
);

BUFx24_ASAP7_75t_SL g436 ( 
.A(n_356),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_369),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_415),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_438),
.B(n_439),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_408),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_410),
.B(n_381),
.Y(n_440)
);

CKINVDCx14_ASAP7_75t_R g498 ( 
.A(n_440),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_442),
.A2(n_407),
.B1(n_400),
.B2(n_432),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_443),
.B(n_460),
.Y(n_478)
);

INVx13_ASAP7_75t_L g444 ( 
.A(n_431),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_415),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_445),
.B(n_456),
.Y(n_505)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_447),
.Y(n_500)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_437),
.Y(n_448)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

A2O1A1O1Ixp25_ASAP7_75t_L g450 ( 
.A1(n_424),
.A2(n_355),
.B(n_357),
.C(n_353),
.D(n_389),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_450),
.A2(n_453),
.B(n_468),
.Y(n_491)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_402),
.Y(n_451)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_451),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_435),
.Y(n_452)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_452),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_409),
.Y(n_456)
);

INVx13_ASAP7_75t_L g457 ( 
.A(n_431),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_457),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_360),
.Y(n_458)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_429),
.B(n_353),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_461),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_413),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_380),
.Y(n_475)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_402),
.Y(n_463)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_463),
.Y(n_496)
);

NAND3xp33_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_466),
.C(n_470),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_403),
.B(n_421),
.Y(n_465)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_465),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_411),
.B(n_358),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_403),
.B(n_365),
.Y(n_467)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_467),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_401),
.A2(n_396),
.B(n_392),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_472),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_428),
.B(n_388),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_421),
.B(n_393),
.Y(n_471)
);

AO21x1_ASAP7_75t_L g473 ( 
.A1(n_471),
.A2(n_399),
.B(n_401),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_399),
.A2(n_386),
.B1(n_382),
.B2(n_367),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_472),
.A2(n_405),
.B1(n_453),
.B2(n_446),
.Y(n_503)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_473),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_446),
.A2(n_422),
.B1(n_434),
.B2(n_417),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_474),
.A2(n_477),
.B1(n_453),
.B2(n_487),
.Y(n_516)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_475),
.Y(n_511)
);

OAI21xp33_ASAP7_75t_SL g476 ( 
.A1(n_449),
.A2(n_422),
.B(n_400),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_476),
.B(n_482),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_418),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_406),
.C(n_427),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_483),
.B(n_485),
.C(n_467),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_441),
.B(n_427),
.C(n_416),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_469),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_416),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_490),
.B(n_497),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_456),
.B(n_439),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_492),
.B(n_493),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_466),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_407),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_460),
.B(n_385),
.Y(n_502)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_502),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_503),
.A2(n_469),
.B1(n_458),
.B2(n_455),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_459),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_504),
.B(n_447),
.Y(n_536)
);

AO22x1_ASAP7_75t_L g506 ( 
.A1(n_454),
.A2(n_433),
.B1(n_419),
.B2(n_420),
.Y(n_506)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_506),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_498),
.A2(n_459),
.B1(n_442),
.B2(n_464),
.Y(n_507)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_507),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_445),
.Y(n_509)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_509),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_479),
.B(n_455),
.Y(n_510)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_510),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_503),
.A2(n_438),
.B1(n_452),
.B2(n_471),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_512),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_513),
.B(n_518),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_505),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_515),
.B(n_536),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_516),
.A2(n_521),
.B1(n_525),
.B2(n_506),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_491),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_517),
.B(n_531),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_483),
.B(n_468),
.Y(n_518)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_520),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_487),
.A2(n_469),
.B1(n_443),
.B2(n_454),
.Y(n_521)
);

XNOR2x1_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_497),
.Y(n_543)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_505),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_524),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_474),
.A2(n_469),
.B1(n_412),
.B2(n_450),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_485),
.B(n_450),
.C(n_451),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_527),
.B(n_491),
.C(n_499),
.Y(n_538)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_481),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_528),
.B(n_529),
.Y(n_554)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_481),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_488),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_530),
.Y(n_555)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_488),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_478),
.B(n_463),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_534),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_489),
.B(n_462),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_533),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_490),
.B(n_448),
.Y(n_534)
);

MAJx2_ASAP7_75t_L g574 ( 
.A(n_538),
.B(n_359),
.C(n_457),
.Y(n_574)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_543),
.Y(n_568)
);

AOI21xp33_ASAP7_75t_L g544 ( 
.A1(n_523),
.A2(n_484),
.B(n_489),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_544),
.B(n_550),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_513),
.B(n_518),
.C(n_527),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_547),
.B(n_549),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_532),
.B(n_473),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_557),
.C(n_558),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_526),
.B(n_499),
.C(n_501),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_535),
.B(n_494),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_551),
.A2(n_522),
.B1(n_520),
.B2(n_509),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_511),
.A2(n_508),
.B1(n_514),
.B2(n_525),
.Y(n_556)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_556),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_526),
.B(n_501),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_517),
.C(n_521),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_519),
.A2(n_494),
.B1(n_480),
.B2(n_496),
.Y(n_561)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_561),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_552),
.A2(n_520),
.B1(n_533),
.B2(n_510),
.Y(n_564)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_564),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_552),
.A2(n_506),
.B1(n_516),
.B2(n_486),
.Y(n_565)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_565),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_553),
.B(n_496),
.Y(n_566)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_566),
.Y(n_594)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_554),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_569),
.A2(n_571),
.B1(n_577),
.B2(n_578),
.Y(n_592)
);

INVx13_ASAP7_75t_L g570 ( 
.A(n_540),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_570),
.B(n_575),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_546),
.A2(n_500),
.B1(n_486),
.B2(n_495),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_560),
.A2(n_495),
.B(n_457),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_572),
.A2(n_542),
.B(n_559),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_574),
.B(n_397),
.Y(n_598)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_545),
.Y(n_575)
);

BUFx12_ASAP7_75t_L g576 ( 
.A(n_543),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_576),
.A2(n_579),
.B(n_539),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_541),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_555),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_541),
.B(n_461),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_559),
.A2(n_382),
.B1(n_404),
.B2(n_394),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_581),
.A2(n_430),
.B1(n_404),
.B2(n_444),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_580),
.A2(n_547),
.B(n_538),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_583),
.A2(n_585),
.B(n_596),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_563),
.B(n_539),
.C(n_558),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_563),
.B(n_537),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_586),
.B(n_588),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_565),
.B(n_537),
.Y(n_588)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_589),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_567),
.A2(n_551),
.B1(n_542),
.B2(n_548),
.Y(n_590)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_590),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_573),
.A2(n_549),
.B1(n_557),
.B2(n_379),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_597),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_SL g610 ( 
.A(n_598),
.B(n_592),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_574),
.B(n_359),
.C(n_444),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_599),
.B(n_579),
.C(n_572),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_568),
.B(n_395),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_600),
.B(n_581),
.Y(n_611)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_601),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_585),
.B(n_562),
.C(n_564),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_608),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_593),
.A2(n_577),
.B1(n_582),
.B2(n_566),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_606),
.A2(n_589),
.B1(n_599),
.B2(n_588),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_568),
.C(n_576),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_610),
.B(n_614),
.Y(n_619)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_611),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_595),
.B(n_569),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_612),
.B(n_364),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_594),
.B(n_590),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_613),
.B(n_601),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_593),
.A2(n_576),
.B1(n_570),
.B2(n_311),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_606),
.A2(n_587),
.B1(n_584),
.B2(n_591),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_616),
.B(n_617),
.Y(n_633)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_618),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_602),
.B(n_600),
.Y(n_620)
);

NOR3xp33_ASAP7_75t_L g629 ( 
.A(n_620),
.B(n_609),
.C(n_610),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_621),
.B(n_371),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_604),
.B(n_364),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_622),
.B(n_625),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_607),
.B(n_598),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_615),
.B(n_605),
.C(n_603),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_627),
.B(n_629),
.Y(n_635)
);

NOR2x1_ASAP7_75t_SL g628 ( 
.A(n_616),
.B(n_608),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_628),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_623),
.B(n_614),
.C(n_339),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_630),
.B(n_631),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_633),
.A2(n_619),
.B(n_624),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_634),
.B(n_636),
.C(n_371),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_626),
.A2(n_620),
.B(n_619),
.Y(n_636)
);

AOI322xp5_ASAP7_75t_L g639 ( 
.A1(n_638),
.A2(n_632),
.A3(n_629),
.B1(n_630),
.B2(n_299),
.C1(n_295),
.C2(n_340),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_639),
.B(n_640),
.C(n_635),
.Y(n_641)
);

OAI211xp5_ASAP7_75t_L g642 ( 
.A1(n_641),
.A2(n_637),
.B(n_373),
.C(n_294),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_373),
.C(n_383),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_643),
.A2(n_294),
.B1(n_383),
.B2(n_638),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_383),
.B(n_294),
.Y(n_645)
);


endmodule