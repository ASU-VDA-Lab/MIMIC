module fake_jpeg_10913_n_575 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_575);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_575;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_8),
.B(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_57),
.Y(n_153)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_59),
.Y(n_157)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g127 ( 
.A(n_64),
.Y(n_127)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_7),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_68),
.B(n_71),
.Y(n_166)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_75),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_7),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_72),
.Y(n_131)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_73),
.Y(n_178)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_81),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_90),
.Y(n_181)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_35),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g150 ( 
.A(n_92),
.Y(n_150)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_31),
.B(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_106),
.Y(n_126)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_55),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_22),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_31),
.B(n_6),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_32),
.B(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_109),
.B(n_44),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_116),
.B(n_124),
.Y(n_210)
);

NAND2x1_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_22),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_118),
.A2(n_136),
.B(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_81),
.B(n_42),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_130),
.B(n_134),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_75),
.A2(n_33),
.B(n_52),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_56),
.A2(n_55),
.B1(n_33),
.B2(n_23),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_137),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_64),
.A2(n_33),
.B(n_82),
.Y(n_140)
);

NAND2xp67_ASAP7_75t_SL g211 ( 
.A(n_140),
.B(n_47),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_73),
.A2(n_55),
.B1(n_51),
.B2(n_50),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_52),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_143),
.B(n_155),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_90),
.B(n_32),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_84),
.A2(n_44),
.B1(n_40),
.B2(n_42),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_18),
.B1(n_34),
.B2(n_29),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_179),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_90),
.B(n_40),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_165),
.B(n_172),
.Y(n_244)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_108),
.B(n_51),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_170),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_72),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_74),
.Y(n_176)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_96),
.A2(n_51),
.B1(n_50),
.B2(n_49),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_25),
.B1(n_18),
.B2(n_28),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_78),
.B(n_30),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_30),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_99),
.Y(n_237)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_186),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_189),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_190),
.Y(n_299)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_191),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_118),
.A2(n_67),
.B1(n_57),
.B2(n_59),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g281 ( 
.A1(n_192),
.A2(n_203),
.B1(n_172),
.B2(n_131),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_193),
.B(n_222),
.Y(n_291)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_197),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_126),
.B(n_85),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_198),
.B(n_237),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_127),
.A2(n_66),
.B1(n_61),
.B2(n_79),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_199),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_202),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_140),
.A2(n_87),
.B1(n_104),
.B2(n_102),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_112),
.Y(n_208)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_208),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_110),
.B1(n_100),
.B2(n_86),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_209),
.A2(n_216),
.B1(n_224),
.B2(n_238),
.Y(n_296)
);

NOR2x1p5_ASAP7_75t_L g287 ( 
.A(n_211),
.B(n_225),
.Y(n_287)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

INVx4_ASAP7_75t_SL g297 ( 
.A(n_212),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_129),
.Y(n_214)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_141),
.A2(n_83),
.B1(n_25),
.B2(n_28),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_215),
.A2(n_182),
.B1(n_138),
.B2(n_178),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_132),
.A2(n_29),
.B1(n_34),
.B2(n_49),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_117),
.Y(n_218)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_121),
.Y(n_219)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

INVx3_ASAP7_75t_SL g302 ( 
.A(n_220),
.Y(n_302)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_113),
.Y(n_221)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_154),
.B(n_99),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_223),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_137),
.A2(n_36),
.B1(n_50),
.B2(n_49),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_SL g225 ( 
.A(n_169),
.B(n_48),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_151),
.A2(n_41),
.B1(n_24),
.B2(n_36),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_123),
.Y(n_227)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_227),
.Y(n_305)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_139),
.Y(n_228)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_228),
.Y(n_309)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_230),
.Y(n_264)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_112),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_231),
.Y(n_266)
);

INVx6_ASAP7_75t_SL g232 ( 
.A(n_150),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_232),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_145),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_234),
.Y(n_273)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_153),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_235),
.A2(n_236),
.B1(n_160),
.B2(n_164),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_153),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_144),
.A2(n_41),
.B1(n_36),
.B2(n_24),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_128),
.B(n_41),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_240),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_133),
.B(n_48),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_243),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_147),
.B(n_48),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_242),
.B(n_247),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_150),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_246),
.Y(n_280)
);

INVx11_ASAP7_75t_L g245 ( 
.A(n_131),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_135),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_149),
.B(n_46),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_145),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_182),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_249),
.B(n_250),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_156),
.B(n_46),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_188),
.B(n_225),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_251),
.B(n_253),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_184),
.B(n_146),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_211),
.A2(n_151),
.B1(n_142),
.B2(n_157),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_254),
.A2(n_279),
.B1(n_285),
.B2(n_298),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_204),
.B(n_114),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_263),
.B(n_265),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_204),
.B(n_114),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_204),
.B(n_195),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_269),
.B(n_270),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_185),
.B(n_120),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_185),
.A2(n_120),
.B1(n_146),
.B2(n_175),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_281),
.A2(n_207),
.B(n_202),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_217),
.B(n_175),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_284),
.B(n_288),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_210),
.B(n_178),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_290),
.B(n_301),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_243),
.B(n_130),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_292),
.B(n_303),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_197),
.A2(n_203),
.B1(n_192),
.B2(n_215),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_218),
.B(n_164),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_243),
.B(n_46),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_203),
.A2(n_157),
.B1(n_160),
.B2(n_47),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_222),
.B1(n_223),
.B2(n_236),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_307),
.A2(n_302),
.B1(n_261),
.B2(n_265),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_192),
.B(n_0),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_308),
.B(n_281),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_222),
.B(n_21),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_200),
.C(n_21),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_299),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_311),
.B(n_332),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_192),
.Y(n_313)
);

XNOR2x1_ASAP7_75t_SL g398 ( 
.A(n_313),
.B(n_297),
.Y(n_398)
);

NAND3xp33_ASAP7_75t_L g314 ( 
.A(n_259),
.B(n_232),
.C(n_212),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_314),
.B(n_350),
.Y(n_386)
);

AO22x1_ASAP7_75t_SL g316 ( 
.A1(n_298),
.A2(n_203),
.B1(n_245),
.B2(n_191),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_343),
.Y(n_365)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_284),
.Y(n_317)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_317),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_283),
.A2(n_293),
.B1(n_272),
.B2(n_279),
.Y(n_318)
);

OAI22x1_ASAP7_75t_L g383 ( 
.A1(n_318),
.A2(n_302),
.B1(n_258),
.B2(n_255),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_319),
.A2(n_321),
.B1(n_325),
.B2(n_348),
.Y(n_364)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_272),
.A2(n_241),
.B1(n_231),
.B2(n_234),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_320),
.A2(n_355),
.B1(n_268),
.B2(n_262),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_308),
.A2(n_205),
.B1(n_201),
.B2(n_206),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_322),
.Y(n_374)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_323),
.Y(n_367)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_296),
.A2(n_235),
.B1(n_220),
.B2(n_194),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_253),
.A2(n_208),
.B1(n_246),
.B2(n_213),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_329),
.A2(n_336),
.B1(n_337),
.B2(n_351),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_330),
.B(n_334),
.Y(n_381)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_331),
.Y(n_396)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_275),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_275),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_335),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_281),
.A2(n_196),
.B1(n_186),
.B2(n_214),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_339),
.B(n_310),
.Y(n_366)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_340),
.B(n_342),
.Y(n_377)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_276),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_256),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_260),
.B(n_8),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_344),
.B(n_347),
.Y(n_361)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_256),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_356),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_346),
.B(n_353),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_280),
.B(n_8),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_291),
.A2(n_21),
.B1(n_9),
.B2(n_11),
.Y(n_348)
);

MAJx2_ASAP7_75t_L g349 ( 
.A(n_269),
.B(n_6),
.C(n_15),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_255),
.C(n_268),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_264),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_293),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_282),
.B(n_6),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_283),
.A2(n_9),
.B(n_14),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_354),
.A2(n_287),
.B(n_291),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_263),
.A2(n_294),
.B1(n_290),
.B2(n_251),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_357),
.B(n_359),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_282),
.B(n_12),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_286),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_309),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_358),
.A2(n_287),
.B(n_291),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_362),
.A2(n_369),
.B(n_370),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_366),
.B(n_390),
.Y(n_415)
);

INVx5_ASAP7_75t_SL g368 ( 
.A(n_330),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_368),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_358),
.A2(n_287),
.B(n_252),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_312),
.A2(n_322),
.B1(n_317),
.B2(n_319),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_371),
.A2(n_384),
.B1(n_389),
.B2(n_336),
.Y(n_403)
);

A2O1A1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_338),
.A2(n_309),
.B(n_305),
.C(n_285),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_373),
.B(n_379),
.Y(n_412)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_354),
.A2(n_305),
.B(n_266),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_376),
.A2(n_402),
.B(n_297),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_315),
.B(n_338),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_329),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_393),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_382),
.A2(n_383),
.B(n_398),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_312),
.A2(n_325),
.B1(n_316),
.B2(n_321),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_395),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_316),
.A2(n_289),
.B1(n_302),
.B2(n_268),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_339),
.B(n_300),
.C(n_258),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_341),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_300),
.C(n_257),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_352),
.B(n_289),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_397),
.B(n_271),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_355),
.B(n_326),
.C(n_313),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_399),
.B(n_350),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_313),
.A2(n_297),
.B(n_257),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_403),
.A2(n_409),
.B1(n_414),
.B2(n_426),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_392),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_365),
.A2(n_333),
.B1(n_356),
.B2(n_348),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_408),
.A2(n_418),
.B1(n_364),
.B2(n_380),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_371),
.A2(n_333),
.B1(n_351),
.B2(n_311),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_410),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_393),
.B(n_360),
.Y(n_411)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_368),
.A2(n_349),
.B(n_328),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_413),
.A2(n_424),
.B(n_428),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_384),
.A2(n_357),
.B1(n_342),
.B2(n_340),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_379),
.B(n_331),
.Y(n_416)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_365),
.A2(n_327),
.B1(n_335),
.B2(n_334),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_375),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_422),
.Y(n_438)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_377),
.Y(n_421)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_421),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_381),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_372),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_433),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_385),
.B(n_324),
.Y(n_425)
);

OAI21xp33_ASAP7_75t_L g457 ( 
.A1(n_425),
.A2(n_401),
.B(n_387),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_392),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_372),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_427),
.B(n_430),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_368),
.A2(n_323),
.B(n_332),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_381),
.A2(n_345),
.B(n_343),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_386),
.B(n_267),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_431),
.A2(n_434),
.B1(n_382),
.B2(n_376),
.Y(n_445)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_389),
.A2(n_306),
.B1(n_267),
.B2(n_271),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_400),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_435),
.B(n_436),
.Y(n_466)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_396),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_1),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_415),
.B(n_399),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_L g478 ( 
.A(n_440),
.B(n_413),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_442),
.A2(n_449),
.B1(n_453),
.B2(n_409),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_366),
.C(n_390),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_447),
.C(n_448),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_445),
.A2(n_446),
.B1(n_461),
.B2(n_463),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_403),
.A2(n_391),
.B1(n_374),
.B2(n_363),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_362),
.C(n_395),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_404),
.B(n_370),
.C(n_398),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_408),
.A2(n_381),
.B1(n_364),
.B2(n_363),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_406),
.B(n_388),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_450),
.B(n_413),
.Y(n_487)
);

OAI32xp33_ASAP7_75t_L g452 ( 
.A1(n_412),
.A2(n_374),
.A3(n_373),
.B1(n_397),
.B2(n_385),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_452),
.B(n_421),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_422),
.A2(n_394),
.B1(n_369),
.B2(n_383),
.Y(n_453)
);

FAx1_ASAP7_75t_SL g454 ( 
.A(n_412),
.B(n_394),
.CI(n_402),
.CON(n_454),
.SN(n_454)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_467),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_411),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_457),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_406),
.B(n_400),
.C(n_378),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_459),
.C(n_464),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_407),
.B(n_391),
.C(n_387),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_414),
.A2(n_361),
.B1(n_367),
.B2(n_4),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_405),
.A2(n_361),
.B1(n_367),
.B2(n_4),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_1),
.C(n_3),
.Y(n_464)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_468),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_451),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_442),
.A2(n_405),
.B1(n_420),
.B2(n_427),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_472),
.A2(n_481),
.B1(n_488),
.B2(n_489),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_475),
.A2(n_493),
.B1(n_425),
.B2(n_454),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_465),
.A2(n_417),
.B(n_419),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_476),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_477),
.A2(n_483),
.B1(n_492),
.B2(n_446),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_478),
.B(n_487),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_440),
.C(n_447),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_479),
.B(n_491),
.C(n_494),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_431),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_480),
.B(n_484),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_456),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_466),
.Y(n_482)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_482),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_449),
.A2(n_453),
.B1(n_459),
.B2(n_438),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_443),
.B(n_416),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_466),
.Y(n_485)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_485),
.Y(n_515)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_460),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_465),
.A2(n_438),
.B(n_417),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_490),
.B(n_428),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_450),
.B(n_410),
.C(n_435),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_451),
.A2(n_423),
.B1(n_424),
.B2(n_433),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_460),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_448),
.B(n_430),
.C(n_419),
.Y(n_494)
);

AND2x2_ASAP7_75t_SL g519 ( 
.A(n_495),
.B(n_483),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_496),
.A2(n_497),
.B1(n_511),
.B2(n_486),
.Y(n_518)
);

NOR2x1_ASAP7_75t_SL g497 ( 
.A(n_491),
.B(n_458),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_498),
.B(n_509),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_441),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_500),
.B(n_502),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_470),
.B(n_479),
.C(n_474),
.Y(n_502)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_503),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g505 ( 
.A(n_471),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_505),
.B(n_513),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_474),
.B(n_439),
.C(n_462),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_507),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_463),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_452),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_477),
.A2(n_454),
.B1(n_461),
.B2(n_462),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_486),
.A2(n_468),
.B1(n_464),
.B2(n_437),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_478),
.B(n_418),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_516),
.C(n_476),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_469),
.B(n_432),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_518),
.A2(n_515),
.B1(n_510),
.B2(n_15),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_524),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_495),
.B(n_490),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_526),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_501),
.A2(n_489),
.B(n_471),
.Y(n_521)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_521),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_508),
.A2(n_493),
.B(n_488),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_523),
.A2(n_527),
.B(n_510),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g526 ( 
.A(n_512),
.Y(n_526)
);

AO21x1_ASAP7_75t_L g527 ( 
.A1(n_508),
.A2(n_472),
.B(n_492),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_502),
.B(n_485),
.C(n_482),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_528),
.B(n_531),
.C(n_533),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_473),
.C(n_436),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_499),
.A2(n_473),
.B1(n_12),
.B2(n_14),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_504),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_501),
.B(n_3),
.C(n_5),
.Y(n_533)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_522),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_535),
.B(n_536),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_520),
.A2(n_496),
.B(n_511),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_523),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_528),
.B(n_509),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_539),
.B(n_540),
.Y(n_550)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_525),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_531),
.B(n_498),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_541),
.B(n_547),
.Y(n_556)
);

AOI21xp33_ASAP7_75t_L g543 ( 
.A1(n_529),
.A2(n_520),
.B(n_530),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_543),
.A2(n_527),
.B(n_532),
.Y(n_553)
);

XNOR2x1_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_533),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_546),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_517),
.B(n_5),
.C(n_14),
.Y(n_547)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_548),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_544),
.B(n_524),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_552),
.B(n_547),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_553),
.A2(n_555),
.B(n_557),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_SL g561 ( 
.A(n_554),
.B(n_534),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_544),
.B(n_517),
.C(n_519),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_542),
.B(n_519),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_550),
.A2(n_538),
.B(n_542),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_558),
.B(n_559),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_555),
.A2(n_546),
.B(n_537),
.Y(n_559)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_561),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_534),
.C(n_545),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_562),
.B(n_563),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_560),
.B(n_556),
.Y(n_568)
);

INVxp33_ASAP7_75t_L g569 ( 
.A(n_568),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_566),
.A2(n_564),
.B(n_548),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_567),
.B(n_565),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_571),
.A2(n_569),
.B(n_557),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_561),
.B(n_551),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_554),
.B(n_5),
.Y(n_574)
);

BUFx24_ASAP7_75t_SL g575 ( 
.A(n_574),
.Y(n_575)
);


endmodule