module fake_jpeg_2682_n_236 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_236);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_235;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_1),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_23),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_7),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_86),
.Y(n_95)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_84),
.Y(n_92)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_79),
.B1(n_77),
.B2(n_73),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_76),
.B1(n_55),
.B2(n_57),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_93),
.B1(n_100),
.B2(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_75),
.B1(n_57),
.B2(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_54),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_75),
.B1(n_67),
.B2(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_61),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_64),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_119),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_85),
.B1(n_67),
.B2(n_73),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_107),
.A2(n_112),
.B1(n_120),
.B2(n_65),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_61),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_66),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

BUFx6f_ASAP7_75t_SL g136 ( 
.A(n_115),
.Y(n_136)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_122),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_79),
.C(n_64),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_82),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_54),
.B1(n_78),
.B2(n_68),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_62),
.B1(n_68),
.B2(n_60),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_88),
.B1(n_59),
.B2(n_72),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_53),
.B1(n_58),
.B2(n_98),
.Y(n_129)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_71),
.B(n_70),
.C(n_56),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_126),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_99),
.B1(n_96),
.B2(n_98),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_139),
.B1(n_131),
.B2(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_133),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_96),
.B(n_81),
.C(n_82),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_134),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_121),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_141),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_81),
.B1(n_101),
.B2(n_62),
.Y(n_137)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_101),
.B1(n_88),
.B2(n_98),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_0),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_1),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_107),
.B1(n_122),
.B2(n_65),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_148),
.B(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_169),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_116),
.C(n_117),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_161),
.C(n_28),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_167),
.B1(n_168),
.B2(n_137),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_81),
.B(n_65),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_29),
.B(n_42),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_65),
.B(n_3),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_123),
.B(n_129),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_51),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_49),
.B1(n_48),
.B2(n_47),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_187),
.B(n_157),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_SL g178 ( 
.A1(n_164),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_180),
.B(n_182),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_137),
.B1(n_10),
.B2(n_12),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_186),
.B1(n_34),
.B2(n_39),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_8),
.B1(n_14),
.B2(n_16),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_18),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_14),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_162),
.B(n_153),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_191),
.B(n_167),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_16),
.B(n_17),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_199),
.B1(n_205),
.B2(n_186),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_146),
.C(n_161),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_188),
.C(n_181),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_197),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

AOI221xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.C(n_20),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_33),
.B(n_40),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_202),
.B(n_177),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_31),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_46),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_215),
.C(n_36),
.Y(n_218)
);

OAI321xp33_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_183),
.A3(n_191),
.B1(n_182),
.B2(n_187),
.C(n_185),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_209),
.B1(n_212),
.B2(n_214),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_172),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_35),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_211),
.B(n_202),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_183),
.B1(n_184),
.B2(n_179),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_204),
.B1(n_196),
.B2(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_219),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_23),
.Y(n_220)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_21),
.B1(n_22),
.B2(n_206),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_219),
.Y(n_227)
);

NOR2xp67_ASAP7_75t_SL g231 ( 
.A(n_227),
.B(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_223),
.B(n_222),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_228),
.A2(n_229),
.B(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_233),
.A2(n_220),
.B(n_225),
.C(n_231),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_234),
.B(n_215),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_235),
.B(n_22),
.Y(n_236)
);


endmodule