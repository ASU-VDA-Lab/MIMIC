module fake_jpeg_22577_n_324 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_39),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_24),
.B1(n_27),
.B2(n_22),
.Y(n_65)
);

AO22x1_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_24),
.B1(n_28),
.B2(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_58),
.B1(n_36),
.B2(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_27),
.B1(n_19),
.B2(n_22),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_18),
.B1(n_29),
.B2(n_33),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_20),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_32),
.A2(n_27),
.B1(n_22),
.B2(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_62),
.Y(n_100)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_38),
.B1(n_36),
.B2(n_30),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_73),
.B1(n_75),
.B2(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_56),
.B1(n_53),
.B2(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_68),
.B(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_74),
.B1(n_77),
.B2(n_80),
.Y(n_96)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_23),
.B1(n_16),
.B2(n_30),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_42),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_16),
.B1(n_29),
.B2(n_18),
.Y(n_79)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_87),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_31),
.B(n_15),
.C(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_85),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_91),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_70),
.B1(n_51),
.B2(n_76),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_72),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_97),
.Y(n_121)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

OR2x4_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_57),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_100),
.B(n_63),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_69),
.A2(n_42),
.B1(n_56),
.B2(n_43),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_59),
.B1(n_62),
.B2(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_114),
.B1(n_116),
.B2(n_102),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_66),
.C(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_112),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_78),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_65),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_52),
.Y(n_144)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_74),
.B1(n_56),
.B2(n_80),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_52),
.B1(n_70),
.B2(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_105),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_123),
.B1(n_47),
.B2(n_49),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_125),
.B(n_84),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_83),
.A2(n_51),
.B1(n_76),
.B2(n_43),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_130),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_77),
.B(n_18),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_42),
.C(n_31),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_84),
.C(n_102),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_40),
.B(n_21),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_87),
.B1(n_94),
.B2(n_95),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_52),
.B1(n_76),
.B2(n_43),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_105),
.B1(n_89),
.B2(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_104),
.B1(n_89),
.B2(n_87),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_136),
.B1(n_137),
.B2(n_148),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_138),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_116),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_147),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_82),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_140),
.B(n_8),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_142),
.B(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_82),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_110),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_104),
.B1(n_91),
.B2(n_40),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_50),
.B(n_90),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_154),
.B(n_155),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_94),
.B1(n_87),
.B2(n_97),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_129),
.B1(n_111),
.B2(n_21),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_49),
.B(n_8),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_161),
.C(n_162),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_120),
.B(n_128),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_159),
.A2(n_170),
.B(n_5),
.Y(n_204)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_164),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_134),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_114),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_143),
.C(n_141),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_140),
.C(n_139),
.Y(n_184)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_109),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_5),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_169),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_145),
.B(n_154),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_126),
.C(n_125),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_126),
.B(n_106),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_149),
.B(n_138),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_150),
.B1(n_137),
.B2(n_148),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_183),
.B1(n_111),
.B2(n_7),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_178),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_7),
.Y(n_197)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_155),
.A2(n_111),
.B1(n_1),
.B2(n_0),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_200),
.C(n_205),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_185),
.A2(n_192),
.B1(n_198),
.B2(n_206),
.Y(n_231)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_209),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_153),
.B(n_152),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_193),
.A2(n_203),
.B1(n_168),
.B2(n_174),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_6),
.B(n_12),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_195),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_6),
.B(n_12),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_0),
.Y(n_196)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_204),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_180),
.A2(n_7),
.B1(n_12),
.B2(n_2),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_173),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_0),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_164),
.B1(n_157),
.B2(n_172),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_0),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_176),
.A2(n_7),
.B(n_2),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_189),
.B(n_165),
.Y(n_214)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_217),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_207),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_168),
.B1(n_172),
.B2(n_166),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_224),
.B1(n_228),
.B2(n_193),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_165),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_223),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_206),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_161),
.C(n_162),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_184),
.C(n_205),
.Y(n_242)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_178),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_229),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_183),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_191),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_232),
.B(n_219),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_187),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_242),
.C(n_244),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_177),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_239),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_231),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_248),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g238 ( 
.A(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_205),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_184),
.C(n_190),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_190),
.C(n_200),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_246),
.C(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_200),
.C(n_202),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_185),
.Y(n_249)
);

XOR2x2_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_204),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_215),
.B(n_195),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_245),
.B(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_231),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_266),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_254),
.A2(n_269),
.B(n_198),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_216),
.B1(n_215),
.B2(n_188),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_258),
.B1(n_211),
.B2(n_213),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_234),
.A2(n_186),
.B1(n_209),
.B2(n_211),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_213),
.Y(n_260)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_263),
.Y(n_270)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_219),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_268),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_220),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_237),
.B1(n_241),
.B2(n_186),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_246),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_191),
.B(n_194),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_233),
.C(n_240),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_274),
.C(n_276),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_247),
.C(n_229),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_260),
.B(n_261),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_197),
.C(n_1),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_266),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_267),
.B(n_9),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_4),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_1),
.C(n_3),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_284),
.C(n_4),
.Y(n_295)
);

INVx11_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_257),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_1),
.C(n_3),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_258),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_256),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_297),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_256),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_291),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_293),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_282),
.B1(n_283),
.B2(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_296),
.B1(n_272),
.B2(n_9),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_273),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_261),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_5),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_270),
.B(n_278),
.C(n_274),
.Y(n_300)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_SL g303 ( 
.A(n_285),
.B(n_278),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_285),
.B(n_293),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_306),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_302),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_310),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_296),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_311),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_287),
.C(n_295),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_314),
.B(n_300),
.C(n_299),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_315),
.B(n_313),
.Y(n_318)
);

O2A1O1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_315),
.B(n_317),
.C(n_316),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_305),
.A3(n_301),
.B1(n_308),
.B2(n_314),
.C1(n_312),
.C2(n_11),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_13),
.Y(n_321)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_13),
.B(n_10),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_13),
.C(n_10),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_10),
.B1(n_11),
.B2(n_321),
.Y(n_324)
);


endmodule