module fake_jpeg_30276_n_64 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_64);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_64;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_3),
.B(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_33),
.B1(n_29),
.B2(n_6),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_29),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_5),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_13),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_5),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_31),
.B(n_16),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_11),
.B(n_18),
.C(n_19),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_15),
.B1(n_21),
.B2(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_50),
.B1(n_7),
.B2(n_10),
.Y(n_56)
);

OA21x2_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_37),
.B(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_52),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_46),
.B(n_49),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_40),
.C(n_22),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_45),
.C(n_53),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_50),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_58),
.A2(n_59),
.B(n_60),
.Y(n_62)
);

AOI222xp33_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.C1(n_59),
.C2(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_62),
.Y(n_64)
);


endmodule