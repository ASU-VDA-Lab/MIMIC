module fake_aes_6357_n_21 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_21;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
NAND2xp5_ASAP7_75t_SL g8 ( .A(n_5), .B(n_1), .Y(n_8) );
INVx1_ASAP7_75t_SL g9 ( .A(n_2), .Y(n_9) );
BUFx10_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_2), .B(n_3), .Y(n_11) );
AND2x6_ASAP7_75t_L g12 ( .A(n_1), .B(n_6), .Y(n_12) );
OAI21xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_7), .B(n_3), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
OAI21x1_ASAP7_75t_SL g15 ( .A1(n_11), .A2(n_0), .B(n_4), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_14), .B(n_10), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_14), .B(n_10), .Y(n_17) );
OAI22xp5_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_13), .B1(n_14), .B2(n_9), .Y(n_18) );
NAND4xp25_ASAP7_75t_L g19 ( .A(n_18), .B(n_8), .C(n_16), .D(n_17), .Y(n_19) );
AOI22x1_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_15), .B1(n_12), .B2(n_6), .Y(n_20) );
AOI22xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_0), .B1(n_5), .B2(n_19), .Y(n_21) );
endmodule