module real_jpeg_16138_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_288;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_249;
wire n_215;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_0),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_0),
.Y(n_108)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_0),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_1),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_1),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_1),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_1),
.Y(n_228)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_2),
.Y(n_130)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_3),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_3),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_4),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_4),
.Y(n_136)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_5),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_6),
.A2(n_279),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_6),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g135 ( 
.A(n_8),
.Y(n_135)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_8),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_49),
.B1(n_55),
.B2(n_59),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_9),
.A2(n_49),
.B1(n_142),
.B2(n_144),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_9),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_9),
.B(n_91),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_9),
.B(n_226),
.C(n_229),
.Y(n_225)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_261),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_180),
.B(n_258),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_168),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_15),
.B(n_168),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_119),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_16),
.B(n_121),
.C(n_163),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_69),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_17),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_52),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_18),
.A2(n_52),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_18),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_26),
.B(n_36),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_24),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B(n_47),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_49),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_49),
.A2(n_113),
.B(n_115),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_49),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_49),
.B(n_148),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_49),
.B(n_244),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_52),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_52),
.A2(n_53),
.B1(n_178),
.B2(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_52),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_52),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_52),
.B(n_237),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g247 ( 
.A(n_52),
.B(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_64),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_54),
.A2(n_123),
.B1(n_131),
.B2(n_132),
.Y(n_122)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_58),
.A2(n_149),
.B1(n_151),
.B2(n_153),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_58),
.Y(n_229)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_62),
.Y(n_242)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_66),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_68),
.Y(n_246)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_70),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_70),
.Y(n_287)
);

XNOR2x1_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_90),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_71),
.B(n_90),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_71),
.B(n_140),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_71),
.B(n_90),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_85),
.Y(n_77)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_78),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_90),
.B(n_140),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_90),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_101),
.B(n_112),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_102),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B1(n_107),
.B2(n_109),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_115),
.A2(n_193),
.A3(n_195),
.B1(n_198),
.B2(n_204),
.Y(n_192)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_163),
.B2(n_164),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_139),
.B1(n_140),
.B2(n_162),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_122),
.B(n_140),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_123),
.A2(n_132),
.B1(n_274),
.B2(n_277),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_135),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_137),
.Y(n_284)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_140),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_139),
.A2(n_140),
.B1(n_190),
.B2(n_191),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_139),
.A2(n_166),
.B(n_172),
.C(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_139),
.A2(n_140),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_139),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_139),
.A2(n_140),
.B1(n_224),
.B2(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_139),
.B(n_175),
.C(n_222),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_139),
.A2(n_140),
.B1(n_273),
.B2(n_285),
.Y(n_272)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_155),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AND3x1_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.C(n_167),
.Y(n_164)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_165),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.C(n_177),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_171),
.A2(n_214),
.B1(n_215),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_171),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_175),
.C(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_172),
.A2(n_173),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_177),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_192),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AO21x2_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_209),
.B(n_257),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_183),
.B(n_185),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.C(n_208),
.Y(n_185)
);

XOR2x2_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

OAI21x1_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_216),
.B(n_256),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21x1_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_251),
.B(n_255),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_232),
.B(n_250),
.Y(n_217)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_223),
.Y(n_250)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2x1_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_247),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_290),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_266),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_286),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_288),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);


endmodule