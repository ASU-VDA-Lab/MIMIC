module real_aes_2308_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_335;
wire n_177;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_0), .B(n_151), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_1), .A2(n_133), .B(n_184), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_2), .A2(n_457), .B1(n_462), .B2(n_807), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_3), .B(n_821), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_4), .A2(n_11), .B1(n_118), .B2(n_119), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_4), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_5), .B(n_141), .Y(n_197) );
INVx1_ASAP7_75t_L g138 ( .A(n_6), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_7), .B(n_141), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_8), .A2(n_113), .B1(n_437), .B2(n_438), .Y(n_112) );
INVxp67_ASAP7_75t_L g438 ( .A(n_8), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_8), .B(n_128), .Y(n_498) );
INVx1_ASAP7_75t_L g526 ( .A(n_9), .Y(n_526) );
CKINVDCx16_ASAP7_75t_R g821 ( .A(n_10), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_11), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_12), .Y(n_541) );
NAND2xp33_ASAP7_75t_L g178 ( .A(n_13), .B(n_145), .Y(n_178) );
INVx2_ASAP7_75t_L g130 ( .A(n_14), .Y(n_130) );
AOI221x1_ASAP7_75t_L g220 ( .A1(n_15), .A2(n_28), .B1(n_133), .B2(n_151), .C(n_221), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g442 ( .A(n_16), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_17), .B(n_151), .Y(n_174) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_18), .A2(n_172), .B(n_173), .Y(n_171) );
INVx1_ASAP7_75t_L g507 ( .A(n_19), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_20), .B(n_164), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_21), .B(n_141), .Y(n_140) );
AO21x1_ASAP7_75t_L g192 ( .A1(n_22), .A2(n_151), .B(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g446 ( .A(n_23), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_24), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g505 ( .A(n_25), .Y(n_505) );
INVx1_ASAP7_75t_SL g491 ( .A(n_26), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_27), .B(n_152), .Y(n_585) );
NAND2x1_ASAP7_75t_L g206 ( .A(n_29), .B(n_141), .Y(n_206) );
AOI33xp33_ASAP7_75t_L g553 ( .A1(n_30), .A2(n_55), .A3(n_481), .B1(n_488), .B2(n_554), .B3(n_555), .Y(n_553) );
NAND2x1_ASAP7_75t_L g160 ( .A(n_31), .B(n_145), .Y(n_160) );
INVx1_ASAP7_75t_L g535 ( .A(n_32), .Y(n_535) );
OR2x2_ASAP7_75t_L g129 ( .A(n_33), .B(n_90), .Y(n_129) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_33), .A2(n_90), .B(n_130), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_34), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_35), .B(n_145), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_36), .B(n_141), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_37), .B(n_145), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_38), .A2(n_133), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g134 ( .A(n_39), .B(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g149 ( .A(n_39), .B(n_138), .Y(n_149) );
INVx1_ASAP7_75t_L g487 ( .A(n_39), .Y(n_487) );
OR2x6_ASAP7_75t_L g444 ( .A(n_40), .B(n_445), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g819 ( .A(n_40), .B(n_820), .C(n_822), .Y(n_819) );
XNOR2xp5_ASAP7_75t_L g458 ( .A(n_41), .B(n_459), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_42), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_43), .B(n_151), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_44), .B(n_479), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_45), .A2(n_128), .B1(n_168), .B2(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_46), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_47), .B(n_152), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_48), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_49), .B(n_145), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_50), .B(n_172), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_51), .B(n_152), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_52), .A2(n_133), .B(n_159), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_53), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_54), .B(n_145), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_56), .B(n_152), .Y(n_565) );
INVx1_ASAP7_75t_L g137 ( .A(n_57), .Y(n_137) );
INVx1_ASAP7_75t_L g147 ( .A(n_57), .Y(n_147) );
AND2x2_ASAP7_75t_L g566 ( .A(n_58), .B(n_164), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g524 ( .A1(n_59), .A2(n_77), .B1(n_479), .B2(n_485), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_60), .B(n_479), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_61), .B(n_141), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_62), .B(n_168), .Y(n_543) );
AOI21xp5_ASAP7_75t_SL g515 ( .A1(n_63), .A2(n_485), .B(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_64), .A2(n_133), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g501 ( .A(n_65), .Y(n_501) );
AO21x1_ASAP7_75t_L g194 ( .A1(n_66), .A2(n_133), .B(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_67), .B(n_151), .Y(n_182) );
INVxp33_ASAP7_75t_L g824 ( .A(n_68), .Y(n_824) );
INVx1_ASAP7_75t_L g564 ( .A(n_69), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_70), .B(n_151), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_71), .A2(n_485), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g243 ( .A(n_72), .B(n_165), .Y(n_243) );
INVx1_ASAP7_75t_L g135 ( .A(n_73), .Y(n_135) );
INVx1_ASAP7_75t_L g143 ( .A(n_73), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_74), .A2(n_100), .B1(n_460), .B2(n_461), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_74), .Y(n_460) );
AND2x2_ASAP7_75t_L g166 ( .A(n_75), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_76), .B(n_479), .Y(n_556) );
AND2x2_ASAP7_75t_L g494 ( .A(n_78), .B(n_167), .Y(n_494) );
INVx1_ASAP7_75t_L g502 ( .A(n_79), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_80), .A2(n_485), .B(n_490), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g583 ( .A1(n_81), .A2(n_485), .B(n_548), .C(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g447 ( .A(n_82), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_83), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g180 ( .A(n_84), .B(n_167), .Y(n_180) );
AND2x2_ASAP7_75t_SL g513 ( .A(n_85), .B(n_167), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_86), .A2(n_485), .B1(n_551), .B2(n_552), .Y(n_550) );
OAI22xp5_ASAP7_75t_SL g114 ( .A1(n_87), .A2(n_115), .B1(n_116), .B2(n_117), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_87), .Y(n_115) );
XNOR2xp5_ASAP7_75t_L g457 ( .A(n_88), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g193 ( .A(n_89), .B(n_128), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_91), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g210 ( .A(n_92), .B(n_167), .Y(n_210) );
INVx1_ASAP7_75t_L g517 ( .A(n_93), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_94), .B(n_141), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_95), .A2(n_133), .B(n_139), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_96), .B(n_145), .Y(n_222) );
AND2x2_ASAP7_75t_L g557 ( .A(n_97), .B(n_167), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_98), .B(n_141), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_99), .A2(n_533), .B(n_534), .C(n_536), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_100), .Y(n_461) );
BUFx2_ASAP7_75t_L g110 ( .A(n_101), .Y(n_110) );
BUFx2_ASAP7_75t_SL g454 ( .A(n_101), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_102), .A2(n_133), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_103), .B(n_152), .Y(n_518) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_815), .B(n_823), .Y(n_104) );
OA22x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B1(n_451), .B2(n_455), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_439), .B(n_448), .Y(n_111) );
INVx1_ASAP7_75t_L g437 ( .A(n_113), .Y(n_437) );
XNOR2x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_120), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_120), .A2(n_463), .B1(n_467), .B2(n_470), .Y(n_462) );
INVx2_ASAP7_75t_L g812 ( .A(n_120), .Y(n_812) );
OR2x6_ASAP7_75t_L g120 ( .A(n_121), .B(n_335), .Y(n_120) );
NAND3xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_247), .C(n_302), .Y(n_121) );
AOI221xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_187), .B1(n_211), .B2(n_215), .C(n_225), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_170), .Y(n_123) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_124), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g246 ( .A(n_124), .Y(n_246) );
AND2x2_ASAP7_75t_L g291 ( .A(n_124), .B(n_228), .Y(n_291) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_155), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g279 ( .A(n_126), .Y(n_279) );
INVx1_ASAP7_75t_L g289 ( .A(n_126), .Y(n_289) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_131), .B(n_153), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_127), .B(n_154), .Y(n_153) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_127), .A2(n_131), .B(n_153), .Y(n_253) );
INVx1_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_128), .A2(n_174), .B(n_175), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_128), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_128), .B(n_148), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_128), .A2(n_515), .B(n_519), .Y(n_514) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_129), .B(n_130), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_150), .Y(n_131) );
AND2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
BUFx3_ASAP7_75t_L g483 ( .A(n_134), .Y(n_483) );
AND2x6_ASAP7_75t_L g145 ( .A(n_135), .B(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g489 ( .A(n_135), .Y(n_489) );
AND2x4_ASAP7_75t_L g485 ( .A(n_136), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x4_ASAP7_75t_L g141 ( .A(n_137), .B(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g481 ( .A(n_137), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_138), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_144), .B(n_148), .Y(n_139) );
INVxp67_ASAP7_75t_L g508 ( .A(n_141), .Y(n_508) );
AND2x4_ASAP7_75t_L g152 ( .A(n_142), .B(n_146), .Y(n_152) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVxp67_ASAP7_75t_L g506 ( .A(n_145), .Y(n_506) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_148), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_148), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_148), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_148), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_148), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_148), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_148), .A2(n_240), .B(n_241), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_148), .A2(n_491), .B(n_492), .C(n_493), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_148), .A2(n_492), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_SL g525 ( .A1(n_148), .A2(n_492), .B(n_526), .C(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g551 ( .A(n_148), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_148), .A2(n_492), .B(n_564), .C(n_565), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_148), .A2(n_585), .B(n_586), .Y(n_584) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g151 ( .A(n_149), .B(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_149), .Y(n_536) );
INVx1_ASAP7_75t_L g503 ( .A(n_152), .Y(n_503) );
OR2x2_ASAP7_75t_L g268 ( .A(n_155), .B(n_171), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_155), .B(n_214), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_155), .B(n_179), .Y(n_312) );
INVx2_ASAP7_75t_L g321 ( .A(n_155), .Y(n_321) );
AND2x2_ASAP7_75t_L g342 ( .A(n_155), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g426 ( .A(n_155), .B(n_245), .Y(n_426) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g254 ( .A(n_156), .B(n_179), .Y(n_254) );
AND2x2_ASAP7_75t_L g387 ( .A(n_156), .B(n_214), .Y(n_387) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_156), .Y(n_413) );
AO21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_163), .B(n_166), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_162), .Y(n_157) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_163), .A2(n_477), .B(n_494), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_164), .A2(n_182), .B(n_183), .Y(n_181) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_164), .A2(n_220), .B(n_224), .Y(n_219) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_164), .A2(n_220), .B(n_224), .Y(n_231) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g209 ( .A(n_167), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_167), .A2(n_209), .B1(n_532), .B2(n_537), .Y(n_531) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_168), .B(n_540), .Y(n_539) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_169), .Y(n_172) );
AND2x4_ASAP7_75t_L g341 ( .A(n_170), .B(n_342), .Y(n_341) );
AOI321xp33_ASAP7_75t_L g355 ( .A1(n_170), .A2(n_284), .A3(n_285), .B1(n_317), .B2(n_356), .C(n_359), .Y(n_355) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_179), .Y(n_170) );
BUFx3_ASAP7_75t_L g212 ( .A(n_171), .Y(n_212) );
INVx2_ASAP7_75t_L g245 ( .A(n_171), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_171), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g278 ( .A(n_171), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g311 ( .A(n_171), .Y(n_311) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_172), .A2(n_524), .B(n_528), .Y(n_523) );
INVx2_ASAP7_75t_SL g548 ( .A(n_172), .Y(n_548) );
INVx5_ASAP7_75t_L g214 ( .A(n_179), .Y(n_214) );
NOR2x1_ASAP7_75t_SL g263 ( .A(n_179), .B(n_253), .Y(n_263) );
BUFx2_ASAP7_75t_L g358 ( .A(n_179), .Y(n_358) );
OR2x6_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVxp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_200), .Y(n_188) );
NOR2xp33_ASAP7_75t_SL g256 ( .A(n_189), .B(n_257), .Y(n_256) );
NOR4xp25_ASAP7_75t_L g359 ( .A(n_189), .B(n_353), .C(n_357), .D(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g397 ( .A(n_189), .Y(n_397) );
AND2x2_ASAP7_75t_L g431 ( .A(n_189), .B(n_371), .Y(n_431) );
BUFx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g232 ( .A(n_190), .Y(n_232) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g286 ( .A(n_191), .Y(n_286) );
OAI21x1_ASAP7_75t_SL g191 ( .A1(n_192), .A2(n_194), .B(n_198), .Y(n_191) );
INVx1_ASAP7_75t_L g199 ( .A(n_193), .Y(n_199) );
AOI33xp33_ASAP7_75t_L g427 ( .A1(n_200), .A2(n_229), .A3(n_260), .B1(n_276), .B2(n_382), .B3(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g217 ( .A(n_201), .B(n_218), .Y(n_217) );
AND2x4_ASAP7_75t_L g227 ( .A(n_201), .B(n_228), .Y(n_227) );
BUFx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g234 ( .A(n_202), .Y(n_234) );
INVxp67_ASAP7_75t_L g315 ( .A(n_202), .Y(n_315) );
AND2x2_ASAP7_75t_L g371 ( .A(n_202), .B(n_236), .Y(n_371) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_209), .B(n_210), .Y(n_202) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_203), .A2(n_209), .B(n_210), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_208), .Y(n_203) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_209), .A2(n_237), .B(n_243), .Y(n_236) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_209), .A2(n_237), .B(n_243), .Y(n_272) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_209), .A2(n_560), .B(n_566), .Y(n_559) );
AO21x2_ASAP7_75t_L g597 ( .A1(n_209), .A2(n_560), .B(n_566), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_211), .A2(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AND2x2_ASAP7_75t_L g380 ( .A(n_212), .B(n_254), .Y(n_380) );
AND3x2_ASAP7_75t_L g382 ( .A(n_212), .B(n_266), .C(n_321), .Y(n_382) );
INVx3_ASAP7_75t_SL g334 ( .A(n_213), .Y(n_334) );
INVx4_ASAP7_75t_L g228 ( .A(n_214), .Y(n_228) );
AND2x2_ASAP7_75t_L g266 ( .A(n_214), .B(n_253), .Y(n_266) );
INVxp67_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g260 ( .A(n_218), .Y(n_260) );
AND2x4_ASAP7_75t_L g285 ( .A(n_218), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g348 ( .A(n_218), .B(n_236), .Y(n_348) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g318 ( .A(n_219), .Y(n_318) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_219), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_R g225 ( .A1(n_226), .A2(n_229), .B(n_233), .C(n_244), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g277 ( .A(n_228), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_228), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_228), .B(n_245), .Y(n_406) );
INVx1_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g388 ( .A(n_230), .B(n_378), .Y(n_388) );
AND2x2_ASAP7_75t_SL g230 ( .A(n_231), .B(n_232), .Y(n_230) );
AND2x2_ASAP7_75t_L g235 ( .A(n_231), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g257 ( .A(n_231), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g273 ( .A(n_231), .B(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g306 ( .A(n_231), .B(n_286), .Y(n_306) );
AND2x4_ASAP7_75t_L g271 ( .A(n_232), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g295 ( .A(n_232), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g333 ( .A(n_232), .B(n_258), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
AND2x2_ASAP7_75t_L g261 ( .A(n_234), .B(n_258), .Y(n_261) );
AND2x2_ASAP7_75t_L g276 ( .A(n_234), .B(n_236), .Y(n_276) );
BUFx2_ASAP7_75t_L g332 ( .A(n_234), .Y(n_332) );
AND2x2_ASAP7_75t_L g346 ( .A(n_234), .B(n_257), .Y(n_346) );
INVx2_ASAP7_75t_L g258 ( .A(n_236), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_238), .B(n_242), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g294 ( .A1(n_244), .A2(n_295), .B1(n_297), .B2(n_301), .Y(n_294) );
INVx2_ASAP7_75t_SL g325 ( .A(n_244), .Y(n_325) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
AND2x2_ASAP7_75t_L g300 ( .A(n_245), .B(n_253), .Y(n_300) );
INVx1_ASAP7_75t_L g407 ( .A(n_246), .Y(n_407) );
NOR3xp33_ASAP7_75t_L g247 ( .A(n_248), .B(n_280), .C(n_294), .Y(n_247) );
OAI221xp5_ASAP7_75t_SL g248 ( .A1(n_249), .A2(n_255), .B1(n_259), .B2(n_262), .C(n_264), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_254), .Y(n_250) );
INVxp67_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g308 ( .A(n_252), .Y(n_308) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_252), .Y(n_436) );
INVx1_ASAP7_75t_L g399 ( .A(n_254), .Y(n_399) );
AND2x2_ASAP7_75t_SL g409 ( .A(n_254), .B(n_278), .Y(n_409) );
INVxp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_258), .B(n_286), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
OR2x2_ASAP7_75t_L g292 ( .A(n_260), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g370 ( .A(n_260), .Y(n_370) );
AND2x2_ASAP7_75t_L g305 ( .A(n_261), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g351 ( .A(n_263), .B(n_311), .Y(n_351) );
AND2x2_ASAP7_75t_L g428 ( .A(n_263), .B(n_426), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_269), .B1(n_276), .B2(n_277), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g287 ( .A(n_268), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx2_ASAP7_75t_L g293 ( .A(n_271), .Y(n_293) );
AND2x4_ASAP7_75t_L g317 ( .A(n_271), .B(n_318), .Y(n_317) );
OAI21xp33_ASAP7_75t_SL g347 ( .A1(n_271), .A2(n_348), .B(n_349), .Y(n_347) );
AND2x2_ASAP7_75t_L g374 ( .A(n_271), .B(n_332), .Y(n_374) );
INVx2_ASAP7_75t_L g296 ( .A(n_272), .Y(n_296) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_272), .Y(n_329) );
INVx1_ASAP7_75t_SL g353 ( .A(n_273), .Y(n_353) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_L g284 ( .A(n_275), .Y(n_284) );
AND2x4_ASAP7_75t_SL g378 ( .A(n_275), .B(n_296), .Y(n_378) );
AND2x2_ASAP7_75t_L g375 ( .A(n_278), .B(n_321), .Y(n_375) );
AND2x2_ASAP7_75t_L g401 ( .A(n_278), .B(n_387), .Y(n_401) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_279), .Y(n_323) );
INVx1_ASAP7_75t_L g343 ( .A(n_279), .Y(n_343) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_287), .B1(n_290), .B2(n_292), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_285), .B(n_296), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_285), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g424 ( .A(n_285), .Y(n_424) );
INVx2_ASAP7_75t_SL g349 ( .A(n_287), .Y(n_349) );
AND2x2_ASAP7_75t_L g361 ( .A(n_289), .B(n_321), .Y(n_361) );
INVx2_ASAP7_75t_L g367 ( .A(n_289), .Y(n_367) );
INVxp33_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g326 ( .A(n_292), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_295), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g417 ( .A(n_295), .Y(n_417) );
INVx1_ASAP7_75t_L g345 ( .A(n_297), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_298), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g356 ( .A(n_300), .B(n_357), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_300), .A2(n_430), .B1(n_431), .B2(n_432), .Y(n_429) );
NOR3xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_324), .C(n_327), .Y(n_302) );
OAI221xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_307), .B1(n_309), .B2(n_313), .C(n_316), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g422 ( .A(n_307), .Y(n_422) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g391 ( .A(n_308), .B(n_357), .Y(n_391) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g322 ( .A(n_311), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g393 ( .A(n_313), .Y(n_393) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g390 ( .A(n_314), .Y(n_390) );
INVx1_ASAP7_75t_L g396 ( .A(n_315), .Y(n_396) );
OR2x2_ASAP7_75t_L g419 ( .A(n_315), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_SL g328 ( .A(n_318), .Y(n_328) );
AND2x2_ASAP7_75t_L g398 ( .A(n_318), .B(n_378), .Y(n_398) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_318), .B(n_331), .Y(n_430) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g435 ( .A(n_321), .Y(n_435) );
INVx1_ASAP7_75t_L g385 ( .A(n_323), .Y(n_385) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_329), .B(n_330), .C(n_334), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_328), .B(n_378), .Y(n_402) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_331), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g339 ( .A(n_333), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g420 ( .A(n_333), .Y(n_420) );
NAND4xp75_ASAP7_75t_L g335 ( .A(n_336), .B(n_392), .C(n_408), .D(n_429), .Y(n_335) );
NOR3x1_ASAP7_75t_L g336 ( .A(n_337), .B(n_354), .C(n_376), .Y(n_336) );
NAND4xp75_ASAP7_75t_L g337 ( .A(n_338), .B(n_344), .C(n_347), .D(n_350), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_339), .B(n_341), .Y(n_338) );
AND2x2_ASAP7_75t_L g389 ( .A(n_340), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g414 ( .A(n_341), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_SL g403 ( .A(n_346), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_362), .Y(n_354) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_358), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_368), .B(n_372), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI322xp33_ASAP7_75t_L g394 ( .A1(n_366), .A2(n_395), .A3(n_399), .B1(n_400), .B2(n_402), .C1(n_403), .C2(n_404), .Y(n_394) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_367), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_370), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_371), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_381), .C(n_383), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_388), .B1(n_389), .B2(n_391), .Y(n_383) );
NOR2xp33_ASAP7_75t_SL g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx2_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_398), .Y(n_395) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_401), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_405), .B(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g411 ( .A(n_406), .B(n_412), .Y(n_411) );
O2A1O1Ixp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_415), .C(n_418), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_411), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_421), .B1(n_423), .B2(n_425), .C(n_427), .Y(n_418) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g450 ( .A(n_441), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
AND2x6_ASAP7_75t_SL g466 ( .A(n_442), .B(n_444), .Y(n_466) );
OR2x6_ASAP7_75t_SL g469 ( .A(n_442), .B(n_443), .Y(n_469) );
OR2x2_ASAP7_75t_L g808 ( .A(n_442), .B(n_444), .Y(n_808) );
CKINVDCx16_ASAP7_75t_R g822 ( .A(n_442), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_446), .B(n_447), .Y(n_818) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_448), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
CKINVDCx11_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
CKINVDCx8_ASAP7_75t_R g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_456), .B(n_809), .Y(n_455) );
INVx1_ASAP7_75t_L g810 ( .A(n_457), .Y(n_810) );
CKINVDCx6p67_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
INVx4_ASAP7_75t_SL g813 ( .A(n_464), .Y(n_813) );
INVx3_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
CKINVDCx11_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
OAI22x1_ASAP7_75t_L g811 ( .A1(n_469), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_811) );
INVx1_ASAP7_75t_L g814 ( .A(n_470), .Y(n_814) );
OR3x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_672), .C(n_743), .Y(n_470) );
NAND3x1_ASAP7_75t_SL g471 ( .A(n_472), .B(n_599), .C(n_621), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_589), .Y(n_472) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_474), .A2(n_520), .B1(n_567), .B2(n_571), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_474), .A2(n_775), .B1(n_776), .B2(n_778), .Y(n_774) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_495), .Y(n_474) );
AND2x2_ASAP7_75t_L g590 ( .A(n_475), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_475), .B(n_637), .Y(n_656) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g574 ( .A(n_476), .Y(n_574) );
AND2x2_ASAP7_75t_L g624 ( .A(n_476), .B(n_497), .Y(n_624) );
INVx1_ASAP7_75t_L g663 ( .A(n_476), .Y(n_663) );
OR2x2_ASAP7_75t_L g700 ( .A(n_476), .B(n_512), .Y(n_700) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_476), .Y(n_712) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_476), .Y(n_736) );
AND2x2_ASAP7_75t_L g793 ( .A(n_476), .B(n_620), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_484), .Y(n_477) );
INVx1_ASAP7_75t_L g544 ( .A(n_479), .Y(n_544) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g580 ( .A(n_480), .Y(n_580) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
OR2x6_ASAP7_75t_L g492 ( .A(n_481), .B(n_489), .Y(n_492) );
INVxp33_ASAP7_75t_L g554 ( .A(n_481), .Y(n_554) );
INVx1_ASAP7_75t_L g581 ( .A(n_483), .Y(n_581) );
INVxp67_ASAP7_75t_L g542 ( .A(n_485), .Y(n_542) );
NOR2x1p5_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g555 ( .A(n_488), .Y(n_555) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_492), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_500) );
INVxp67_ASAP7_75t_L g533 ( .A(n_492), .Y(n_533) );
INVx2_ASAP7_75t_L g587 ( .A(n_492), .Y(n_587) );
NOR2x1_ASAP7_75t_L g495 ( .A(n_496), .B(n_510), .Y(n_495) );
INVx1_ASAP7_75t_L g668 ( .A(n_496), .Y(n_668) );
AND2x2_ASAP7_75t_L g694 ( .A(n_496), .B(n_512), .Y(n_694) );
NAND2x1_ASAP7_75t_L g710 ( .A(n_496), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g591 ( .A(n_497), .B(n_577), .Y(n_591) );
INVx3_ASAP7_75t_L g620 ( .A(n_497), .Y(n_620) );
NOR2x1_ASAP7_75t_SL g739 ( .A(n_497), .B(n_512), .Y(n_739) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_504), .B(n_509), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_503), .B(n_535), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B1(n_507), .B2(n_508), .Y(n_504) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_510), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g618 ( .A(n_511), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx4_ASAP7_75t_L g588 ( .A(n_512), .Y(n_588) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_512), .Y(n_633) );
AND2x2_ASAP7_75t_L g705 ( .A(n_512), .B(n_577), .Y(n_705) );
AND2x4_ASAP7_75t_L g722 ( .A(n_512), .B(n_666), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g769 ( .A(n_512), .B(n_664), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_512), .B(n_573), .Y(n_798) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_520), .A2(n_615), .B1(n_686), .B2(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_545), .Y(n_520) );
INVx2_ASAP7_75t_L g688 ( .A(n_521), .Y(n_688) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_529), .Y(n_521) );
BUFx3_ASAP7_75t_L g678 ( .A(n_522), .Y(n_678) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_523), .B(n_547), .Y(n_570) );
INVx2_ASAP7_75t_L g594 ( .A(n_523), .Y(n_594) );
INVx1_ASAP7_75t_L g606 ( .A(n_523), .Y(n_606) );
AND2x4_ASAP7_75t_L g613 ( .A(n_523), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g630 ( .A(n_523), .B(n_530), .Y(n_630) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_523), .Y(n_644) );
INVxp67_ASAP7_75t_L g652 ( .A(n_523), .Y(n_652) );
AND2x2_ASAP7_75t_L g681 ( .A(n_529), .B(n_597), .Y(n_681) );
AND2x2_ASAP7_75t_L g697 ( .A(n_529), .B(n_598), .Y(n_697) );
NOR2xp67_ASAP7_75t_L g784 ( .A(n_529), .B(n_597), .Y(n_784) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g593 ( .A(n_530), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g604 ( .A(n_530), .Y(n_604) );
INVx1_ASAP7_75t_L g617 ( .A(n_530), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_530), .B(n_559), .Y(n_654) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_538), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_542), .B1(n_543), .B2(n_544), .Y(n_538) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g777 ( .A(n_545), .Y(n_777) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_558), .Y(n_545) );
AND2x2_ASAP7_75t_L g651 ( .A(n_546), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g680 ( .A(n_546), .Y(n_680) );
AND2x2_ASAP7_75t_L g782 ( .A(n_546), .B(n_597), .Y(n_782) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_547), .B(n_559), .Y(n_642) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B(n_557), .Y(n_547) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_548), .A2(n_549), .B(n_557), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_550), .B(n_556), .Y(n_549) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g568 ( .A(n_558), .Y(n_568) );
NAND2x1p5_ASAP7_75t_L g757 ( .A(n_558), .B(n_678), .Y(n_757) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_559), .Y(n_671) );
AND2x2_ASAP7_75t_L g698 ( .A(n_559), .B(n_644), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g612 ( .A(n_568), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g628 ( .A(n_568), .Y(n_628) );
AND2x2_ASAP7_75t_L g716 ( .A(n_568), .B(n_593), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_568), .B(n_736), .Y(n_741) );
AND2x2_ASAP7_75t_L g751 ( .A(n_568), .B(n_630), .Y(n_751) );
OR2x2_ASAP7_75t_L g788 ( .A(n_568), .B(n_688), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_569), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g748 ( .A(n_569), .B(n_604), .Y(n_748) );
AND2x2_ASAP7_75t_L g764 ( .A(n_569), .B(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g758 ( .A(n_570), .B(n_654), .Y(n_758) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
INVx1_ASAP7_75t_L g640 ( .A(n_572), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_572), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g738 ( .A(n_572), .B(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_572), .B(n_619), .Y(n_763) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_573), .Y(n_610) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_574), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_575), .A2(n_608), .B1(n_626), .B2(n_629), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_575), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g742 ( .A(n_575), .Y(n_742) );
AND2x4_ASAP7_75t_SL g575 ( .A(n_576), .B(n_588), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g619 ( .A(n_577), .B(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g639 ( .A(n_577), .Y(n_639) );
INVx1_ASAP7_75t_L g666 ( .A(n_577), .Y(n_666) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .C(n_582), .Y(n_579) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_588), .Y(n_608) );
AND2x4_ASAP7_75t_L g665 ( .A(n_588), .B(n_666), .Y(n_665) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_588), .B(n_695), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
AND2x2_ASAP7_75t_L g690 ( .A(n_590), .B(n_633), .Y(n_690) );
OAI21xp5_ASAP7_75t_L g770 ( .A1(n_590), .A2(n_771), .B(n_772), .Y(n_770) );
INVx2_ASAP7_75t_L g648 ( .A(n_591), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_592), .A2(n_702), .B1(n_706), .B2(n_709), .Y(n_701) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_593), .Y(n_659) );
AND2x2_ASAP7_75t_L g669 ( .A(n_593), .B(n_670), .Y(n_669) );
INVx3_ASAP7_75t_L g708 ( .A(n_593), .Y(n_708) );
NAND2x1_ASAP7_75t_SL g733 ( .A(n_593), .B(n_602), .Y(n_733) );
AND2x2_ASAP7_75t_L g629 ( .A(n_595), .B(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_597), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g602 ( .A(n_598), .Y(n_602) );
INVx2_ASAP7_75t_L g614 ( .A(n_598), .Y(n_614) );
AOI21xp5_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_607), .B(n_611), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_602), .B(n_796), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_603), .A2(n_692), .B1(n_696), .B2(n_699), .Y(n_691) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
BUFx2_ASAP7_75t_L g796 ( .A(n_604), .Y(n_796) );
INVx1_ASAP7_75t_SL g803 ( .A(n_604), .Y(n_803) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_605), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OA21x2_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .B(n_618), .Y(n_611) );
AND2x2_ASAP7_75t_L g615 ( .A(n_613), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g657 ( .A(n_613), .B(n_653), .Y(n_657) );
AND2x2_ASAP7_75t_L g772 ( .A(n_613), .B(n_670), .Y(n_772) );
AND2x2_ASAP7_75t_L g775 ( .A(n_613), .B(n_681), .Y(n_775) );
AND2x4_ASAP7_75t_L g783 ( .A(n_613), .B(n_784), .Y(n_783) );
OAI21xp33_ASAP7_75t_L g737 ( .A1(n_615), .A2(n_738), .B(n_740), .Y(n_737) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g765 ( .A(n_617), .Y(n_765) );
AND2x2_ASAP7_75t_L g781 ( .A(n_617), .B(n_782), .Y(n_781) );
INVx4_ASAP7_75t_L g695 ( .A(n_619), .Y(n_695) );
INVx1_ASAP7_75t_L g664 ( .A(n_620), .Y(n_664) );
AND2x2_ASAP7_75t_L g686 ( .A(n_620), .B(n_639), .Y(n_686) );
NOR2x1_ASAP7_75t_L g621 ( .A(n_622), .B(n_645), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B(n_631), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_624), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_SL g785 ( .A(n_624), .B(n_637), .Y(n_785) );
AND2x2_ASAP7_75t_L g806 ( .A(n_624), .B(n_722), .Y(n_806) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g732 ( .A(n_629), .Y(n_732) );
OAI21xp5_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_634), .B(n_641), .Y(n_631) );
OR2x6_ASAP7_75t_L g684 ( .A(n_633), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_640), .Y(n_635) );
INVx2_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OR2x2_ASAP7_75t_L g707 ( .A(n_642), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g804 ( .A(n_642), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_643), .B(n_777), .Y(n_776) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_658), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_655), .B2(n_657), .Y(n_646) );
OR2x2_ASAP7_75t_L g718 ( .A(n_648), .B(n_719), .Y(n_718) );
INVx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_650), .Y(n_675) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g724 ( .A(n_653), .Y(n_724) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_667), .B2(n_669), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .Y(n_661) );
AND2x4_ASAP7_75t_SL g662 ( .A(n_663), .B(n_664), .Y(n_662) );
AND2x2_ASAP7_75t_L g667 ( .A(n_665), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g728 ( .A(n_668), .B(n_722), .Y(n_728) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_673), .B(n_713), .Y(n_672) );
NOR2xp67_ASAP7_75t_L g673 ( .A(n_674), .B(n_687), .Y(n_673) );
AOI21xp33_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_676), .B(n_682), .Y(n_674) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2x1p5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI22xp33_ASAP7_75t_SL g752 ( .A1(n_684), .A2(n_753), .B1(n_755), .B2(n_758), .Y(n_752) );
NOR2x1_ASAP7_75t_L g699 ( .A(n_685), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g735 ( .A(n_686), .B(n_736), .Y(n_735) );
OAI211xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B(n_691), .C(n_701), .Y(n_687) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp33_ASAP7_75t_SL g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVxp33_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g704 ( .A(n_695), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_696), .A2(n_716), .B1(n_717), .B2(n_720), .C(n_723), .Y(n_715) );
AND2x4_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g756 ( .A(n_697), .Y(n_756) );
INVx2_ASAP7_75t_SL g754 ( .A(n_700), .Y(n_754) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
NAND2x1_ASAP7_75t_L g753 ( .A(n_704), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g750 ( .A(n_710), .Y(n_750) );
INVx1_ASAP7_75t_L g779 ( .A(n_711), .Y(n_779) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NOR2x1_ASAP7_75t_L g713 ( .A(n_714), .B(n_729), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_727), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g768 ( .A(n_719), .Y(n_768) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g789 ( .A(n_722), .B(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g794 ( .A(n_722), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVxp33_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
BUFx2_ASAP7_75t_L g747 ( .A(n_726), .Y(n_747) );
OAI21xp5_ASAP7_75t_SL g729 ( .A1(n_730), .A2(n_734), .B(n_737), .Y(n_729) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx2_ASAP7_75t_L g790 ( .A(n_736), .Y(n_790) );
AND2x2_ASAP7_75t_L g778 ( .A(n_739), .B(n_779), .Y(n_778) );
NOR2xp33_ASAP7_75t_R g740 ( .A(n_741), .B(n_742), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_759), .C(n_786), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_752), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_746), .B(n_749), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
OR2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_773), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_761), .B(n_770), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_764), .B1(n_766), .B2(n_767), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NOR2x1_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_769), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g773 ( .A(n_774), .B(n_780), .Y(n_773) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_783), .B(n_785), .Y(n_780) );
INVx1_ASAP7_75t_L g799 ( .A(n_783), .Y(n_799) );
AOI211xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_789), .B(n_791), .C(n_800), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_795), .B1(n_797), .B2(n_799), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_805), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
INVxp67_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g825 ( .A(n_816), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
AND2x4_ASAP7_75t_SL g817 ( .A(n_818), .B(n_819), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
endmodule