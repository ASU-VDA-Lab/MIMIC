module fake_jpeg_16892_n_378 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_40),
.B(n_51),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_17),
.B(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_22),
.Y(n_56)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_14),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_37),
.Y(n_93)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_29),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_35),
.B(n_26),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_68),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_69),
.B(n_71),
.Y(n_166)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_73),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_38),
.B(n_18),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_36),
.Y(n_79)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_35),
.B(n_33),
.C(n_31),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_82),
.A2(n_24),
.B(n_3),
.C(n_4),
.Y(n_149)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_16),
.B1(n_27),
.B2(n_29),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_111),
.B1(n_23),
.B2(n_21),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_43),
.B(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_1),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_42),
.B(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

CKINVDCx9p33_ASAP7_75t_R g99 ( 
.A(n_50),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_56),
.A2(n_58),
.B1(n_49),
.B2(n_61),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_112),
.B1(n_25),
.B2(n_21),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_56),
.A2(n_26),
.B1(n_37),
.B2(n_30),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_41),
.A2(n_37),
.B1(n_30),
.B2(n_19),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_39),
.A2(n_16),
.B1(n_27),
.B2(n_30),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_19),
.Y(n_122)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_121),
.A2(n_136),
.B1(n_163),
.B2(n_9),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_122),
.B(n_11),
.Y(n_178)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_125),
.A2(n_75),
.B1(n_83),
.B2(n_106),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_63),
.B1(n_60),
.B2(n_59),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_127),
.A2(n_129),
.B1(n_134),
.B2(n_141),
.Y(n_174)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_111),
.B1(n_112),
.B2(n_91),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_72),
.A2(n_54),
.B1(n_25),
.B2(n_23),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_23),
.B1(n_21),
.B2(n_19),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_143),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_96),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_28),
.B1(n_24),
.B2(n_4),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_77),
.B(n_45),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_145),
.B(n_9),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_153),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_150),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_77),
.B(n_45),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_154),
.A2(n_94),
.B1(n_105),
.B2(n_89),
.Y(n_186)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_75),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_159)
);

OAI22x1_ASAP7_75t_L g202 ( 
.A1(n_159),
.A2(n_12),
.B1(n_154),
.B2(n_134),
.Y(n_202)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_73),
.B(n_5),
.C(n_6),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_107),
.C(n_110),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_83),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_96),
.B(n_7),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_145),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_108),
.Y(n_181)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_74),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_120),
.A2(n_90),
.B(n_10),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_169),
.A2(n_196),
.B(n_198),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_172),
.A2(n_175),
.B1(n_202),
.B2(n_198),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_179),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_177),
.B(n_197),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_178),
.B(n_199),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_SL g180 ( 
.A(n_131),
.B(n_74),
.C(n_70),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g244 ( 
.A(n_180),
.B(n_213),
.C(n_171),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_193),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_118),
.A2(n_108),
.B1(n_106),
.B2(n_94),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_182),
.A2(n_140),
.B1(n_162),
.B2(n_132),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_70),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_183),
.B(n_190),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_202),
.B1(n_126),
.B2(n_135),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_120),
.B(n_89),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_213),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_133),
.B(n_105),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_107),
.B(n_110),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_192),
.A2(n_210),
.B(n_178),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_129),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_125),
.A2(n_102),
.B(n_12),
.C(n_13),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_11),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_102),
.C(n_11),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_151),
.C(n_147),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_205),
.B(n_206),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_138),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_153),
.A2(n_119),
.B1(n_165),
.B2(n_155),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_210),
.B1(n_142),
.B2(n_123),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_145),
.A2(n_160),
.B1(n_157),
.B2(n_156),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_179),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_124),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_215),
.A2(n_217),
.B1(n_222),
.B2(n_228),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_161),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_216),
.B(n_226),
.C(n_208),
.Y(n_266)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_219),
.B(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_142),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_235),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_167),
.B(n_152),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_244),
.B(n_253),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_174),
.A2(n_126),
.B1(n_135),
.B2(n_158),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_174),
.A2(n_152),
.B1(n_140),
.B2(n_150),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_232),
.B1(n_228),
.B2(n_209),
.Y(n_265)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_230),
.Y(n_255)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_234),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_132),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_241),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_201),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_242),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_189),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_247),
.B(n_215),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_169),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_250),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_249),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_193),
.Y(n_248)
);

INVx13_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_251),
.Y(n_280)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_241),
.Y(n_283)
);

A2O1A1O1Ixp25_ASAP7_75t_L g253 ( 
.A1(n_196),
.A2(n_180),
.B(n_172),
.C(n_175),
.D(n_177),
.Y(n_253)
);

AND2x6_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_197),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_256),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_258),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_186),
.B(n_194),
.C(n_191),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_259),
.A2(n_265),
.B1(n_249),
.B2(n_260),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_178),
.B1(n_173),
.B2(n_176),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_200),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_262),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_173),
.B(n_194),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_286),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_267),
.C(n_282),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_204),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_275),
.B1(n_277),
.B2(n_286),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_223),
.B(n_204),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_270),
.A2(n_278),
.B1(n_261),
.B2(n_263),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_203),
.B(n_208),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_240),
.A2(n_203),
.B1(n_229),
.B2(n_223),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_224),
.A2(n_235),
.B1(n_236),
.B2(n_214),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_220),
.A2(n_230),
.B1(n_238),
.B2(n_221),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_216),
.A2(n_231),
.B(n_226),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_225),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_252),
.A2(n_233),
.B1(n_234),
.B2(n_237),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_303),
.C(n_306),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_280),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_283),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_302),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_293),
.A2(n_299),
.B1(n_310),
.B2(n_312),
.Y(n_314)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_295),
.B(n_296),
.Y(n_320)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_297),
.A2(n_304),
.B(n_291),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_276),
.B1(n_256),
.B2(n_269),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_301),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_279),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_305),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_266),
.C(n_278),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_275),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_254),
.C(n_255),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_272),
.B1(n_259),
.B2(n_263),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_264),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_258),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_272),
.A2(n_259),
.B1(n_262),
.B2(n_271),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_259),
.A2(n_284),
.B1(n_257),
.B2(n_255),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_310),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_254),
.C(n_273),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_316),
.B(n_324),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_322),
.C(n_323),
.Y(n_338)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_319),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_321),
.A2(n_329),
.B(n_327),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_257),
.C(n_284),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_280),
.C(n_259),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_301),
.Y(n_324)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_281),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_328),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_281),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_305),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_298),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_299),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_304),
.C(n_307),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_294),
.B1(n_300),
.B2(n_308),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_334),
.A2(n_339),
.B1(n_341),
.B2(n_344),
.Y(n_352)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_327),
.A2(n_293),
.B1(n_294),
.B2(n_313),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_323),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_329),
.A2(n_289),
.B(n_308),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_289),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_347),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_314),
.A2(n_291),
.B1(n_295),
.B2(n_296),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_333),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_287),
.C(n_317),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_338),
.C(n_317),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_331),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_326),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_325),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_315),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_350),
.B(n_353),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_355),
.C(n_359),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_341),
.A2(n_318),
.B1(n_314),
.B2(n_333),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_340),
.B(n_332),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_360),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_358),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_328),
.Y(n_359)
);

NOR3xp33_ASAP7_75t_L g364 ( 
.A(n_357),
.B(n_348),
.C(n_334),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_364),
.B(n_365),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_356),
.Y(n_365)
);

AOI21x1_ASAP7_75t_L g367 ( 
.A1(n_363),
.A2(n_352),
.B(n_345),
.Y(n_367)
);

AOI322xp5_ASAP7_75t_L g372 ( 
.A1(n_367),
.A2(n_369),
.A3(n_342),
.B1(n_335),
.B2(n_343),
.C1(n_344),
.C2(n_354),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_362),
.A2(n_349),
.B1(n_360),
.B2(n_347),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_361),
.B(n_336),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_370),
.B(n_366),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_371),
.B(n_372),
.Y(n_373)
);

NAND4xp25_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_368),
.C(n_367),
.D(n_355),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_359),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_375),
.B(n_346),
.C(n_351),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_335),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_343),
.Y(n_378)
);


endmodule