module fake_aes_4794_n_476 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_476);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_476;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_73;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g71 ( .A(n_17), .Y(n_71) );
INVxp33_ASAP7_75t_L g72 ( .A(n_44), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_16), .Y(n_73) );
CKINVDCx20_ASAP7_75t_R g74 ( .A(n_58), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_60), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_18), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_64), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_67), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_32), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_51), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_25), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_17), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_63), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_50), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_42), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_31), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_15), .Y(n_87) );
INVx2_ASAP7_75t_SL g88 ( .A(n_33), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_21), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_8), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_46), .Y(n_91) );
OR2x2_ASAP7_75t_L g92 ( .A(n_0), .B(n_66), .Y(n_92) );
INVx2_ASAP7_75t_SL g93 ( .A(n_11), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_43), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_24), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_3), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_4), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_5), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_15), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_56), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_20), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_62), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_52), .Y(n_103) );
AND2x2_ASAP7_75t_L g104 ( .A(n_90), .B(n_0), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_93), .B(n_1), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g106 ( .A(n_88), .B(n_1), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_74), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_87), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_89), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_102), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_102), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_88), .B(n_2), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_82), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_75), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_82), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_77), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_77), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_71), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_71), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_72), .B(n_2), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_79), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_99), .B(n_3), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_93), .B(n_4), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_80), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_110), .B(n_86), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_111), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_120), .B(n_99), .Y(n_129) );
INVx2_ASAP7_75t_SL g130 ( .A(n_120), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_119), .B(n_101), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_112), .B(n_91), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_119), .B(n_124), .Y(n_133) );
INVxp67_ASAP7_75t_SL g134 ( .A(n_104), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_111), .Y(n_135) );
NAND3x1_ASAP7_75t_L g136 ( .A(n_104), .B(n_73), .C(n_98), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_124), .B(n_73), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_111), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_124), .B(n_76), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_115), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_104), .B(n_76), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_117), .B(n_97), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_116), .B(n_94), .Y(n_143) );
AO22x2_ASAP7_75t_L g144 ( .A1(n_106), .A2(n_92), .B1(n_103), .B2(n_100), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_115), .Y(n_145) );
INVx4_ASAP7_75t_SL g146 ( .A(n_117), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_116), .A2(n_98), .B1(n_97), .B2(n_96), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_118), .B(n_92), .Y(n_148) );
INVx4_ASAP7_75t_L g149 ( .A(n_115), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_118), .B(n_85), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_123), .B(n_103), .Y(n_151) );
NOR3xp33_ASAP7_75t_SL g152 ( .A(n_127), .B(n_114), .C(n_107), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_134), .B(n_126), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_128), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_133), .B(n_125), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_135), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_133), .B(n_122), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_128), .Y(n_158) );
BUFx10_ASAP7_75t_L g159 ( .A(n_133), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_133), .B(n_126), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_128), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_135), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_148), .B(n_123), .Y(n_163) );
NOR2xp33_ASAP7_75t_R g164 ( .A(n_130), .B(n_108), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_138), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_128), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_151), .B(n_121), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
NAND2x1p5_ASAP7_75t_L g169 ( .A(n_149), .B(n_106), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_130), .B(n_105), .Y(n_170) );
NOR2x1_ASAP7_75t_L g171 ( .A(n_143), .B(n_125), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_151), .B(n_121), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
INVx5_ASAP7_75t_L g174 ( .A(n_128), .Y(n_174) );
INVx4_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_151), .B(n_121), .Y(n_176) );
INVxp67_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
NOR2xp67_ASAP7_75t_L g179 ( .A(n_151), .B(n_113), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_145), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_138), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_132), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_131), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_184), .A2(n_136), .B1(n_144), .B2(n_141), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_157), .A2(n_144), .B1(n_137), .B2(n_141), .Y(n_186) );
OR2x6_ASAP7_75t_L g187 ( .A(n_163), .B(n_136), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_167), .A2(n_137), .B(n_139), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_177), .A2(n_147), .B(n_122), .C(n_105), .Y(n_189) );
BUFx2_ASAP7_75t_L g190 ( .A(n_173), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_173), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_173), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_177), .Y(n_193) );
OR2x2_ASAP7_75t_L g194 ( .A(n_163), .B(n_109), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_SL g195 ( .A1(n_167), .A2(n_140), .B(n_80), .C(n_81), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_153), .B(n_137), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_160), .B(n_139), .Y(n_198) );
NOR2xp67_ASAP7_75t_L g199 ( .A(n_183), .B(n_129), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_164), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_153), .B(n_129), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_160), .B(n_142), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_171), .B(n_129), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_168), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_168), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_172), .A2(n_176), .B(n_170), .Y(n_206) );
INVx1_ASAP7_75t_SL g207 ( .A(n_159), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_157), .B(n_139), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_171), .B(n_139), .Y(n_209) );
BUFx2_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_157), .B(n_142), .Y(n_211) );
BUFx2_ASAP7_75t_L g212 ( .A(n_168), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_157), .A2(n_144), .B1(n_142), .B2(n_113), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_159), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_159), .B(n_142), .Y(n_215) );
OR2x2_ASAP7_75t_L g216 ( .A(n_155), .B(n_150), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_196), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_191), .Y(n_218) );
OAI21x1_ASAP7_75t_L g219 ( .A1(n_213), .A2(n_161), .B(n_154), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_202), .B(n_159), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g221 ( .A1(n_185), .A2(n_179), .B1(n_172), .B2(n_176), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_200), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g223 ( .A1(n_187), .A2(n_144), .B1(n_169), .B2(n_156), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_187), .A2(n_179), .B1(n_169), .B2(n_165), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_204), .Y(n_225) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_186), .A2(n_161), .B(n_166), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_195), .A2(n_156), .B(n_162), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_205), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_194), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_191), .Y(n_230) );
CKINVDCx14_ASAP7_75t_R g231 ( .A(n_194), .Y(n_231) );
INVx6_ASAP7_75t_L g232 ( .A(n_191), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_201), .B(n_181), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_210), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_190), .Y(n_235) );
NAND3xp33_ASAP7_75t_SL g236 ( .A(n_189), .B(n_152), .C(n_169), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_210), .Y(n_237) );
BUFx4f_ASAP7_75t_SL g238 ( .A(n_198), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_202), .B(n_181), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_212), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_225), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_239), .B(n_208), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_239), .B(n_208), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_228), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_217), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_233), .B(n_187), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_233), .B(n_208), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_228), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_225), .Y(n_249) );
OAI221xp5_ASAP7_75t_SL g250 ( .A1(n_231), .A2(n_187), .B1(n_201), .B2(n_197), .C(n_193), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_222), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_217), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_225), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_227), .A2(n_195), .B(n_206), .Y(n_254) );
AOI221xp5_ASAP7_75t_SL g255 ( .A1(n_221), .A2(n_188), .B1(n_203), .B2(n_209), .C(n_211), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_217), .Y(n_256) );
AOI21x1_ASAP7_75t_L g257 ( .A1(n_227), .A2(n_162), .B(n_165), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_223), .A2(n_198), .B1(n_199), .B2(n_190), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_218), .B(n_191), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_234), .Y(n_260) );
NAND3xp33_ASAP7_75t_L g261 ( .A(n_255), .B(n_224), .C(n_152), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_241), .B(n_230), .Y(n_262) );
OAI332xp33_ASAP7_75t_L g263 ( .A1(n_244), .A2(n_216), .A3(n_81), .B1(n_100), .B2(n_84), .B3(n_83), .C1(n_229), .C2(n_95), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_241), .B(n_230), .Y(n_264) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_254), .A2(n_226), .B(n_219), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_241), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_249), .B(n_230), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_257), .A2(n_226), .B(n_219), .Y(n_268) );
NOR3xp33_ASAP7_75t_SL g269 ( .A(n_250), .B(n_236), .C(n_83), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_249), .Y(n_270) );
OAI321xp33_ASAP7_75t_L g271 ( .A1(n_250), .A2(n_236), .A3(n_235), .B1(n_84), .B2(n_237), .C(n_234), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_244), .B(n_237), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_249), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_246), .B(n_235), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_253), .B(n_226), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_253), .Y(n_276) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_257), .A2(n_219), .B(n_218), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_251), .B(n_238), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_246), .B(n_240), .Y(n_279) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_247), .A2(n_198), .B1(n_220), .B2(n_216), .C(n_240), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_253), .Y(n_281) );
INVx5_ASAP7_75t_L g282 ( .A(n_245), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_273), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_270), .B(n_248), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_263), .B(n_260), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_270), .B(n_248), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_266), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_275), .B(n_252), .Y(n_288) );
NAND3xp33_ASAP7_75t_SL g289 ( .A(n_269), .B(n_258), .C(n_261), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_273), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_263), .B(n_242), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_273), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_276), .B(n_256), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_281), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_269), .A2(n_258), .B1(n_246), .B2(n_247), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_272), .B(n_242), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_281), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_272), .B(n_242), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_280), .B(n_243), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_280), .A2(n_243), .B1(n_220), .B2(n_259), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_281), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_274), .B(n_256), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_262), .B(n_264), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_262), .B(n_256), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_262), .B(n_252), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_275), .B(n_252), .Y(n_306) );
INVxp67_ASAP7_75t_L g307 ( .A(n_278), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_275), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_264), .B(n_267), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_279), .B(n_243), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_277), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_282), .B(n_252), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_313), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_284), .B(n_279), .Y(n_315) );
NOR2xp33_ASAP7_75t_R g316 ( .A(n_289), .B(n_5), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_308), .B(n_282), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_308), .B(n_265), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_303), .B(n_274), .Y(n_319) );
OR2x4_ASAP7_75t_L g320 ( .A(n_302), .B(n_271), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_303), .B(n_265), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_284), .B(n_264), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_286), .B(n_267), .Y(n_323) );
INVx1_ASAP7_75t_SL g324 ( .A(n_309), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_309), .B(n_265), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_286), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_285), .A2(n_261), .B(n_271), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_297), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_287), .Y(n_329) );
NOR3xp33_ASAP7_75t_SL g330 ( .A(n_295), .B(n_78), .C(n_254), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_288), .B(n_265), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_283), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_288), .B(n_265), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_288), .B(n_268), .Y(n_334) );
NOR2xp67_ASAP7_75t_SL g335 ( .A(n_290), .B(n_282), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_302), .B(n_268), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_292), .Y(n_337) );
OAI33xp33_ASAP7_75t_L g338 ( .A1(n_307), .A2(n_6), .A3(n_7), .B1(n_8), .B2(n_9), .B3(n_10), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_313), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_296), .B(n_255), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_291), .A2(n_259), .B1(n_169), .B2(n_252), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_292), .B(n_268), .Y(n_342) );
NOR2xp67_ASAP7_75t_L g343 ( .A(n_283), .B(n_282), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_298), .B(n_282), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_294), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_294), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_288), .B(n_277), .Y(n_347) );
AOI221xp5_ASAP7_75t_SL g348 ( .A1(n_310), .A2(n_6), .B1(n_7), .B2(n_9), .C(n_10), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_306), .B(n_282), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_306), .B(n_282), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_299), .B(n_259), .Y(n_351) );
INVx3_ASAP7_75t_SL g352 ( .A(n_313), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_283), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_301), .B(n_245), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_313), .Y(n_355) );
NOR3xp33_ASAP7_75t_L g356 ( .A(n_338), .B(n_218), .C(n_311), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_324), .B(n_306), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_316), .A2(n_300), .B1(n_306), .B2(n_305), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_326), .B(n_305), .Y(n_359) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_320), .A2(n_301), .B1(n_245), .B2(n_312), .Y(n_360) );
AOI32xp33_ASAP7_75t_L g361 ( .A1(n_321), .A2(n_293), .A3(n_304), .B1(n_311), .B2(n_312), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_328), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_335), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_329), .Y(n_364) );
AOI322xp5_ASAP7_75t_L g365 ( .A1(n_348), .A2(n_304), .A3(n_293), .B1(n_13), .B2(n_14), .C1(n_16), .C2(n_18), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_327), .A2(n_259), .B1(n_218), .B2(n_232), .Y(n_366) );
AOI321xp33_ASAP7_75t_SL g367 ( .A1(n_355), .A2(n_11), .A3(n_12), .B1(n_13), .B2(n_14), .C(n_19), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_352), .B(n_12), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_346), .Y(n_369) );
OAI322xp33_ASAP7_75t_SL g370 ( .A1(n_315), .A2(n_181), .A3(n_180), .B1(n_178), .B2(n_214), .C1(n_28), .C2(n_29), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_319), .B(n_259), .Y(n_371) );
NAND2x1_ASAP7_75t_L g372 ( .A(n_335), .B(n_245), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_322), .B(n_245), .Y(n_373) );
NOR3xp33_ASAP7_75t_L g374 ( .A(n_340), .B(n_207), .C(n_212), .Y(n_374) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_351), .A2(n_245), .B(n_217), .Y(n_375) );
NOR2x1_ASAP7_75t_L g376 ( .A(n_343), .B(n_217), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_332), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g378 ( .A1(n_320), .A2(n_217), .B1(n_232), .B2(n_192), .Y(n_378) );
NAND2x1_ASAP7_75t_L g379 ( .A(n_314), .B(n_232), .Y(n_379) );
OAI21xp5_ASAP7_75t_L g380 ( .A1(n_330), .A2(n_215), .B(n_180), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_337), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_345), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_352), .B(n_232), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_323), .B(n_180), .Y(n_384) );
AOI322xp5_ASAP7_75t_L g385 ( .A1(n_321), .A2(n_215), .A3(n_178), .B1(n_192), .B2(n_182), .C1(n_166), .C2(n_161), .Y(n_385) );
NOR3xp33_ASAP7_75t_L g386 ( .A(n_344), .B(n_178), .C(n_166), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_349), .Y(n_387) );
OAI21xp33_ASAP7_75t_L g388 ( .A1(n_325), .A2(n_192), .B(n_154), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_320), .B(n_22), .Y(n_389) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_332), .Y(n_390) );
OAI311xp33_ASAP7_75t_L g391 ( .A1(n_341), .A2(n_23), .A3(n_26), .B1(n_27), .C1(n_30), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_336), .Y(n_392) );
A2O1A1Ixp33_ASAP7_75t_L g393 ( .A1(n_314), .A2(n_192), .B(n_196), .C(n_182), .Y(n_393) );
OAI211xp5_ASAP7_75t_SL g394 ( .A1(n_314), .A2(n_154), .B(n_35), .C(n_36), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_317), .A2(n_232), .B1(n_182), .B2(n_196), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_339), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_339), .A2(n_196), .B1(n_182), .B2(n_174), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_325), .B(n_182), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_377), .Y(n_399) );
NOR2xp33_ASAP7_75t_R g400 ( .A(n_396), .B(n_339), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_362), .B(n_318), .Y(n_401) );
A2O1A1Ixp33_ASAP7_75t_L g402 ( .A1(n_361), .A2(n_317), .B(n_350), .C(n_349), .Y(n_402) );
NOR3xp33_ASAP7_75t_SL g403 ( .A(n_368), .B(n_317), .C(n_350), .Y(n_403) );
OAI33xp33_ASAP7_75t_L g404 ( .A1(n_392), .A2(n_342), .A3(n_354), .B1(n_353), .B2(n_318), .B3(n_333), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_387), .B(n_334), .Y(n_405) );
NAND3xp33_ASAP7_75t_L g406 ( .A(n_374), .B(n_342), .C(n_347), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_357), .B(n_334), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_359), .B(n_347), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_390), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_363), .B(n_331), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_364), .Y(n_411) );
NAND2x1_ASAP7_75t_L g412 ( .A(n_376), .B(n_175), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_381), .B(n_34), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_374), .A2(n_182), .B1(n_158), .B2(n_174), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_382), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_369), .B(n_37), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_383), .Y(n_417) );
NOR3xp33_ASAP7_75t_SL g418 ( .A(n_389), .B(n_38), .C(n_39), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_390), .B(n_40), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_358), .B(n_41), .Y(n_420) );
NOR2xp33_ASAP7_75t_SL g421 ( .A(n_386), .B(n_175), .Y(n_421) );
NAND2x1p5_ASAP7_75t_L g422 ( .A(n_372), .B(n_174), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_398), .Y(n_423) );
NOR2xp33_ASAP7_75t_R g424 ( .A(n_370), .B(n_45), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_393), .A2(n_174), .B(n_158), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_386), .A2(n_174), .B1(n_158), .B2(n_49), .Y(n_426) );
INVx3_ASAP7_75t_SL g427 ( .A(n_384), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_373), .B(n_47), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_371), .B(n_48), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_356), .B(n_53), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_400), .B(n_360), .Y(n_431) );
XOR2x2_ASAP7_75t_L g432 ( .A(n_427), .B(n_367), .Y(n_432) );
AOI322xp5_ASAP7_75t_L g433 ( .A1(n_403), .A2(n_356), .A3(n_378), .B1(n_366), .B2(n_388), .C1(n_375), .C2(n_365), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_411), .Y(n_434) );
NAND4xp75_ASAP7_75t_L g435 ( .A(n_403), .B(n_395), .C(n_380), .D(n_391), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g436 ( .A(n_430), .B(n_394), .C(n_397), .Y(n_436) );
OA22x2_ASAP7_75t_L g437 ( .A1(n_427), .A2(n_379), .B1(n_385), .B2(n_394), .Y(n_437) );
XOR2xp5_ASAP7_75t_L g438 ( .A(n_417), .B(n_54), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_402), .B(n_158), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_414), .B(n_158), .C(n_175), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_420), .B(n_55), .C(n_57), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_415), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_423), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_423), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_404), .A2(n_59), .B1(n_61), .B2(n_65), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_399), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_401), .B(n_68), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_445), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_445), .B(n_444), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_444), .B(n_401), .Y(n_451) );
NAND3x1_ASAP7_75t_SL g452 ( .A(n_437), .B(n_424), .C(n_404), .Y(n_452) );
AOI21xp33_ASAP7_75t_SL g453 ( .A1(n_437), .A2(n_420), .B(n_422), .Y(n_453) );
AOI221xp5_ASAP7_75t_SL g454 ( .A1(n_439), .A2(n_414), .B1(n_405), .B2(n_424), .C(n_407), .Y(n_454) );
NOR2xp33_ASAP7_75t_R g455 ( .A(n_448), .B(n_421), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_438), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_431), .B(n_408), .Y(n_457) );
OA22x2_ASAP7_75t_L g458 ( .A1(n_446), .A2(n_410), .B1(n_408), .B2(n_428), .Y(n_458) );
OAI31xp33_ASAP7_75t_L g459 ( .A1(n_436), .A2(n_410), .A3(n_422), .B(n_419), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_432), .A2(n_429), .B1(n_413), .B2(n_416), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_436), .A2(n_426), .B1(n_425), .B2(n_412), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_435), .A2(n_418), .B1(n_70), .B2(n_69), .Y(n_462) );
OAI221xp5_ASAP7_75t_L g463 ( .A1(n_433), .A2(n_146), .B1(n_441), .B2(n_442), .C(n_440), .Y(n_463) );
AO22x2_ASAP7_75t_L g464 ( .A1(n_443), .A2(n_444), .B1(n_406), .B2(n_434), .Y(n_464) );
OAI22xp33_ASAP7_75t_L g465 ( .A1(n_447), .A2(n_437), .B1(n_446), .B2(n_427), .Y(n_465) );
NOR3xp33_ASAP7_75t_SL g466 ( .A(n_465), .B(n_463), .C(n_459), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_453), .B(n_454), .Y(n_467) );
OAI221xp5_ASAP7_75t_R g468 ( .A1(n_460), .A2(n_454), .B1(n_452), .B2(n_462), .C(n_458), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_450), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_469), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_467), .B(n_449), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_470), .Y(n_472) );
INVxp33_ASAP7_75t_L g473 ( .A(n_471), .Y(n_473) );
XNOR2x1_ASAP7_75t_L g474 ( .A(n_473), .B(n_456), .Y(n_474) );
AOI322xp5_ASAP7_75t_L g475 ( .A1(n_474), .A2(n_472), .A3(n_466), .B1(n_468), .B2(n_457), .C1(n_451), .C2(n_461), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_475), .A2(n_472), .B1(n_464), .B2(n_459), .C(n_455), .Y(n_476) );
endmodule