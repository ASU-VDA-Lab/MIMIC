module fake_jpeg_1927_n_134 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_0),
.Y(n_55)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_47),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_39),
.C(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_42),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_53),
.B1(n_49),
.B2(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_53),
.B1(n_49),
.B2(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_67),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_59),
.Y(n_67)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_40),
.B(n_38),
.C(n_36),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_41),
.B(n_37),
.C(n_3),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_46),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_82),
.B1(n_83),
.B2(n_89),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_51),
.B(n_52),
.C(n_33),
.Y(n_81)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_18),
.B(n_30),
.C(n_28),
.D(n_27),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_49),
.B1(n_48),
.B2(n_52),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_52),
.B1(n_38),
.B2(n_46),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_1),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_78),
.C(n_69),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_31),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.C(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_104),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_73),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_105),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_2),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_8),
.B(n_9),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_5),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_16),
.B1(n_26),
.B2(n_25),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_6),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_7),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_113),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_8),
.C(n_9),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_11),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_122),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_126),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_112),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_107),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_114),
.B(n_115),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_125),
.B(n_124),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_128),
.B(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_118),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_SL g132 ( 
.A(n_131),
.B(n_118),
.C(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_12),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_12),
.Y(n_134)
);


endmodule