module fake_netlist_5_1441_n_2953 (n_137, n_294, n_431, n_318, n_380, n_419, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_631, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_637, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_644, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_639, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2953);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_644;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_639;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2953;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_2899;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_1462;
wire n_854;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1547;
wire n_1070;
wire n_777;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1561;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_1600;
wire n_845;
wire n_663;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_1587;
wire n_680;
wire n_1473;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2932;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_2919;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_2930;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_870;
wire n_931;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_744;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_2320;
wire n_2339;
wire n_1045;
wire n_1208;
wire n_2473;
wire n_2038;
wire n_2137;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_2941;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_1119;
wire n_2261;
wire n_1240;
wire n_2156;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_2929;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2933;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_912;
wire n_968;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_2916;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_1636;
wire n_894;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_2935;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_2722;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_2924;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2926;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_698;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_2284;
wire n_2187;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_2654;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_2884;
wire n_1268;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_2950;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2774;
wire n_2726;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_2208;
wire n_1404;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_2809;
wire n_2050;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_722;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_2940;
wire n_1546;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_2918;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1996;
wire n_1879;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_2938;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_1089;
wire n_927;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_33),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_610),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_523),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_369),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_535),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_505),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_9),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_492),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_360),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_532),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_376),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_489),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_210),
.Y(n_657)
);

BUFx8_ASAP7_75t_SL g658 ( 
.A(n_437),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_431),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_276),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_177),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_387),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_497),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_495),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_358),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_75),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_498),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_379),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_4),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_206),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_217),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_166),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_637),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_256),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_153),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_237),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_611),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_496),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_415),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_121),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_328),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_133),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_467),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_89),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_506),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_487),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_500),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_597),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_551),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_569),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_338),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_98),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_493),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_496),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_393),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_358),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_507),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_511),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_322),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_438),
.Y(n_700)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_243),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_192),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_372),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_112),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_105),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_403),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_330),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_57),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_448),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_472),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_506),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_455),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_477),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_570),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_188),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_522),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_356),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_604),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_415),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_147),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_471),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_482),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_318),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_526),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_449),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_223),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_493),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_464),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_275),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_275),
.Y(n_730)
);

BUFx2_ASAP7_75t_R g731 ( 
.A(n_262),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_240),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_503),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_371),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_102),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_91),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_305),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_491),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_123),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_179),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_355),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_625),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_113),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_592),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_434),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_502),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_573),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_151),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_288),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_212),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_642),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_489),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_368),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_240),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_245),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_425),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_114),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_209),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_345),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_398),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_43),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_494),
.Y(n_762)
);

BUFx5_ASAP7_75t_L g763 ( 
.A(n_445),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_37),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_101),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_508),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_95),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_350),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_344),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_328),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_377),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_582),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_346),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_56),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_453),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_201),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_466),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_639),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_55),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_261),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_4),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_410),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_488),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_374),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_143),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_290),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_386),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_562),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_614),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_218),
.Y(n_790)
);

CKINVDCx12_ASAP7_75t_R g791 ( 
.A(n_579),
.Y(n_791)
);

BUFx5_ASAP7_75t_L g792 ( 
.A(n_224),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_312),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_464),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_8),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_435),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_147),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_330),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_237),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_563),
.Y(n_800)
);

CKINVDCx14_ASAP7_75t_R g801 ( 
.A(n_601),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_499),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_137),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_209),
.Y(n_804)
);

BUFx10_ASAP7_75t_L g805 ( 
.A(n_636),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_507),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_47),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_557),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_207),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_96),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_494),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_276),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_635),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_131),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_16),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_512),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_590),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_351),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_504),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_185),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_195),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_406),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_450),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_298),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_41),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_266),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_588),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_381),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_501),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_71),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_302),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_174),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_431),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_251),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_626),
.Y(n_835)
);

BUFx5_ASAP7_75t_L g836 ( 
.A(n_138),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_142),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_215),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_78),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_15),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_121),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_435),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_43),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_24),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_519),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_280),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_509),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_583),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_398),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_543),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_51),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_7),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_295),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_368),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_476),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_287),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_386),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_333),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_134),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_333),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_619),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_490),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_153),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_411),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_388),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_640),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_164),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_524),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_552),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_404),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_229),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_528),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_227),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_297),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_14),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_172),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_124),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_424),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_248),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_403),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_353),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_111),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_515),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_20),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_621),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_497),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_279),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_484),
.Y(n_888)
);

CKINVDCx16_ASAP7_75t_R g889 ( 
.A(n_317),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_176),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_427),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_215),
.Y(n_892)
);

BUFx10_ASAP7_75t_L g893 ( 
.A(n_542),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_424),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_7),
.Y(n_895)
);

CKINVDCx16_ASAP7_75t_R g896 ( 
.A(n_701),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_763),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_763),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_658),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_763),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_763),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_763),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_885),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_763),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_763),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_658),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_889),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_645),
.Y(n_908)
);

CKINVDCx16_ASAP7_75t_R g909 ( 
.A(n_801),
.Y(n_909)
);

INVxp33_ASAP7_75t_L g910 ( 
.A(n_785),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_792),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_648),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_736),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_792),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_651),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_792),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_792),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_649),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_677),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_690),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_792),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_792),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_657),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_792),
.Y(n_924)
);

CKINVDCx16_ASAP7_75t_R g925 ( 
.A(n_801),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_836),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_836),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_724),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_742),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_836),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_688),
.B(n_1),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_744),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_836),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_836),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_747),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_772),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_683),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_800),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_836),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_827),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_797),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_835),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_845),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_848),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_850),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_836),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_832),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_735),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_735),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_861),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_736),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_735),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_866),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_773),
.Y(n_954)
);

INVxp33_ASAP7_75t_SL g955 ( 
.A(n_652),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_773),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_657),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_726),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_653),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_660),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_781),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_781),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_662),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_663),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_664),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_654),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_654),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_669),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_671),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_674),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_798),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_676),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_735),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_868),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_798),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_874),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_874),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_659),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_746),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_878),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_878),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_720),
.B(n_729),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_678),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_872),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_869),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_869),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_737),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_737),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_718),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_737),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_737),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_679),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_666),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_829),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_829),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_659),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_829),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_987),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_988),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_994),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_918),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_919),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_983),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_995),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_948),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_948),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_949),
.Y(n_1007)
);

INVxp33_ASAP7_75t_SL g1008 ( 
.A(n_899),
.Y(n_1008)
);

INVxp67_ASAP7_75t_SL g1009 ( 
.A(n_966),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_907),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_989),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_923),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_981),
.Y(n_1013)
);

CKINVDCx16_ASAP7_75t_R g1014 ( 
.A(n_896),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_949),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_920),
.B(n_778),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_952),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_923),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_952),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_973),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_973),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_990),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_957),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_928),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_957),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_990),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_955),
.B(n_647),
.Y(n_1027)
);

CKINVDCx16_ASAP7_75t_R g1028 ( 
.A(n_909),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_991),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_978),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_991),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_929),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_978),
.Y(n_1033)
);

INVxp33_ASAP7_75t_SL g1034 ( 
.A(n_906),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_955),
.B(n_778),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_996),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_996),
.Y(n_1037)
);

INVxp67_ASAP7_75t_SL g1038 ( 
.A(n_966),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_906),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_R g1040 ( 
.A(n_932),
.B(n_718),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_907),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_935),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_997),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_936),
.B(n_673),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_938),
.Y(n_1045)
);

INVxp33_ASAP7_75t_SL g1046 ( 
.A(n_940),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_997),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_951),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_954),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_942),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_956),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_943),
.Y(n_1052)
);

NOR2xp67_ASAP7_75t_L g1053 ( 
.A(n_944),
.B(n_646),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_958),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_945),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_950),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_953),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_974),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_961),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_979),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_962),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_971),
.Y(n_1062)
);

INVxp33_ASAP7_75t_SL g1063 ( 
.A(n_984),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1009),
.B(n_967),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1048),
.Y(n_1065)
);

AND2x2_ASAP7_75t_R g1066 ( 
.A(n_1040),
.B(n_731),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1019),
.B(n_897),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_1019),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_998),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1013),
.B(n_1038),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1049),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1051),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_1044),
.B(n_1016),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1059),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_999),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_1061),
.Y(n_1076)
);

AOI22x1_ASAP7_75t_SL g1077 ( 
.A1(n_1018),
.A2(n_675),
.B1(n_770),
.B2(n_712),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_1062),
.B(n_967),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1000),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_1054),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1004),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_1005),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_1006),
.Y(n_1083)
);

CKINVDCx11_ASAP7_75t_R g1084 ( 
.A(n_1018),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_1007),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1015),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1017),
.Y(n_1087)
);

CKINVDCx8_ASAP7_75t_R g1088 ( 
.A(n_1014),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1020),
.B(n_901),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1021),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1022),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_SL g1092 ( 
.A(n_1027),
.B(n_883),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1026),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_1029),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_1003),
.B(n_925),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1031),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_1053),
.B(n_913),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_1043),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_1054),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_1001),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1047),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1035),
.B(n_908),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1010),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1002),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_1046),
.B(n_908),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_1028),
.B(n_941),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1024),
.A2(n_712),
.B1(n_770),
.B2(n_675),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1032),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1045),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_1052),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1055),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1056),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_1057),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1058),
.B(n_913),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_1060),
.Y(n_1115)
);

AND2x6_ASAP7_75t_L g1116 ( 
.A(n_1063),
.B(n_673),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1042),
.B(n_902),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1050),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1060),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1041),
.B(n_975),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1008),
.B(n_904),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_L g1122 ( 
.A(n_1041),
.B(n_883),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_1011),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1039),
.B(n_947),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1039),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1034),
.B(n_905),
.Y(n_1126)
);

INVx4_ASAP7_75t_L g1127 ( 
.A(n_1012),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1023),
.B(n_976),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1023),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1025),
.B(n_903),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1025),
.B(n_977),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1030),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1030),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_1033),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_1033),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1036),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_1036),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1037),
.B(n_980),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1037),
.A2(n_810),
.B1(n_814),
.B2(n_783),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_1019),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1048),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1019),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1019),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1009),
.B(n_982),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1019),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1048),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1019),
.B(n_911),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_1001),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1019),
.Y(n_1149)
);

AOI22x1_ASAP7_75t_SL g1150 ( 
.A1(n_1018),
.A2(n_810),
.B1(n_814),
.B2(n_783),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1048),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1019),
.Y(n_1152)
);

INVxp33_ASAP7_75t_SL g1153 ( 
.A(n_1040),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1065),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1073),
.B(n_992),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1064),
.B(n_689),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1071),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1149),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1072),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_1128),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1074),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1141),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1152),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1143),
.Y(n_1164)
);

OA21x2_ASAP7_75t_L g1165 ( 
.A1(n_1067),
.A2(n_916),
.B(n_914),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1146),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1114),
.B(n_869),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1080),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1068),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1073),
.B(n_912),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1151),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1106),
.B(n_912),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1143),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1145),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1102),
.B(n_915),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1145),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1068),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1079),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1102),
.B(n_915),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1094),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1064),
.B(n_959),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1068),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1094),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1070),
.B(n_959),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1097),
.B(n_1144),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1140),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1097),
.B(n_960),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1099),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1076),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1076),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1115),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1114),
.B(n_869),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1140),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1126),
.B(n_1121),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1144),
.B(n_960),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1078),
.B(n_716),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1075),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1140),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1067),
.A2(n_921),
.B(n_917),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1119),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1142),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1142),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1142),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1075),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1147),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1078),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1147),
.A2(n_1089),
.B(n_1081),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1126),
.A2(n_788),
.B1(n_751),
.B2(n_931),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1121),
.B(n_963),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_1116),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1069),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1086),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1087),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1075),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1090),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1091),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1093),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1116),
.B(n_969),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1096),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1092),
.B(n_751),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_1124),
.Y(n_1221)
);

AND2x6_ASAP7_75t_L g1222 ( 
.A(n_1111),
.B(n_788),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1101),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1089),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1082),
.B(n_1098),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1082),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1082),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1098),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1098),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1083),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1083),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1083),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1083),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1085),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1085),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1085),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1085),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1117),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1117),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1116),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1110),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1116),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1116),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1110),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1103),
.Y(n_1245)
);

NAND2xp33_ASAP7_75t_L g1246 ( 
.A(n_1110),
.B(n_789),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1128),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1131),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1131),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1120),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1110),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1138),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1138),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1120),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1112),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1132),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1092),
.B(n_992),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1130),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1153),
.B(n_963),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1104),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1108),
.Y(n_1261)
);

XNOR2xp5_ASAP7_75t_L g1262 ( 
.A(n_1134),
.B(n_964),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1095),
.A2(n_900),
.B(n_898),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1080),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1105),
.B(n_964),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1095),
.B(n_965),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1105),
.B(n_965),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1109),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1113),
.B(n_808),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1153),
.B(n_968),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1113),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1113),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1113),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1100),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1122),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1100),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1088),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1132),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1118),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1107),
.B(n_968),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1129),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1084),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1136),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1148),
.Y(n_1284)
);

AND2x6_ASAP7_75t_L g1285 ( 
.A(n_1132),
.B(n_813),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1107),
.B(n_969),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1132),
.B(n_817),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1133),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1133),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1133),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1139),
.A2(n_840),
.B1(n_860),
.B2(n_818),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1133),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1262),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1158),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1224),
.B(n_1205),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1225),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1220),
.A2(n_1238),
.B1(n_1239),
.B2(n_1194),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1205),
.B(n_922),
.Y(n_1298)
);

OAI22x1_ASAP7_75t_L g1299 ( 
.A1(n_1175),
.A2(n_1125),
.B1(n_1127),
.B2(n_1123),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_1241),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1244),
.Y(n_1301)
);

AND2x6_ASAP7_75t_L g1302 ( 
.A(n_1243),
.B(n_1137),
.Y(n_1302)
);

BUFx10_ASAP7_75t_L g1303 ( 
.A(n_1209),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1158),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1225),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1163),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1163),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1220),
.A2(n_686),
.B1(n_762),
.B2(n_668),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1264),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1225),
.Y(n_1310)
);

XOR2xp5_ASAP7_75t_R g1311 ( 
.A(n_1291),
.B(n_1066),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1154),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1212),
.Y(n_1313)
);

NAND2xp33_ASAP7_75t_L g1314 ( 
.A(n_1243),
.B(n_1244),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1244),
.B(n_1127),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1197),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1188),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1194),
.B(n_924),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1197),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1157),
.Y(n_1320)
);

NAND3xp33_ASAP7_75t_L g1321 ( 
.A(n_1175),
.B(n_972),
.C(n_970),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1179),
.B(n_970),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1155),
.B(n_1139),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1159),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_SL g1325 ( 
.A(n_1241),
.B(n_818),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1212),
.Y(n_1326)
);

AND2x6_ASAP7_75t_L g1327 ( 
.A(n_1243),
.B(n_1137),
.Y(n_1327)
);

OR2x6_ASAP7_75t_L g1328 ( 
.A(n_1244),
.B(n_937),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1251),
.Y(n_1329)
);

OAI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1170),
.A2(n_972),
.B1(n_910),
.B2(n_860),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1251),
.B(n_805),
.Y(n_1331)
);

NAND2xp33_ASAP7_75t_L g1332 ( 
.A(n_1243),
.B(n_927),
.Y(n_1332)
);

AND2x2_ASAP7_75t_SL g1333 ( 
.A(n_1179),
.B(n_1077),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1209),
.B(n_1135),
.Y(n_1334)
);

XNOR2xp5_ASAP7_75t_L g1335 ( 
.A(n_1282),
.B(n_1150),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1161),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1251),
.B(n_805),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1251),
.B(n_805),
.Y(n_1338)
);

AND2x6_ASAP7_75t_L g1339 ( 
.A(n_1240),
.B(n_1242),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1162),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1216),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1216),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1260),
.B(n_893),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1168),
.B(n_993),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1180),
.B(n_930),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1180),
.B(n_933),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1278),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1183),
.B(n_934),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1219),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1208),
.A2(n_714),
.B1(n_946),
.B2(n_939),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1166),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1260),
.B(n_893),
.Y(n_1352)
);

AND2x6_ASAP7_75t_L g1353 ( 
.A(n_1240),
.B(n_1242),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1267),
.B(n_1084),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1171),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1178),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1268),
.B(n_893),
.Y(n_1357)
);

NOR3xp33_ASAP7_75t_L g1358 ( 
.A(n_1259),
.B(n_1135),
.C(n_719),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1219),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1278),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1164),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1183),
.B(n_1255),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1213),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1164),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1215),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1265),
.B(n_759),
.Y(n_1366)
);

INVx6_ASAP7_75t_L g1367 ( 
.A(n_1278),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1217),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1223),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1173),
.Y(n_1370)
);

OAI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1268),
.A2(n_840),
.B1(n_765),
.B2(n_710),
.Y(n_1371)
);

BUFx4f_ASAP7_75t_L g1372 ( 
.A(n_1278),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1197),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1288),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1258),
.B(n_666),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1173),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1174),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1266),
.B(n_733),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1185),
.A2(n_768),
.B1(n_825),
.B2(n_771),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1174),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1176),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1197),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1204),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1176),
.Y(n_1384)
);

INVx4_ASAP7_75t_L g1385 ( 
.A(n_1288),
.Y(n_1385)
);

INVxp33_ASAP7_75t_L g1386 ( 
.A(n_1172),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1288),
.Y(n_1387)
);

BUFx4f_ASAP7_75t_L g1388 ( 
.A(n_1288),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1195),
.B(n_666),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1255),
.B(n_985),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1191),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1177),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1287),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1177),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1204),
.Y(n_1395)
);

BUFx4f_ASAP7_75t_L g1396 ( 
.A(n_1284),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1211),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1206),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1261),
.B(n_985),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1182),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1184),
.B(n_985),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1182),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1165),
.B(n_898),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1186),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1204),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1165),
.B(n_900),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1156),
.A2(n_926),
.B1(n_829),
.B2(n_769),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1156),
.A2(n_926),
.B1(n_791),
.B2(n_839),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1156),
.A2(n_794),
.B1(n_864),
.B2(n_754),
.Y(n_1409)
);

AOI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1230),
.A2(n_655),
.B(n_650),
.Y(n_1410)
);

BUFx10_ASAP7_75t_L g1411 ( 
.A(n_1269),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1186),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1165),
.B(n_831),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1198),
.Y(n_1414)
);

NOR3xp33_ASAP7_75t_L g1415 ( 
.A(n_1259),
.B(n_681),
.C(n_680),
.Y(n_1415)
);

BUFx4f_ASAP7_75t_L g1416 ( 
.A(n_1277),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1198),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1201),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1201),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1256),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1204),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1226),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1287),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1271),
.B(n_656),
.Y(n_1424)
);

INVx8_ASAP7_75t_L g1425 ( 
.A(n_1285),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1189),
.A2(n_884),
.B1(n_754),
.B2(n_887),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1256),
.B(n_884),
.Y(n_1427)
);

INVx5_ASAP7_75t_L g1428 ( 
.A(n_1285),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1207),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1227),
.Y(n_1430)
);

OR2x6_ASAP7_75t_L g1431 ( 
.A(n_1249),
.B(n_661),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1228),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1160),
.Y(n_1433)
);

INVxp33_ASAP7_75t_L g1434 ( 
.A(n_1200),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1287),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1190),
.A2(n_891),
.B1(n_892),
.B2(n_890),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1289),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1229),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1289),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1214),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1221),
.B(n_682),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1207),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1232),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1196),
.A2(n_667),
.B1(n_670),
.B2(n_665),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1232),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1236),
.Y(n_1446)
);

INVx5_ASAP7_75t_L g1447 ( 
.A(n_1285),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1257),
.B(n_685),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1214),
.B(n_985),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1236),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1231),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1199),
.B(n_672),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1169),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1214),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1214),
.B(n_986),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1233),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1237),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1199),
.B(n_684),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1234),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1181),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1290),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1199),
.B(n_691),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1235),
.B(n_693),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1234),
.Y(n_1464)
);

INVx4_ASAP7_75t_L g1465 ( 
.A(n_1234),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1269),
.B(n_986),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1292),
.Y(n_1467)
);

CKINVDCx11_ASAP7_75t_R g1468 ( 
.A(n_1281),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1169),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1169),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1202),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1279),
.Y(n_1472)
);

NOR3xp33_ASAP7_75t_L g1473 ( 
.A(n_1270),
.B(n_692),
.C(n_687),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1202),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1270),
.B(n_695),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1235),
.B(n_694),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1234),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1202),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1250),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1203),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1249),
.B(n_1252),
.Y(n_1481)
);

INVx6_ASAP7_75t_L g1482 ( 
.A(n_1269),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1203),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1167),
.B(n_700),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1203),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1193),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1193),
.Y(n_1487)
);

INVxp67_ASAP7_75t_SL g1488 ( 
.A(n_1250),
.Y(n_1488)
);

INVxp33_ASAP7_75t_SL g1489 ( 
.A(n_1160),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1280),
.B(n_696),
.Y(n_1490)
);

CKINVDCx11_ASAP7_75t_R g1491 ( 
.A(n_1281),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1245),
.B(n_1250),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1283),
.B(n_702),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1167),
.B(n_704),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1329),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1313),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1312),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1326),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1320),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1309),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1341),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1295),
.B(n_1272),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1344),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1342),
.Y(n_1504)
);

NOR3xp33_ASAP7_75t_L g1505 ( 
.A(n_1366),
.B(n_1275),
.C(n_1286),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1295),
.B(n_1297),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1347),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1317),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1322),
.B(n_1460),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1324),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1347),
.Y(n_1511)
);

NOR2xp67_ASAP7_75t_L g1512 ( 
.A(n_1428),
.B(n_1447),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1336),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1323),
.B(n_1283),
.C(n_1187),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1349),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1340),
.Y(n_1516)
);

NOR3xp33_ASAP7_75t_L g1517 ( 
.A(n_1330),
.B(n_1254),
.C(n_1274),
.Y(n_1517)
);

NAND2xp33_ASAP7_75t_L g1518 ( 
.A(n_1302),
.B(n_1210),
.Y(n_1518)
);

NAND2xp33_ASAP7_75t_L g1519 ( 
.A(n_1302),
.B(n_1210),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1378),
.B(n_1273),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1460),
.B(n_1276),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1303),
.B(n_1252),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1303),
.B(n_1247),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1325),
.B(n_1248),
.Y(n_1524)
);

NOR3xp33_ASAP7_75t_L g1525 ( 
.A(n_1321),
.B(n_1253),
.C(n_1218),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1492),
.B(n_1192),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1361),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1325),
.B(n_1210),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1321),
.B(n_1192),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1362),
.B(n_1285),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1411),
.B(n_1210),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1386),
.B(n_1196),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1364),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1362),
.B(n_1285),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1489),
.B(n_1196),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1370),
.Y(n_1536)
);

NAND3xp33_ASAP7_75t_L g1537 ( 
.A(n_1490),
.B(n_1246),
.C(n_708),
.Y(n_1537)
);

XOR2xp5_ASAP7_75t_L g1538 ( 
.A(n_1293),
.B(n_516),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1376),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1351),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1377),
.Y(n_1541)
);

INVx8_ASAP7_75t_L g1542 ( 
.A(n_1302),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1448),
.B(n_1222),
.Y(n_1543)
);

NAND2xp33_ASAP7_75t_SL g1544 ( 
.A(n_1300),
.B(n_1246),
.Y(n_1544)
);

AO221x1_ASAP7_75t_L g1545 ( 
.A1(n_1371),
.A2(n_721),
.B1(n_723),
.B2(n_713),
.C(n_705),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1355),
.B(n_1222),
.Y(n_1546)
);

NOR2xp67_ASAP7_75t_L g1547 ( 
.A(n_1428),
.B(n_517),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1347),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1356),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1372),
.A2(n_1263),
.B(n_986),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1363),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1294),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1459),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1365),
.B(n_1222),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1368),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1411),
.B(n_1263),
.Y(n_1556)
);

NOR3xp33_ASAP7_75t_L g1557 ( 
.A(n_1334),
.B(n_698),
.C(n_697),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1369),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1493),
.B(n_702),
.Y(n_1559)
);

NOR2xp67_ASAP7_75t_L g1560 ( 
.A(n_1428),
.B(n_1447),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1393),
.B(n_699),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1296),
.B(n_1222),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1359),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1475),
.A2(n_732),
.B(n_734),
.C(n_727),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1434),
.B(n_703),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1304),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1296),
.B(n_1222),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1391),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1305),
.B(n_706),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1306),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1307),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1433),
.B(n_709),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1305),
.B(n_711),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1328),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1310),
.B(n_715),
.Y(n_1575)
);

INVxp33_ASAP7_75t_L g1576 ( 
.A(n_1468),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1420),
.Y(n_1577)
);

NOR2xp67_ASAP7_75t_L g1578 ( 
.A(n_1447),
.B(n_518),
.Y(n_1578)
);

INVx4_ASAP7_75t_L g1579 ( 
.A(n_1374),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1380),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1441),
.B(n_752),
.C(n_743),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1472),
.B(n_717),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1310),
.B(n_722),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1423),
.B(n_725),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1435),
.B(n_728),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1328),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1318),
.B(n_730),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1372),
.B(n_738),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1318),
.B(n_739),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1381),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_L g1591 ( 
.A(n_1415),
.B(n_786),
.C(n_784),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1389),
.B(n_1375),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1488),
.B(n_1298),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1328),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1298),
.B(n_740),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1354),
.B(n_741),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1374),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1463),
.B(n_745),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1473),
.A2(n_822),
.B1(n_824),
.B2(n_815),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1463),
.B(n_748),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1384),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1379),
.B(n_749),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1443),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1374),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1476),
.B(n_750),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1481),
.B(n_826),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1476),
.B(n_753),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1398),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_SL g1609 ( 
.A(n_1396),
.B(n_702),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1343),
.B(n_755),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1461),
.B(n_756),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1416),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1467),
.B(n_757),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1427),
.B(n_707),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1345),
.B(n_758),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1481),
.B(n_828),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1352),
.B(n_760),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_L g1618 ( 
.A(n_1302),
.B(n_886),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1357),
.B(n_761),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1427),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1416),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1345),
.B(n_764),
.Y(n_1622)
);

NOR2xp67_ASAP7_75t_L g1623 ( 
.A(n_1301),
.B(n_520),
.Y(n_1623)
);

A2O1A1Ixp33_ASAP7_75t_L g1624 ( 
.A1(n_1397),
.A2(n_833),
.B(n_843),
.C(n_830),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1388),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1445),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1491),
.B(n_766),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1446),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1388),
.Y(n_1629)
);

OAI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1482),
.A2(n_767),
.B1(n_775),
.B2(n_774),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1402),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1395),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1404),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1412),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1346),
.B(n_776),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1346),
.B(n_777),
.Y(n_1636)
);

BUFx5_ASAP7_75t_L g1637 ( 
.A(n_1339),
.Y(n_1637)
);

NOR3xp33_ASAP7_75t_L g1638 ( 
.A(n_1358),
.B(n_780),
.C(n_779),
.Y(n_1638)
);

NOR3xp33_ASAP7_75t_L g1639 ( 
.A(n_1331),
.B(n_787),
.C(n_782),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1427),
.B(n_1431),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1348),
.B(n_790),
.Y(n_1641)
);

NOR2xp67_ASAP7_75t_L g1642 ( 
.A(n_1301),
.B(n_521),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1479),
.B(n_793),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_L g1644 ( 
.A(n_1408),
.B(n_858),
.C(n_856),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1482),
.B(n_795),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1450),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1348),
.B(n_796),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1431),
.B(n_707),
.Y(n_1648)
);

NAND3xp33_ASAP7_75t_L g1649 ( 
.A(n_1408),
.B(n_802),
.C(n_799),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1417),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1392),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1419),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1394),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1431),
.B(n_707),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1424),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1395),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1400),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1395),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1422),
.B(n_803),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1413),
.B(n_804),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1424),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1414),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1337),
.B(n_807),
.C(n_806),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1418),
.Y(n_1664)
);

NOR2x1p5_ASAP7_75t_L g1665 ( 
.A(n_1437),
.B(n_809),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1413),
.B(n_811),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1479),
.B(n_1484),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1479),
.B(n_812),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1430),
.B(n_816),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_L g1670 ( 
.A(n_1350),
.B(n_1494),
.C(n_1484),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1453),
.Y(n_1671)
);

NOR3xp33_ASAP7_75t_L g1672 ( 
.A(n_1338),
.B(n_820),
.C(n_819),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1494),
.B(n_821),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1469),
.Y(n_1674)
);

INVx4_ASAP7_75t_L g1675 ( 
.A(n_1385),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1432),
.B(n_823),
.Y(n_1676)
);

NOR3xp33_ASAP7_75t_L g1677 ( 
.A(n_1315),
.B(n_837),
.C(n_834),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1396),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1451),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1299),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1385),
.B(n_1421),
.Y(n_1681)
);

NAND2x1p5_ASAP7_75t_L g1682 ( 
.A(n_1405),
.B(n_873),
.Y(n_1682)
);

INVx4_ASAP7_75t_L g1683 ( 
.A(n_1367),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1438),
.B(n_838),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1333),
.B(n_841),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1439),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1481),
.B(n_1444),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1456),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1457),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1360),
.B(n_876),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1471),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1421),
.B(n_842),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_SL g1693 ( 
.A(n_1327),
.Y(n_1693)
);

AO221x1_ASAP7_75t_L g1694 ( 
.A1(n_1316),
.A2(n_1373),
.B1(n_1383),
.B2(n_1382),
.C(n_1319),
.Y(n_1694)
);

AND2x2_ASAP7_75t_SL g1695 ( 
.A(n_1314),
.B(n_851),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1470),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1480),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1485),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1409),
.B(n_851),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1474),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1478),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1483),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1486),
.B(n_844),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1487),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1678),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1602),
.A2(n_1327),
.B1(n_1401),
.B2(n_1436),
.Y(n_1706)
);

NOR2xp67_ASAP7_75t_L g1707 ( 
.A(n_1514),
.B(n_1452),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1509),
.B(n_1520),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1505),
.A2(n_1327),
.B1(n_1308),
.B2(n_1466),
.Y(n_1709)
);

INVx4_ASAP7_75t_L g1710 ( 
.A(n_1625),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1521),
.B(n_1335),
.Y(n_1711)
);

BUFx8_ASAP7_75t_L g1712 ( 
.A(n_1693),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1625),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1595),
.B(n_1327),
.Y(n_1714)
);

NOR2xp67_ASAP7_75t_L g1715 ( 
.A(n_1568),
.B(n_1452),
.Y(n_1715)
);

NAND2xp33_ASAP7_75t_L g1716 ( 
.A(n_1625),
.B(n_1425),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1497),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1499),
.Y(n_1718)
);

A2O1A1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1529),
.A2(n_1458),
.B(n_1462),
.C(n_1425),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1510),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1577),
.Y(n_1721)
);

OR2x2_ASAP7_75t_SL g1722 ( 
.A(n_1649),
.B(n_1311),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1592),
.B(n_1421),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1587),
.B(n_1426),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1513),
.Y(n_1725)
);

INVx5_ASAP7_75t_L g1726 ( 
.A(n_1542),
.Y(n_1726)
);

AND2x2_ASAP7_75t_SL g1727 ( 
.A(n_1695),
.B(n_1609),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1589),
.B(n_1506),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1535),
.B(n_1440),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1502),
.B(n_1308),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1612),
.B(n_1387),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1500),
.B(n_1440),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1503),
.B(n_1440),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1508),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1516),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1540),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1598),
.B(n_1407),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1600),
.B(n_1454),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1596),
.B(n_1367),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1605),
.B(n_1458),
.Y(n_1740)
);

OAI21xp33_ASAP7_75t_L g1741 ( 
.A1(n_1524),
.A2(n_847),
.B(n_846),
.Y(n_1741)
);

INVxp67_ASAP7_75t_SL g1742 ( 
.A(n_1593),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1532),
.B(n_1459),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1670),
.A2(n_1462),
.B(n_1406),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1607),
.B(n_1403),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1615),
.B(n_1403),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1549),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1551),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_1544),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1495),
.B(n_1399),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1622),
.B(n_1406),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1555),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1537),
.B(n_852),
.C(n_849),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1537),
.A2(n_1353),
.B1(n_1339),
.B2(n_1425),
.Y(n_1754)
);

CKINVDCx20_ASAP7_75t_R g1755 ( 
.A(n_1538),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1517),
.A2(n_853),
.B1(n_855),
.B2(n_854),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1687),
.A2(n_857),
.B1(n_862),
.B2(n_859),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1545),
.A2(n_863),
.B1(n_867),
.B2(n_865),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1495),
.B(n_1316),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1635),
.B(n_1319),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1621),
.B(n_1459),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1559),
.B(n_1410),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1558),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1636),
.B(n_1373),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1608),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1572),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1665),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1570),
.Y(n_1768)
);

INVxp67_ASAP7_75t_SL g1769 ( 
.A(n_1518),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1571),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1655),
.B(n_1382),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1641),
.B(n_1647),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1660),
.B(n_1383),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1666),
.B(n_1464),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1673),
.B(n_1464),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1563),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1638),
.A2(n_1525),
.B1(n_1661),
.B2(n_1659),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1669),
.A2(n_870),
.B1(n_875),
.B2(n_871),
.Y(n_1778)
);

OR2x6_ASAP7_75t_L g1779 ( 
.A(n_1542),
.B(n_1405),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1557),
.A2(n_1353),
.B1(n_1339),
.B2(n_1390),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1668),
.B(n_1449),
.Y(n_1781)
);

INVxp33_ASAP7_75t_L g1782 ( 
.A(n_1565),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1522),
.B(n_1339),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1582),
.B(n_1465),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1679),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1552),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1526),
.B(n_1353),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1566),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1620),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1591),
.A2(n_1353),
.B1(n_1477),
.B2(n_1465),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1629),
.B(n_1477),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1591),
.A2(n_1332),
.B1(n_1455),
.B2(n_1442),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1688),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1580),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1590),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_SL g1796 ( 
.A(n_1693),
.B(n_1542),
.Y(n_1796)
);

NAND2x1p5_ASAP7_75t_L g1797 ( 
.A(n_1629),
.B(n_1429),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1629),
.B(n_851),
.Y(n_1798)
);

INVxp33_ASAP7_75t_L g1799 ( 
.A(n_1645),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1684),
.B(n_877),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1523),
.B(n_879),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1667),
.B(n_880),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1689),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1690),
.B(n_881),
.Y(n_1804)
);

NOR2x1_ASAP7_75t_L g1805 ( 
.A(n_1675),
.B(n_986),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1601),
.Y(n_1806)
);

BUFx12f_ASAP7_75t_L g1807 ( 
.A(n_1586),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1610),
.B(n_882),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1631),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1640),
.B(n_525),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1496),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1611),
.B(n_888),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1519),
.A2(n_529),
.B(n_527),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1690),
.B(n_894),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1685),
.A2(n_895),
.B1(n_2),
.B2(n_0),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1569),
.B(n_0),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1617),
.B(n_1),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1573),
.B(n_2),
.Y(n_1818)
);

AO22x1_ASAP7_75t_L g1819 ( 
.A1(n_1576),
.A2(n_6),
.B1(n_3),
.B2(n_5),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1633),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1575),
.B(n_3),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1594),
.B(n_5),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1686),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1574),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1630),
.B(n_6),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1583),
.B(n_8),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1543),
.A2(n_1556),
.B(n_1534),
.Y(n_1827)
);

OR2x6_ASAP7_75t_L g1828 ( 
.A(n_1675),
.B(n_530),
.Y(n_1828)
);

AND2x6_ASAP7_75t_SL g1829 ( 
.A(n_1627),
.B(n_9),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1530),
.A2(n_533),
.B(n_531),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1680),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1634),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1613),
.B(n_10),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1650),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1599),
.B(n_10),
.Y(n_1835)
);

INVx4_ASAP7_75t_L g1836 ( 
.A(n_1632),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1619),
.B(n_11),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1606),
.Y(n_1838)
);

INVx8_ASAP7_75t_L g1839 ( 
.A(n_1507),
.Y(n_1839)
);

OR2x6_ASAP7_75t_L g1840 ( 
.A(n_1512),
.B(n_534),
.Y(n_1840)
);

BUFx4_ASAP7_75t_L g1841 ( 
.A(n_1584),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1699),
.B(n_11),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1606),
.B(n_12),
.Y(n_1843)
);

NAND3xp33_ASAP7_75t_L g1844 ( 
.A(n_1581),
.B(n_12),
.C(n_13),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_R g1845 ( 
.A(n_1618),
.B(n_536),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1652),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1616),
.B(n_13),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1498),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1616),
.B(n_14),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1676),
.B(n_15),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1648),
.B(n_16),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1654),
.B(n_17),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1644),
.B(n_17),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1501),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1581),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1683),
.B(n_1704),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1644),
.A2(n_1639),
.B1(n_1672),
.B2(n_1663),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1614),
.B(n_18),
.Y(n_1858)
);

NAND2x1p5_ASAP7_75t_L g1859 ( 
.A(n_1683),
.B(n_539),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1682),
.B(n_19),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1504),
.B(n_21),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1528),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1862)
);

O2A1O1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1564),
.A2(n_1624),
.B(n_1588),
.C(n_1692),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1677),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1864)
);

AOI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1670),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1561),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1515),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1585),
.B(n_28),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1527),
.Y(n_1869)
);

INVx3_ASAP7_75t_L g1870 ( 
.A(n_1579),
.Y(n_1870)
);

O2A1O1Ixp33_ASAP7_75t_L g1871 ( 
.A1(n_1643),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1703),
.B(n_29),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1533),
.B(n_30),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1536),
.B(n_31),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1653),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1539),
.B(n_32),
.Y(n_1876)
);

NAND3xp33_ASAP7_75t_L g1877 ( 
.A(n_1546),
.B(n_34),
.C(n_35),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1541),
.B(n_34),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1651),
.B(n_35),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1664),
.B(n_1603),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1671),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1657),
.Y(n_1882)
);

AOI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1554),
.A2(n_1701),
.B1(n_1700),
.B2(n_1567),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1662),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1626),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1628),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1674),
.B(n_1696),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1646),
.B(n_36),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1691),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1632),
.B(n_38),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1702),
.B(n_39),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1632),
.B(n_39),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1697),
.B(n_40),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1656),
.B(n_40),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1698),
.A2(n_44),
.B1(n_41),
.B2(n_42),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1553),
.B(n_42),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1553),
.B(n_44),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1579),
.Y(n_1898)
);

AND2x2_ASAP7_75t_SL g1899 ( 
.A(n_1562),
.B(n_45),
.Y(n_1899)
);

INVx6_ASAP7_75t_L g1900 ( 
.A(n_1656),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1681),
.B(n_45),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1766),
.A2(n_1560),
.B1(n_1512),
.B2(n_1623),
.Y(n_1902)
);

OAI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1815),
.A2(n_1642),
.B1(n_1623),
.B2(n_1578),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1717),
.Y(n_1904)
);

A2O1A1Ixp33_ASAP7_75t_L g1905 ( 
.A1(n_1808),
.A2(n_1642),
.B(n_1547),
.C(n_1578),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1719),
.A2(n_1550),
.B(n_1531),
.Y(n_1906)
);

A2O1A1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1817),
.A2(n_1547),
.B(n_1560),
.C(n_1656),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1708),
.A2(n_1658),
.B1(n_1511),
.B2(n_1548),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1735),
.Y(n_1909)
);

AOI21x1_ASAP7_75t_L g1910 ( 
.A1(n_1707),
.A2(n_1694),
.B(n_1637),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1740),
.A2(n_1637),
.B(n_1511),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1742),
.A2(n_1637),
.B(n_1511),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1769),
.A2(n_1637),
.B(n_1548),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1802),
.B(n_1658),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1782),
.B(n_1658),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1728),
.A2(n_1637),
.B(n_1548),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1784),
.B(n_1507),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1746),
.A2(n_1597),
.B(n_1507),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1777),
.B(n_1597),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1710),
.B(n_1597),
.Y(n_1920)
);

AO21x1_ASAP7_75t_L g1921 ( 
.A1(n_1865),
.A2(n_46),
.B(n_47),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1799),
.B(n_1604),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1842),
.B(n_1604),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1899),
.B(n_1604),
.Y(n_1924)
);

AOI21x1_ASAP7_75t_L g1925 ( 
.A1(n_1827),
.A2(n_538),
.B(n_537),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1721),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1711),
.B(n_540),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1734),
.Y(n_1928)
);

INVx4_ASAP7_75t_L g1929 ( 
.A(n_1726),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1772),
.B(n_46),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1801),
.B(n_48),
.Y(n_1931)
);

AOI21x1_ASAP7_75t_L g1932 ( 
.A1(n_1751),
.A2(n_544),
.B(n_541),
.Y(n_1932)
);

O2A1O1Ixp33_ASAP7_75t_L g1933 ( 
.A1(n_1837),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_1933)
);

OAI21xp33_ASAP7_75t_L g1934 ( 
.A1(n_1850),
.A2(n_49),
.B(n_50),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1777),
.B(n_51),
.Y(n_1935)
);

AO21x2_ASAP7_75t_L g1936 ( 
.A1(n_1744),
.A2(n_546),
.B(n_545),
.Y(n_1936)
);

BUFx3_ASAP7_75t_L g1937 ( 
.A(n_1823),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1745),
.A2(n_629),
.B(n_628),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1738),
.A2(n_631),
.B(n_630),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1739),
.B(n_52),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1763),
.Y(n_1941)
);

INVx4_ASAP7_75t_L g1942 ( 
.A(n_1726),
.Y(n_1942)
);

AOI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1714),
.A2(n_633),
.B(n_632),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1810),
.B(n_52),
.Y(n_1944)
);

INVx4_ASAP7_75t_SL g1945 ( 
.A(n_1840),
.Y(n_1945)
);

AOI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1774),
.A2(n_641),
.B(n_638),
.Y(n_1946)
);

OAI21xp33_ASAP7_75t_L g1947 ( 
.A1(n_1800),
.A2(n_53),
.B(n_54),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1727),
.B(n_53),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1715),
.B(n_54),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_SL g1950 ( 
.A(n_1796),
.B(n_1712),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1872),
.B(n_55),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1863),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1705),
.B(n_547),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1726),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1749),
.B(n_548),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1779),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1773),
.A2(n_617),
.B(n_616),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1724),
.B(n_58),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1756),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1857),
.B(n_59),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1833),
.B(n_549),
.Y(n_1961)
);

O2A1O1Ixp33_ASAP7_75t_L g1962 ( 
.A1(n_1825),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1962)
);

OAI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1737),
.A2(n_553),
.B(n_550),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1810),
.B(n_62),
.Y(n_1964)
);

OAI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1787),
.A2(n_555),
.B(n_554),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1779),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1712),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1760),
.A2(n_608),
.B(n_607),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1803),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1775),
.B(n_63),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1757),
.B(n_63),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1755),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1806),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1786),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1812),
.B(n_556),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1764),
.B(n_64),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1798),
.B(n_558),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1730),
.B(n_64),
.Y(n_1978)
);

O2A1O1Ixp33_ASAP7_75t_L g1979 ( 
.A1(n_1851),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1838),
.B(n_65),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1788),
.Y(n_1981)
);

INVx2_ASAP7_75t_SL g1982 ( 
.A(n_1713),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1757),
.B(n_1741),
.Y(n_1983)
);

A2O1A1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1756),
.A2(n_1818),
.B(n_1821),
.C(n_1816),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1718),
.Y(n_1985)
);

AOI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1813),
.A2(n_622),
.B(n_620),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1868),
.B(n_559),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1824),
.B(n_1722),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1754),
.A2(n_627),
.B(n_624),
.Y(n_1989)
);

INVx4_ASAP7_75t_L g1990 ( 
.A(n_1713),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_SL g1991 ( 
.A(n_1828),
.B(n_66),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1720),
.Y(n_1992)
);

OAI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1753),
.A2(n_67),
.B(n_68),
.Y(n_1993)
);

O2A1O1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1852),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1778),
.B(n_69),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1725),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1830),
.A2(n_644),
.B(n_561),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1783),
.A2(n_643),
.B(n_564),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1706),
.A2(n_634),
.B(n_565),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1716),
.A2(n_623),
.B(n_566),
.Y(n_2000)
);

A2O1A1Ixp33_ASAP7_75t_L g2001 ( 
.A1(n_1826),
.A2(n_1758),
.B(n_1865),
.C(n_1871),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1789),
.B(n_1729),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1713),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1794),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1743),
.A2(n_618),
.B(n_567),
.Y(n_2005)
);

AO21x1_ASAP7_75t_L g2006 ( 
.A1(n_1758),
.A2(n_1853),
.B(n_1883),
.Y(n_2006)
);

AOI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_1790),
.A2(n_615),
.B(n_568),
.Y(n_2007)
);

OAI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_1709),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1778),
.B(n_72),
.Y(n_2009)
);

AOI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1792),
.A2(n_571),
.B(n_560),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1795),
.B(n_73),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1835),
.B(n_73),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1723),
.A2(n_613),
.B(n_574),
.Y(n_2013)
);

AOI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1762),
.A2(n_612),
.B(n_575),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1804),
.B(n_74),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1807),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1814),
.B(n_74),
.Y(n_2017)
);

O2A1O1Ixp33_ASAP7_75t_L g2018 ( 
.A1(n_1858),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_2018)
);

OAI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1877),
.A2(n_576),
.B(n_572),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1840),
.A2(n_609),
.B(n_578),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1840),
.A2(n_606),
.B(n_580),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1828),
.A2(n_605),
.B(n_581),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1831),
.B(n_577),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1736),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1889),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1828),
.A2(n_585),
.B(n_584),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1779),
.A2(n_587),
.B(n_586),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1856),
.B(n_76),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1747),
.Y(n_2029)
);

A2O1A1Ixp33_ASAP7_75t_L g2030 ( 
.A1(n_1864),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1748),
.B(n_79),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_1710),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1732),
.B(n_1781),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1752),
.B(n_80),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1767),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1860),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1780),
.A2(n_603),
.B(n_591),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1765),
.B(n_1785),
.Y(n_2038)
);

NOR3xp33_ASAP7_75t_L g2039 ( 
.A(n_1819),
.B(n_81),
.C(n_82),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1811),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_1844),
.A2(n_83),
.B(n_84),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1759),
.A2(n_1791),
.B(n_1887),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1797),
.A2(n_602),
.B(n_593),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_1768),
.A2(n_1776),
.B(n_1770),
.Y(n_2044)
);

INVxp67_ASAP7_75t_SL g2045 ( 
.A(n_1793),
.Y(n_2045)
);

AOI21xp33_ASAP7_75t_L g2046 ( 
.A1(n_1891),
.A2(n_83),
.B(n_84),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1809),
.A2(n_600),
.B(n_594),
.Y(n_2047)
);

BUFx8_ASAP7_75t_L g2048 ( 
.A(n_1856),
.Y(n_2048)
);

OAI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_1861),
.A2(n_85),
.B(n_86),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_1839),
.Y(n_2050)
);

O2A1O1Ixp33_ASAP7_75t_L g2051 ( 
.A1(n_1822),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1854),
.B(n_87),
.Y(n_2052)
);

CKINVDCx20_ASAP7_75t_R g2053 ( 
.A(n_1839),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1869),
.B(n_88),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1820),
.Y(n_2055)
);

INVx4_ASAP7_75t_L g2056 ( 
.A(n_1839),
.Y(n_2056)
);

INVx3_ASAP7_75t_SL g2057 ( 
.A(n_1900),
.Y(n_2057)
);

NOR3xp33_ASAP7_75t_L g2058 ( 
.A(n_1843),
.B(n_88),
.C(n_89),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1885),
.B(n_90),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1832),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1834),
.Y(n_2061)
);

NOR3xp33_ASAP7_75t_L g2062 ( 
.A(n_1847),
.B(n_90),
.C(n_91),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1846),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1880),
.A2(n_595),
.B(n_589),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1849),
.B(n_92),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_1731),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1733),
.B(n_1771),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1882),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1848),
.B(n_92),
.Y(n_2069)
);

A2O1A1Ixp33_ASAP7_75t_L g2070 ( 
.A1(n_1750),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_1972),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1937),
.Y(n_2072)
);

NAND3xp33_ASAP7_75t_SL g2073 ( 
.A(n_1984),
.B(n_1875),
.C(n_1866),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1945),
.B(n_1836),
.Y(n_2074)
);

AOI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_1905),
.A2(n_1903),
.B(n_1906),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_2042),
.B(n_1845),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2045),
.Y(n_2077)
);

AND2x4_ASAP7_75t_L g2078 ( 
.A(n_1945),
.B(n_1836),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1909),
.Y(n_2079)
);

AOI22x1_ASAP7_75t_L g2080 ( 
.A1(n_2019),
.A2(n_1859),
.B1(n_1884),
.B2(n_1867),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1978),
.B(n_1901),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1969),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1973),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1985),
.Y(n_2084)
);

INVx1_ASAP7_75t_SL g2085 ( 
.A(n_1928),
.Y(n_2085)
);

BUFx2_ASAP7_75t_L g2086 ( 
.A(n_2048),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_1927),
.B(n_1829),
.Y(n_2087)
);

HB1xp67_ASAP7_75t_SL g2088 ( 
.A(n_2048),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2025),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2060),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2061),
.Y(n_2091)
);

BUFx6f_ASAP7_75t_L g2092 ( 
.A(n_2057),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2033),
.B(n_1930),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1974),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1923),
.B(n_1897),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1958),
.B(n_1886),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1992),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1981),
.Y(n_2098)
);

INVx1_ASAP7_75t_SL g2099 ( 
.A(n_1926),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1967),
.Y(n_2100)
);

OR2x2_ASAP7_75t_SL g2101 ( 
.A(n_1951),
.B(n_1931),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1970),
.B(n_1875),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1996),
.Y(n_2103)
);

INVx3_ASAP7_75t_L g2104 ( 
.A(n_1954),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1976),
.B(n_1893),
.Y(n_2105)
);

CKINVDCx20_ASAP7_75t_R g2106 ( 
.A(n_2053),
.Y(n_2106)
);

BUFx2_ASAP7_75t_L g2107 ( 
.A(n_2066),
.Y(n_2107)
);

HB1xp67_ASAP7_75t_L g2108 ( 
.A(n_2002),
.Y(n_2108)
);

CKINVDCx11_ASAP7_75t_R g2109 ( 
.A(n_2035),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1954),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1924),
.B(n_1896),
.Y(n_2111)
);

NAND2x1p5_ASAP7_75t_L g2112 ( 
.A(n_2056),
.B(n_1870),
.Y(n_2112)
);

BUFx3_ASAP7_75t_L g2113 ( 
.A(n_1922),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1935),
.B(n_1890),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1983),
.B(n_1892),
.Y(n_2115)
);

OAI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_2001),
.A2(n_1855),
.B1(n_1862),
.B2(n_1895),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2024),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1934),
.B(n_1894),
.Y(n_2118)
);

AO22x1_ASAP7_75t_L g2119 ( 
.A1(n_2039),
.A2(n_1874),
.B1(n_1876),
.B2(n_1873),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1971),
.B(n_1878),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2029),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2055),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_R g2123 ( 
.A(n_1950),
.B(n_1870),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2063),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2068),
.Y(n_2125)
);

AND2x4_ASAP7_75t_SL g2126 ( 
.A(n_2056),
.B(n_1731),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2004),
.B(n_1904),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1941),
.B(n_1879),
.Y(n_2128)
);

BUFx3_ASAP7_75t_L g2129 ( 
.A(n_1915),
.Y(n_2129)
);

BUFx6f_ASAP7_75t_L g2130 ( 
.A(n_2003),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2038),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_1914),
.B(n_2012),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_1945),
.B(n_1898),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2065),
.B(n_1888),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1948),
.B(n_1771),
.Y(n_2135)
);

INVx1_ASAP7_75t_SL g2136 ( 
.A(n_1917),
.Y(n_2136)
);

INVx6_ASAP7_75t_L g2137 ( 
.A(n_2003),
.Y(n_2137)
);

AND2x6_ASAP7_75t_L g2138 ( 
.A(n_1956),
.B(n_1805),
.Y(n_2138)
);

INVxp67_ASAP7_75t_L g2139 ( 
.A(n_2067),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2044),
.Y(n_2140)
);

AOI22x1_ASAP7_75t_L g2141 ( 
.A1(n_2019),
.A2(n_1898),
.B1(n_1881),
.B2(n_1841),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2040),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_1975),
.B(n_1900),
.Y(n_2143)
);

INVx2_ASAP7_75t_SL g2144 ( 
.A(n_2003),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1960),
.B(n_1761),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2031),
.Y(n_2146)
);

BUFx6f_ASAP7_75t_L g2147 ( 
.A(n_1920),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1995),
.B(n_93),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2052),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2034),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2054),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2059),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_SL g2153 ( 
.A1(n_2009),
.A2(n_97),
.B1(n_94),
.B2(n_96),
.Y(n_2153)
);

AOI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_1991),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_2154)
);

BUFx8_ASAP7_75t_L g2155 ( 
.A(n_1944),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_L g2156 ( 
.A(n_1920),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1961),
.B(n_1987),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2011),
.Y(n_2158)
);

AOI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_1991),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_2159)
);

INVx2_ASAP7_75t_SL g2160 ( 
.A(n_1982),
.Y(n_2160)
);

AND2x2_ASAP7_75t_SL g2161 ( 
.A(n_1950),
.B(n_100),
.Y(n_2161)
);

CKINVDCx8_ASAP7_75t_R g2162 ( 
.A(n_2016),
.Y(n_2162)
);

AOI221xp5_ASAP7_75t_L g2163 ( 
.A1(n_1933),
.A2(n_2062),
.B1(n_2058),
.B2(n_1947),
.C(n_2049),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_1940),
.B(n_102),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_L g2165 ( 
.A(n_2050),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1919),
.B(n_103),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_1956),
.B(n_596),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2032),
.Y(n_2168)
);

AND2x2_ASAP7_75t_SL g2169 ( 
.A(n_1929),
.B(n_103),
.Y(n_2169)
);

OR2x6_ASAP7_75t_L g2170 ( 
.A(n_2022),
.B(n_2026),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2032),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_1966),
.B(n_598),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_2006),
.B(n_599),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_R g2174 ( 
.A(n_2050),
.B(n_104),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2069),
.Y(n_2175)
);

OR2x2_ASAP7_75t_SL g2176 ( 
.A(n_2015),
.B(n_104),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1990),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1936),
.Y(n_2178)
);

INVx3_ASAP7_75t_L g2179 ( 
.A(n_1929),
.Y(n_2179)
);

INVxp67_ASAP7_75t_L g2180 ( 
.A(n_1988),
.Y(n_2180)
);

BUFx3_ASAP7_75t_L g2181 ( 
.A(n_1990),
.Y(n_2181)
);

BUFx8_ASAP7_75t_L g2182 ( 
.A(n_1964),
.Y(n_2182)
);

AOI21xp5_ASAP7_75t_L g2183 ( 
.A1(n_2076),
.A2(n_1963),
.B(n_1999),
.Y(n_2183)
);

NOR2x1_ASAP7_75t_L g2184 ( 
.A(n_2140),
.B(n_1936),
.Y(n_2184)
);

BUFx2_ASAP7_75t_R g2185 ( 
.A(n_2162),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2108),
.B(n_2093),
.Y(n_2186)
);

BUFx3_ASAP7_75t_L g2187 ( 
.A(n_2092),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_2157),
.B(n_1955),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2131),
.B(n_2017),
.Y(n_2189)
);

NAND2x1p5_ASAP7_75t_L g2190 ( 
.A(n_2133),
.B(n_1966),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2090),
.Y(n_2191)
);

CKINVDCx6p67_ASAP7_75t_R g2192 ( 
.A(n_2109),
.Y(n_2192)
);

AND2x6_ASAP7_75t_SL g2193 ( 
.A(n_2087),
.B(n_1953),
.Y(n_2193)
);

OAI22xp5_ASAP7_75t_L g2194 ( 
.A1(n_2101),
.A2(n_1959),
.B1(n_2030),
.B2(n_2036),
.Y(n_2194)
);

INVx2_ASAP7_75t_SL g2195 ( 
.A(n_2072),
.Y(n_2195)
);

O2A1O1Ixp5_ASAP7_75t_L g2196 ( 
.A1(n_2173),
.A2(n_1921),
.B(n_1952),
.C(n_2041),
.Y(n_2196)
);

OAI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_2141),
.A2(n_2070),
.B1(n_2008),
.B2(n_1993),
.Y(n_2197)
);

BUFx12f_ASAP7_75t_L g2198 ( 
.A(n_2071),
.Y(n_2198)
);

O2A1O1Ixp33_ASAP7_75t_L g2199 ( 
.A1(n_2073),
.A2(n_1962),
.B(n_1994),
.C(n_1979),
.Y(n_2199)
);

O2A1O1Ixp33_ASAP7_75t_SL g2200 ( 
.A1(n_2163),
.A2(n_1949),
.B(n_2046),
.C(n_2018),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2091),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2122),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2122),
.Y(n_2203)
);

O2A1O1Ixp5_ASAP7_75t_L g2204 ( 
.A1(n_2119),
.A2(n_1963),
.B(n_1997),
.C(n_2010),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_2092),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2084),
.Y(n_2206)
);

A2O1A1Ixp33_ASAP7_75t_L g2207 ( 
.A1(n_2075),
.A2(n_1977),
.B(n_2051),
.C(n_2021),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_2077),
.B(n_2124),
.Y(n_2208)
);

INVx2_ASAP7_75t_SL g2209 ( 
.A(n_2072),
.Y(n_2209)
);

BUFx6f_ASAP7_75t_L g2210 ( 
.A(n_2092),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2124),
.Y(n_2211)
);

A2O1A1Ixp33_ASAP7_75t_L g2212 ( 
.A1(n_2116),
.A2(n_2102),
.B(n_2159),
.C(n_2154),
.Y(n_2212)
);

HAxp5_ASAP7_75t_L g2213 ( 
.A(n_2176),
.B(n_1980),
.CON(n_2213),
.SN(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2125),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_2072),
.Y(n_2215)
);

A2O1A1Ixp33_ASAP7_75t_L g2216 ( 
.A1(n_2081),
.A2(n_2020),
.B(n_2037),
.C(n_2007),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2125),
.Y(n_2217)
);

HB1xp67_ASAP7_75t_L g2218 ( 
.A(n_2107),
.Y(n_2218)
);

A2O1A1Ixp33_ASAP7_75t_SL g2219 ( 
.A1(n_2143),
.A2(n_2023),
.B(n_1965),
.C(n_1998),
.Y(n_2219)
);

BUFx2_ASAP7_75t_L g2220 ( 
.A(n_2123),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_2141),
.A2(n_2028),
.B1(n_1907),
.B2(n_1902),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2099),
.B(n_2146),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2150),
.B(n_1918),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_L g2224 ( 
.A(n_2139),
.B(n_105),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2175),
.B(n_1911),
.Y(n_2225)
);

AOI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2170),
.A2(n_1986),
.B(n_1912),
.Y(n_2226)
);

BUFx10_ASAP7_75t_L g2227 ( 
.A(n_2100),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2153),
.A2(n_1965),
.B1(n_1989),
.B2(n_1908),
.Y(n_2228)
);

INVxp33_ASAP7_75t_L g2229 ( 
.A(n_2095),
.Y(n_2229)
);

NAND3xp33_ASAP7_75t_L g2230 ( 
.A(n_2148),
.B(n_1939),
.C(n_1938),
.Y(n_2230)
);

A2O1A1Ixp33_ASAP7_75t_L g2231 ( 
.A1(n_2118),
.A2(n_2000),
.B(n_2014),
.C(n_2027),
.Y(n_2231)
);

BUFx3_ASAP7_75t_L g2232 ( 
.A(n_2113),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2097),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2103),
.Y(n_2234)
);

A2O1A1Ixp33_ASAP7_75t_L g2235 ( 
.A1(n_2114),
.A2(n_1957),
.B(n_1968),
.C(n_1946),
.Y(n_2235)
);

A2O1A1Ixp33_ASAP7_75t_L g2236 ( 
.A1(n_2105),
.A2(n_2047),
.B(n_2005),
.C(n_2013),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_2117),
.B(n_1942),
.Y(n_2237)
);

A2O1A1Ixp33_ASAP7_75t_L g2238 ( 
.A1(n_2135),
.A2(n_1943),
.B(n_2064),
.C(n_2043),
.Y(n_2238)
);

OAI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_2161),
.A2(n_1942),
.B1(n_1913),
.B2(n_1916),
.Y(n_2239)
);

BUFx3_ASAP7_75t_L g2240 ( 
.A(n_2129),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2121),
.Y(n_2241)
);

INVxp67_ASAP7_75t_SL g2242 ( 
.A(n_2178),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_SL g2243 ( 
.A(n_2169),
.Y(n_2243)
);

BUFx2_ASAP7_75t_L g2244 ( 
.A(n_2074),
.Y(n_2244)
);

CKINVDCx14_ASAP7_75t_R g2245 ( 
.A(n_2106),
.Y(n_2245)
);

OAI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_2180),
.A2(n_1910),
.B1(n_1925),
.B2(n_1932),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2149),
.B(n_106),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2202),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2186),
.B(n_2132),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2208),
.B(n_2111),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2203),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2208),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_2218),
.B(n_2074),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2223),
.B(n_2136),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_2244),
.Y(n_2255)
);

NOR2x1p5_ASAP7_75t_L g2256 ( 
.A(n_2192),
.B(n_2120),
.Y(n_2256)
);

INVxp67_ASAP7_75t_L g2257 ( 
.A(n_2241),
.Y(n_2257)
);

INVx4_ASAP7_75t_L g2258 ( 
.A(n_2215),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2211),
.Y(n_2259)
);

BUFx2_ASAP7_75t_L g2260 ( 
.A(n_2190),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2229),
.B(n_2085),
.Y(n_2261)
);

BUFx3_ASAP7_75t_L g2262 ( 
.A(n_2205),
.Y(n_2262)
);

AND2x4_ASAP7_75t_L g2263 ( 
.A(n_2214),
.B(n_2078),
.Y(n_2263)
);

AOI22xp33_ASAP7_75t_L g2264 ( 
.A1(n_2194),
.A2(n_2080),
.B1(n_2164),
.B2(n_2115),
.Y(n_2264)
);

AOI22xp33_ASAP7_75t_L g2265 ( 
.A1(n_2243),
.A2(n_2080),
.B1(n_2166),
.B2(n_2170),
.Y(n_2265)
);

OAI321xp33_ASAP7_75t_L g2266 ( 
.A1(n_2197),
.A2(n_2145),
.A3(n_2178),
.B1(n_2096),
.B2(n_2128),
.C(n_2152),
.Y(n_2266)
);

CKINVDCx14_ASAP7_75t_R g2267 ( 
.A(n_2245),
.Y(n_2267)
);

AOI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_2243),
.A2(n_2134),
.B1(n_2172),
.B2(n_2167),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2217),
.Y(n_2269)
);

AOI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_2183),
.A2(n_2207),
.B(n_2204),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2206),
.Y(n_2271)
);

AOI21xp5_ASAP7_75t_L g2272 ( 
.A1(n_2226),
.A2(n_2133),
.B(n_2151),
.Y(n_2272)
);

INVx2_ASAP7_75t_SL g2273 ( 
.A(n_2205),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2225),
.B(n_2158),
.Y(n_2274)
);

NOR2x1_ASAP7_75t_SL g2275 ( 
.A(n_2221),
.B(n_2177),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2222),
.B(n_2142),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2233),
.Y(n_2277)
);

OAI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2228),
.A2(n_2212),
.B1(n_2188),
.B2(n_2220),
.Y(n_2278)
);

OAI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_2228),
.A2(n_2088),
.B1(n_2086),
.B2(n_2078),
.Y(n_2279)
);

BUFx3_ASAP7_75t_L g2280 ( 
.A(n_2205),
.Y(n_2280)
);

HB1xp67_ASAP7_75t_L g2281 ( 
.A(n_2242),
.Y(n_2281)
);

AOI22xp33_ASAP7_75t_SL g2282 ( 
.A1(n_2230),
.A2(n_2174),
.B1(n_2182),
.B2(n_2155),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2234),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_2237),
.B(n_2104),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2191),
.Y(n_2285)
);

OAI21xp5_ASAP7_75t_L g2286 ( 
.A1(n_2270),
.A2(n_2196),
.B(n_2216),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2281),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2254),
.B(n_2201),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_2263),
.B(n_2237),
.Y(n_2289)
);

OAI21x1_ASAP7_75t_L g2290 ( 
.A1(n_2272),
.A2(n_2184),
.B(n_2239),
.Y(n_2290)
);

AOI22xp33_ASAP7_75t_SL g2291 ( 
.A1(n_2278),
.A2(n_2275),
.B1(n_2279),
.B2(n_2267),
.Y(n_2291)
);

OAI21x1_ASAP7_75t_L g2292 ( 
.A1(n_2265),
.A2(n_2184),
.B(n_2199),
.Y(n_2292)
);

AND2x4_ASAP7_75t_L g2293 ( 
.A(n_2263),
.B(n_2195),
.Y(n_2293)
);

BUFx3_ASAP7_75t_L g2294 ( 
.A(n_2262),
.Y(n_2294)
);

AO21x2_ASAP7_75t_L g2295 ( 
.A1(n_2266),
.A2(n_2246),
.B(n_2235),
.Y(n_2295)
);

OAI21x1_ASAP7_75t_L g2296 ( 
.A1(n_2265),
.A2(n_2189),
.B(n_2179),
.Y(n_2296)
);

OAI21x1_ASAP7_75t_L g2297 ( 
.A1(n_2274),
.A2(n_2179),
.B(n_2127),
.Y(n_2297)
);

BUFx3_ASAP7_75t_L g2298 ( 
.A(n_2262),
.Y(n_2298)
);

OAI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_2264),
.A2(n_2231),
.B1(n_2236),
.B2(n_2238),
.Y(n_2299)
);

BUFx2_ASAP7_75t_L g2300 ( 
.A(n_2281),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2254),
.B(n_2249),
.Y(n_2301)
);

O2A1O1Ixp5_ASAP7_75t_L g2302 ( 
.A1(n_2276),
.A2(n_2219),
.B(n_2247),
.C(n_2224),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2250),
.B(n_2209),
.Y(n_2303)
);

CKINVDCx20_ASAP7_75t_R g2304 ( 
.A(n_2267),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2255),
.B(n_2232),
.Y(n_2305)
);

BUFx2_ASAP7_75t_R g2306 ( 
.A(n_2280),
.Y(n_2306)
);

O2A1O1Ixp33_ASAP7_75t_L g2307 ( 
.A1(n_2264),
.A2(n_2200),
.B(n_2213),
.C(n_2160),
.Y(n_2307)
);

INVx3_ASAP7_75t_L g2308 ( 
.A(n_2248),
.Y(n_2308)
);

AOI22xp33_ASAP7_75t_L g2309 ( 
.A1(n_2299),
.A2(n_2282),
.B1(n_2256),
.B2(n_2260),
.Y(n_2309)
);

OAI21x1_ASAP7_75t_L g2310 ( 
.A1(n_2290),
.A2(n_2259),
.B(n_2251),
.Y(n_2310)
);

AND2x4_ASAP7_75t_L g2311 ( 
.A(n_2308),
.B(n_2284),
.Y(n_2311)
);

INVx2_ASAP7_75t_SL g2312 ( 
.A(n_2308),
.Y(n_2312)
);

BUFx3_ASAP7_75t_L g2313 ( 
.A(n_2304),
.Y(n_2313)
);

NAND2x1p5_ASAP7_75t_L g2314 ( 
.A(n_2290),
.B(n_2253),
.Y(n_2314)
);

INVx2_ASAP7_75t_SL g2315 ( 
.A(n_2294),
.Y(n_2315)
);

CKINVDCx20_ASAP7_75t_R g2316 ( 
.A(n_2305),
.Y(n_2316)
);

BUFx3_ASAP7_75t_L g2317 ( 
.A(n_2294),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2287),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2312),
.Y(n_2319)
);

BUFx2_ASAP7_75t_L g2320 ( 
.A(n_2316),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2312),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2318),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2315),
.B(n_2301),
.Y(n_2323)
);

BUFx3_ASAP7_75t_L g2324 ( 
.A(n_2313),
.Y(n_2324)
);

CKINVDCx5p33_ASAP7_75t_R g2325 ( 
.A(n_2324),
.Y(n_2325)
);

OAI21x1_ASAP7_75t_L g2326 ( 
.A1(n_2319),
.A2(n_2310),
.B(n_2314),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2322),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_2324),
.Y(n_2328)
);

INVx3_ASAP7_75t_L g2329 ( 
.A(n_2319),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_2320),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2323),
.Y(n_2331)
);

OAI21x1_ASAP7_75t_SL g2332 ( 
.A1(n_2321),
.A2(n_2315),
.B(n_2309),
.Y(n_2332)
);

OAI22xp33_ASAP7_75t_L g2333 ( 
.A1(n_2321),
.A2(n_2286),
.B1(n_2317),
.B2(n_2314),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_2330),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2330),
.B(n_2325),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2325),
.B(n_2328),
.Y(n_2336)
);

OR2x2_ASAP7_75t_L g2337 ( 
.A(n_2331),
.B(n_2288),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2328),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2328),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2328),
.B(n_2313),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2327),
.Y(n_2341)
);

INVxp67_ASAP7_75t_SL g2342 ( 
.A(n_2329),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2329),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2329),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_2334),
.B(n_2313),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2335),
.B(n_2340),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2336),
.B(n_2317),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2338),
.B(n_2339),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2342),
.B(n_2339),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2343),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2337),
.B(n_2342),
.Y(n_2351)
);

INVx1_ASAP7_75t_SL g2352 ( 
.A(n_2344),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2344),
.B(n_2317),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2349),
.Y(n_2354)
);

NOR2xp67_ASAP7_75t_L g2355 ( 
.A(n_2345),
.B(n_2343),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2349),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2345),
.B(n_2333),
.Y(n_2357)
);

OAI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2357),
.A2(n_2345),
.B(n_2346),
.Y(n_2358)
);

AND2x4_ASAP7_75t_L g2359 ( 
.A(n_2355),
.B(n_2349),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2354),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2356),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_2359),
.B(n_2346),
.Y(n_2362)
);

AND2x2_ASAP7_75t_SL g2363 ( 
.A(n_2359),
.B(n_2347),
.Y(n_2363)
);

INVxp67_ASAP7_75t_SL g2364 ( 
.A(n_2358),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2361),
.Y(n_2365)
);

OR2x2_ASAP7_75t_L g2366 ( 
.A(n_2360),
.B(n_2351),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2359),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2363),
.B(n_2348),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2366),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2362),
.B(n_2348),
.Y(n_2370)
);

OR2x2_ASAP7_75t_L g2371 ( 
.A(n_2367),
.B(n_2352),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2362),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2364),
.B(n_2347),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2365),
.B(n_2353),
.Y(n_2374)
);

INVx1_ASAP7_75t_SL g2375 ( 
.A(n_2363),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_2362),
.Y(n_2376)
);

INVxp67_ASAP7_75t_SL g2377 ( 
.A(n_2364),
.Y(n_2377)
);

AOI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2375),
.A2(n_2350),
.B1(n_2341),
.B2(n_2291),
.Y(n_2378)
);

OAI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2368),
.A2(n_2350),
.B(n_2326),
.Y(n_2379)
);

OA222x2_ASAP7_75t_L g2380 ( 
.A1(n_2376),
.A2(n_2332),
.B1(n_2187),
.B2(n_2193),
.C1(n_2185),
.C2(n_2240),
.Y(n_2380)
);

NAND4xp75_ASAP7_75t_L g2381 ( 
.A(n_2373),
.B(n_2302),
.C(n_2286),
.D(n_2312),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2368),
.B(n_2318),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_2376),
.B(n_2326),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2372),
.B(n_2261),
.Y(n_2384)
);

OAI21xp5_ASAP7_75t_L g2385 ( 
.A1(n_2377),
.A2(n_2370),
.B(n_2371),
.Y(n_2385)
);

O2A1O1Ixp33_ASAP7_75t_L g2386 ( 
.A1(n_2377),
.A2(n_2307),
.B(n_2193),
.C(n_2314),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2370),
.Y(n_2387)
);

AOI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_2369),
.A2(n_2282),
.B1(n_2210),
.B2(n_2198),
.Y(n_2388)
);

OAI31xp33_ASAP7_75t_L g2389 ( 
.A1(n_2374),
.A2(n_2305),
.A3(n_2300),
.B(n_2294),
.Y(n_2389)
);

NAND2xp33_ASAP7_75t_SL g2390 ( 
.A(n_2368),
.B(n_2210),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2387),
.B(n_2227),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2384),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_SL g2393 ( 
.A(n_2385),
.B(n_2306),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2382),
.Y(n_2394)
);

OAI31xp33_ASAP7_75t_SL g2395 ( 
.A1(n_2379),
.A2(n_2292),
.A3(n_2227),
.B(n_2310),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2383),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2378),
.B(n_2310),
.Y(n_2397)
);

CKINVDCx16_ASAP7_75t_R g2398 ( 
.A(n_2390),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2380),
.B(n_2311),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2388),
.B(n_2311),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2386),
.Y(n_2401)
);

NOR2x1_ASAP7_75t_L g2402 ( 
.A(n_2381),
.B(n_2210),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2389),
.B(n_2300),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2383),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2387),
.B(n_2287),
.Y(n_2405)
);

AOI22xp33_ASAP7_75t_L g2406 ( 
.A1(n_2399),
.A2(n_2292),
.B1(n_2295),
.B2(n_2215),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2393),
.B(n_2398),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2391),
.B(n_2155),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2396),
.Y(n_2409)
);

BUFx3_ASAP7_75t_L g2410 ( 
.A(n_2392),
.Y(n_2410)
);

HB1xp67_ASAP7_75t_L g2411 ( 
.A(n_2402),
.Y(n_2411)
);

INVxp67_ASAP7_75t_L g2412 ( 
.A(n_2393),
.Y(n_2412)
);

INVx1_ASAP7_75t_SL g2413 ( 
.A(n_2404),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2400),
.B(n_2311),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2401),
.B(n_2182),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2403),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2405),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2394),
.B(n_2311),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2397),
.B(n_2303),
.Y(n_2419)
);

OAI22xp5_ASAP7_75t_L g2420 ( 
.A1(n_2406),
.A2(n_2395),
.B1(n_2298),
.B2(n_2215),
.Y(n_2420)
);

OAI322xp33_ASAP7_75t_L g2421 ( 
.A1(n_2412),
.A2(n_2395),
.A3(n_111),
.B1(n_108),
.B2(n_110),
.C1(n_106),
.C2(n_107),
.Y(n_2421)
);

AOI21xp33_ASAP7_75t_L g2422 ( 
.A1(n_2407),
.A2(n_107),
.B(n_108),
.Y(n_2422)
);

NAND3xp33_ASAP7_75t_L g2423 ( 
.A(n_2411),
.B(n_109),
.C(n_110),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2413),
.B(n_2298),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2410),
.Y(n_2425)
);

NAND3xp33_ASAP7_75t_SL g2426 ( 
.A(n_2415),
.B(n_2268),
.C(n_2112),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2409),
.B(n_109),
.Y(n_2427)
);

OAI21xp5_ASAP7_75t_L g2428 ( 
.A1(n_2408),
.A2(n_2416),
.B(n_2418),
.Y(n_2428)
);

OAI32xp33_ASAP7_75t_L g2429 ( 
.A1(n_2419),
.A2(n_2298),
.A3(n_2181),
.B1(n_2280),
.B2(n_2258),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2417),
.Y(n_2430)
);

INVx2_ASAP7_75t_SL g2431 ( 
.A(n_2414),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2417),
.B(n_2295),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2413),
.B(n_2295),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2410),
.Y(n_2434)
);

OAI322xp33_ASAP7_75t_SL g2435 ( 
.A1(n_2416),
.A2(n_2252),
.A3(n_2285),
.B1(n_2271),
.B2(n_2283),
.C1(n_2277),
.C2(n_2269),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2413),
.B(n_2308),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2414),
.B(n_2289),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2409),
.Y(n_2438)
);

INVx3_ASAP7_75t_L g2439 ( 
.A(n_2410),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_L g2440 ( 
.A(n_2413),
.B(n_112),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2409),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2431),
.B(n_113),
.Y(n_2442)
);

AOI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2439),
.A2(n_2273),
.B1(n_2258),
.B2(n_2172),
.Y(n_2443)
);

OAI21xp33_ASAP7_75t_L g2444 ( 
.A1(n_2424),
.A2(n_2296),
.B(n_2253),
.Y(n_2444)
);

OR2x2_ASAP7_75t_L g2445 ( 
.A(n_2439),
.B(n_114),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2440),
.B(n_115),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2437),
.B(n_115),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2427),
.B(n_116),
.Y(n_2448)
);

AOI21xp5_ASAP7_75t_L g2449 ( 
.A1(n_2421),
.A2(n_2167),
.B(n_116),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2428),
.A2(n_117),
.B(n_118),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2425),
.B(n_117),
.Y(n_2451)
);

A2O1A1Ixp33_ASAP7_75t_L g2452 ( 
.A1(n_2423),
.A2(n_2296),
.B(n_2308),
.C(n_120),
.Y(n_2452)
);

OAI33xp33_ASAP7_75t_L g2453 ( 
.A1(n_2438),
.A2(n_120),
.A3(n_123),
.B1(n_118),
.B2(n_119),
.B3(n_122),
.Y(n_2453)
);

AOI21xp33_ASAP7_75t_SL g2454 ( 
.A1(n_2422),
.A2(n_119),
.B(n_122),
.Y(n_2454)
);

NAND3xp33_ASAP7_75t_SL g2455 ( 
.A(n_2434),
.B(n_2441),
.C(n_2430),
.Y(n_2455)
);

O2A1O1Ixp33_ASAP7_75t_L g2456 ( 
.A1(n_2433),
.A2(n_2432),
.B(n_2436),
.C(n_2429),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2420),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2426),
.Y(n_2458)
);

OAI21xp33_ASAP7_75t_L g2459 ( 
.A1(n_2435),
.A2(n_2293),
.B(n_2126),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2439),
.B(n_2289),
.Y(n_2460)
);

NAND2xp33_ASAP7_75t_SL g2461 ( 
.A(n_2439),
.B(n_2177),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2431),
.B(n_124),
.Y(n_2462)
);

AOI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_2431),
.A2(n_2293),
.B1(n_2137),
.B2(n_2177),
.Y(n_2463)
);

AOI221xp5_ASAP7_75t_L g2464 ( 
.A1(n_2421),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.C(n_128),
.Y(n_2464)
);

OAI322xp33_ASAP7_75t_L g2465 ( 
.A1(n_2424),
.A2(n_130),
.A3(n_129),
.B1(n_127),
.B2(n_125),
.C1(n_126),
.C2(n_128),
.Y(n_2465)
);

OAI321xp33_ASAP7_75t_L g2466 ( 
.A1(n_2424),
.A2(n_2144),
.A3(n_2257),
.B1(n_2130),
.B2(n_131),
.C(n_133),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2424),
.Y(n_2467)
);

AOI221x1_ASAP7_75t_L g2468 ( 
.A1(n_2440),
.A2(n_132),
.B1(n_129),
.B2(n_130),
.C(n_134),
.Y(n_2468)
);

OAI21xp5_ASAP7_75t_L g2469 ( 
.A1(n_2440),
.A2(n_2297),
.B(n_2257),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2431),
.B(n_132),
.Y(n_2470)
);

AOI211x1_ASAP7_75t_L g2471 ( 
.A1(n_2429),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2424),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2431),
.B(n_135),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2431),
.B(n_136),
.Y(n_2474)
);

AOI21xp5_ASAP7_75t_L g2475 ( 
.A1(n_2431),
.A2(n_138),
.B(n_139),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2431),
.B(n_139),
.Y(n_2476)
);

INVxp67_ASAP7_75t_L g2477 ( 
.A(n_2440),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2431),
.B(n_140),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2460),
.B(n_140),
.Y(n_2479)
);

OAI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2463),
.A2(n_2137),
.B1(n_2130),
.B2(n_2293),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2464),
.B(n_2130),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2445),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2467),
.B(n_2289),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2442),
.Y(n_2484)
);

INVx2_ASAP7_75t_SL g2485 ( 
.A(n_2478),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2462),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2475),
.B(n_141),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2468),
.B(n_141),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2449),
.B(n_142),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2472),
.B(n_2289),
.Y(n_2490)
);

OR2x2_ASAP7_75t_L g2491 ( 
.A(n_2470),
.B(n_143),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2471),
.B(n_2450),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2473),
.Y(n_2493)
);

NOR2x1_ASAP7_75t_L g2494 ( 
.A(n_2455),
.B(n_144),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2457),
.B(n_2293),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2474),
.Y(n_2496)
);

INVxp67_ASAP7_75t_L g2497 ( 
.A(n_2476),
.Y(n_2497)
);

OAI321xp33_ASAP7_75t_L g2498 ( 
.A1(n_2458),
.A2(n_146),
.A3(n_149),
.B1(n_144),
.B2(n_145),
.C(n_148),
.Y(n_2498)
);

NOR2xp33_ASAP7_75t_L g2499 ( 
.A(n_2447),
.B(n_145),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2477),
.B(n_2451),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2448),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2454),
.B(n_2284),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2446),
.B(n_146),
.Y(n_2503)
);

OR2x6_ASAP7_75t_L g2504 ( 
.A(n_2456),
.B(n_2165),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_SL g2505 ( 
.A(n_2466),
.B(n_2165),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2459),
.B(n_2297),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2443),
.B(n_148),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2461),
.B(n_149),
.Y(n_2508)
);

INVx2_ASAP7_75t_SL g2509 ( 
.A(n_2453),
.Y(n_2509)
);

AND2x4_ASAP7_75t_L g2510 ( 
.A(n_2452),
.B(n_150),
.Y(n_2510)
);

NAND2x1_ASAP7_75t_L g2511 ( 
.A(n_2469),
.B(n_2165),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2444),
.B(n_150),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2465),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2460),
.B(n_151),
.Y(n_2514)
);

INVxp67_ASAP7_75t_L g2515 ( 
.A(n_2445),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2460),
.B(n_152),
.Y(n_2516)
);

INVx2_ASAP7_75t_SL g2517 ( 
.A(n_2494),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2488),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2495),
.Y(n_2519)
);

INVx1_ASAP7_75t_SL g2520 ( 
.A(n_2491),
.Y(n_2520)
);

NOR2xp33_ASAP7_75t_L g2521 ( 
.A(n_2479),
.B(n_152),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2516),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2514),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2483),
.B(n_154),
.Y(n_2524)
);

AOI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2509),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2490),
.B(n_155),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2499),
.B(n_156),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2508),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2502),
.B(n_157),
.Y(n_2529)
);

NOR2xp33_ASAP7_75t_L g2530 ( 
.A(n_2515),
.B(n_157),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2487),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2489),
.Y(n_2532)
);

XNOR2xp5_ASAP7_75t_L g2533 ( 
.A(n_2513),
.B(n_158),
.Y(n_2533)
);

NOR2xp33_ASAP7_75t_L g2534 ( 
.A(n_2482),
.B(n_158),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2512),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2482),
.B(n_2510),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2504),
.Y(n_2537)
);

NAND2x1p5_ASAP7_75t_SL g2538 ( 
.A(n_2485),
.B(n_159),
.Y(n_2538)
);

BUFx2_ASAP7_75t_L g2539 ( 
.A(n_2504),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2492),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2503),
.Y(n_2541)
);

NOR3xp33_ASAP7_75t_L g2542 ( 
.A(n_2497),
.B(n_2486),
.C(n_2484),
.Y(n_2542)
);

OAI21xp33_ASAP7_75t_L g2543 ( 
.A1(n_2507),
.A2(n_159),
.B(n_160),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2510),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2481),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2496),
.B(n_160),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2505),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2500),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2501),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_L g2550 ( 
.A(n_2498),
.B(n_161),
.Y(n_2550)
);

NAND3xp33_ASAP7_75t_SL g2551 ( 
.A(n_2493),
.B(n_2511),
.C(n_2506),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2480),
.Y(n_2552)
);

OAI21xp5_ASAP7_75t_SL g2553 ( 
.A1(n_2495),
.A2(n_161),
.B(n_162),
.Y(n_2553)
);

INVxp67_ASAP7_75t_L g2554 ( 
.A(n_2494),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2495),
.B(n_162),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2495),
.B(n_163),
.Y(n_2556)
);

NAND2x1_ASAP7_75t_L g2557 ( 
.A(n_2494),
.B(n_163),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2488),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2488),
.Y(n_2559)
);

CKINVDCx20_ASAP7_75t_R g2560 ( 
.A(n_2509),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2488),
.Y(n_2561)
);

NAND2xp33_ASAP7_75t_L g2562 ( 
.A(n_2494),
.B(n_164),
.Y(n_2562)
);

INVx2_ASAP7_75t_SL g2563 ( 
.A(n_2494),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2495),
.B(n_165),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_2479),
.B(n_165),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_R g2566 ( 
.A(n_2488),
.B(n_166),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_2515),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2495),
.B(n_167),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_2479),
.B(n_167),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2495),
.B(n_168),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2495),
.B(n_168),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2495),
.B(n_169),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2495),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2495),
.B(n_169),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2495),
.B(n_170),
.Y(n_2575)
);

XNOR2xp5_ASAP7_75t_L g2576 ( 
.A(n_2495),
.B(n_170),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2488),
.Y(n_2577)
);

INVx3_ASAP7_75t_SL g2578 ( 
.A(n_2491),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_2515),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2495),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2555),
.B(n_171),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2576),
.Y(n_2582)
);

AOI22xp5_ASAP7_75t_L g2583 ( 
.A1(n_2560),
.A2(n_2110),
.B1(n_2104),
.B2(n_2138),
.Y(n_2583)
);

NOR3xp33_ASAP7_75t_L g2584 ( 
.A(n_2551),
.B(n_171),
.C(n_172),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2572),
.B(n_173),
.Y(n_2585)
);

AOI211xp5_ASAP7_75t_L g2586 ( 
.A1(n_2550),
.A2(n_175),
.B(n_173),
.C(n_174),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2526),
.B(n_175),
.Y(n_2587)
);

OAI211xp5_ASAP7_75t_L g2588 ( 
.A1(n_2553),
.A2(n_178),
.B(n_176),
.C(n_177),
.Y(n_2588)
);

AOI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_2567),
.A2(n_2110),
.B1(n_2138),
.B2(n_2168),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2533),
.Y(n_2590)
);

OAI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2554),
.A2(n_2171),
.B1(n_2156),
.B2(n_2147),
.Y(n_2591)
);

AOI211xp5_ASAP7_75t_L g2592 ( 
.A1(n_2562),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2525),
.B(n_2530),
.Y(n_2593)
);

NOR3x1_ASAP7_75t_L g2594 ( 
.A(n_2556),
.B(n_180),
.C(n_181),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2564),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2568),
.Y(n_2596)
);

OAI211xp5_ASAP7_75t_L g2597 ( 
.A1(n_2566),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_2597)
);

INVx1_ASAP7_75t_SL g2598 ( 
.A(n_2557),
.Y(n_2598)
);

OAI21xp5_ASAP7_75t_L g2599 ( 
.A1(n_2529),
.A2(n_182),
.B(n_183),
.Y(n_2599)
);

AOI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2536),
.A2(n_2563),
.B(n_2517),
.Y(n_2600)
);

OAI211xp5_ASAP7_75t_SL g2601 ( 
.A1(n_2547),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_2601)
);

AOI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2579),
.A2(n_2138),
.B1(n_2156),
.B2(n_2147),
.Y(n_2602)
);

AOI22xp5_ASAP7_75t_L g2603 ( 
.A1(n_2519),
.A2(n_2138),
.B1(n_2156),
.B2(n_2147),
.Y(n_2603)
);

O2A1O1Ixp33_ASAP7_75t_L g2604 ( 
.A1(n_2570),
.A2(n_2574),
.B(n_2575),
.C(n_2571),
.Y(n_2604)
);

INVxp67_ASAP7_75t_L g2605 ( 
.A(n_2534),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2525),
.B(n_184),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2521),
.B(n_186),
.Y(n_2607)
);

AOI21xp5_ASAP7_75t_L g2608 ( 
.A1(n_2527),
.A2(n_187),
.B(n_188),
.Y(n_2608)
);

AND2x2_ASAP7_75t_L g2609 ( 
.A(n_2573),
.B(n_187),
.Y(n_2609)
);

AOI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2580),
.A2(n_2082),
.B1(n_2083),
.B2(n_2079),
.Y(n_2610)
);

OA22x2_ASAP7_75t_L g2611 ( 
.A1(n_2537),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_2611)
);

AND4x1_ASAP7_75t_L g2612 ( 
.A(n_2542),
.B(n_191),
.C(n_189),
.D(n_190),
.Y(n_2612)
);

NAND3xp33_ASAP7_75t_L g2613 ( 
.A(n_2543),
.B(n_192),
.C(n_193),
.Y(n_2613)
);

NOR2xp33_ASAP7_75t_L g2614 ( 
.A(n_2543),
.B(n_193),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2546),
.Y(n_2615)
);

AOI22xp5_ASAP7_75t_L g2616 ( 
.A1(n_2548),
.A2(n_2089),
.B1(n_2098),
.B2(n_2094),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2538),
.Y(n_2617)
);

OAI211xp5_ASAP7_75t_SL g2618 ( 
.A1(n_2540),
.A2(n_196),
.B(n_194),
.C(n_195),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2549),
.A2(n_197),
.B1(n_194),
.B2(n_196),
.Y(n_2619)
);

NOR4xp25_ASAP7_75t_L g2620 ( 
.A(n_2545),
.B(n_199),
.C(n_197),
.D(n_198),
.Y(n_2620)
);

OAI21xp33_ASAP7_75t_SL g2621 ( 
.A1(n_2524),
.A2(n_198),
.B(n_199),
.Y(n_2621)
);

NOR2x1_ASAP7_75t_L g2622 ( 
.A(n_2539),
.B(n_2565),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2569),
.B(n_200),
.Y(n_2623)
);

NOR2x1_ASAP7_75t_L g2624 ( 
.A(n_2544),
.B(n_200),
.Y(n_2624)
);

OAI211xp5_ASAP7_75t_SL g2625 ( 
.A1(n_2518),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_2625)
);

AOI22xp5_ASAP7_75t_L g2626 ( 
.A1(n_2558),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_2626)
);

OAI22xp5_ASAP7_75t_L g2627 ( 
.A1(n_2559),
.A2(n_2577),
.B1(n_2561),
.B2(n_2535),
.Y(n_2627)
);

NOR3xp33_ASAP7_75t_SL g2628 ( 
.A(n_2552),
.B(n_204),
.C(n_205),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2522),
.Y(n_2629)
);

OAI21xp5_ASAP7_75t_L g2630 ( 
.A1(n_2523),
.A2(n_205),
.B(n_206),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2528),
.Y(n_2631)
);

OAI21xp33_ASAP7_75t_SL g2632 ( 
.A1(n_2520),
.A2(n_207),
.B(n_208),
.Y(n_2632)
);

INVx1_ASAP7_75t_SL g2633 ( 
.A(n_2578),
.Y(n_2633)
);

NOR2x1_ASAP7_75t_L g2634 ( 
.A(n_2531),
.B(n_208),
.Y(n_2634)
);

OA22x2_ASAP7_75t_L g2635 ( 
.A1(n_2532),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2541),
.B(n_211),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2576),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2555),
.B(n_213),
.Y(n_2638)
);

NAND3xp33_ASAP7_75t_L g2639 ( 
.A(n_2562),
.B(n_213),
.C(n_214),
.Y(n_2639)
);

AOI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_2560),
.A2(n_217),
.B1(n_214),
.B2(n_216),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2576),
.Y(n_2641)
);

NOR3xp33_ASAP7_75t_L g2642 ( 
.A(n_2551),
.B(n_216),
.C(n_218),
.Y(n_2642)
);

AO22x2_ASAP7_75t_L g2643 ( 
.A1(n_2517),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2576),
.Y(n_2644)
);

OAI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_2560),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2555),
.B(n_222),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2555),
.B(n_222),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2576),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2555),
.B(n_223),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2576),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2576),
.Y(n_2651)
);

NAND3xp33_ASAP7_75t_L g2652 ( 
.A(n_2562),
.B(n_224),
.C(n_225),
.Y(n_2652)
);

OAI22xp33_ASAP7_75t_L g2653 ( 
.A1(n_2529),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2576),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2576),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2576),
.Y(n_2656)
);

OAI21xp33_ASAP7_75t_L g2657 ( 
.A1(n_2633),
.A2(n_226),
.B(n_228),
.Y(n_2657)
);

INVxp67_ASAP7_75t_L g2658 ( 
.A(n_2649),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2624),
.Y(n_2659)
);

INVxp67_ASAP7_75t_L g2660 ( 
.A(n_2609),
.Y(n_2660)
);

AOI21xp33_ASAP7_75t_L g2661 ( 
.A1(n_2621),
.A2(n_228),
.B(n_229),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2628),
.B(n_230),
.Y(n_2662)
);

AOI21xp5_ASAP7_75t_L g2663 ( 
.A1(n_2600),
.A2(n_230),
.B(n_231),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_R g2664 ( 
.A(n_2598),
.B(n_2581),
.Y(n_2664)
);

INVxp67_ASAP7_75t_L g2665 ( 
.A(n_2634),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2611),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2612),
.B(n_231),
.Y(n_2667)
);

AOI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2584),
.A2(n_2642),
.B1(n_2614),
.B2(n_2588),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2617),
.B(n_232),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2585),
.Y(n_2670)
);

NOR2xp33_ASAP7_75t_L g2671 ( 
.A(n_2587),
.B(n_232),
.Y(n_2671)
);

OR2x2_ASAP7_75t_L g2672 ( 
.A(n_2620),
.B(n_233),
.Y(n_2672)
);

INVx2_ASAP7_75t_SL g2673 ( 
.A(n_2635),
.Y(n_2673)
);

A2O1A1Ixp33_ASAP7_75t_L g2674 ( 
.A1(n_2632),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2643),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2594),
.B(n_234),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2638),
.Y(n_2677)
);

AOI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2622),
.A2(n_514),
.B1(n_238),
.B2(n_235),
.Y(n_2678)
);

A2O1A1Ixp33_ASAP7_75t_L g2679 ( 
.A1(n_2608),
.A2(n_239),
.B(n_236),
.C(n_238),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2646),
.Y(n_2680)
);

OAI21xp5_ASAP7_75t_L g2681 ( 
.A1(n_2639),
.A2(n_236),
.B(n_239),
.Y(n_2681)
);

OAI21xp33_ASAP7_75t_L g2682 ( 
.A1(n_2590),
.A2(n_241),
.B(n_242),
.Y(n_2682)
);

OAI21xp5_ASAP7_75t_L g2683 ( 
.A1(n_2652),
.A2(n_241),
.B(n_242),
.Y(n_2683)
);

INVxp67_ASAP7_75t_L g2684 ( 
.A(n_2636),
.Y(n_2684)
);

AOI21xp5_ASAP7_75t_SL g2685 ( 
.A1(n_2645),
.A2(n_514),
.B(n_243),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2647),
.Y(n_2686)
);

AOI211xp5_ASAP7_75t_L g2687 ( 
.A1(n_2613),
.A2(n_246),
.B(n_244),
.C(n_245),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2643),
.Y(n_2688)
);

OAI221xp5_ASAP7_75t_L g2689 ( 
.A1(n_2592),
.A2(n_247),
.B1(n_244),
.B2(n_246),
.C(n_248),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2606),
.Y(n_2690)
);

NOR2x1_ASAP7_75t_L g2691 ( 
.A(n_2597),
.B(n_247),
.Y(n_2691)
);

AOI211xp5_ASAP7_75t_L g2692 ( 
.A1(n_2627),
.A2(n_2601),
.B(n_2618),
.C(n_2625),
.Y(n_2692)
);

OR2x2_ASAP7_75t_L g2693 ( 
.A(n_2607),
.B(n_249),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2623),
.Y(n_2694)
);

AOI221xp5_ASAP7_75t_L g2695 ( 
.A1(n_2586),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.C(n_252),
.Y(n_2695)
);

OAI21xp5_ASAP7_75t_SL g2696 ( 
.A1(n_2629),
.A2(n_250),
.B(n_252),
.Y(n_2696)
);

AOI21xp33_ASAP7_75t_L g2697 ( 
.A1(n_2604),
.A2(n_253),
.B(n_254),
.Y(n_2697)
);

AOI322xp5_ASAP7_75t_L g2698 ( 
.A1(n_2631),
.A2(n_253),
.A3(n_254),
.B1(n_255),
.B2(n_256),
.C1(n_257),
.C2(n_258),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2599),
.Y(n_2699)
);

AOI322xp5_ASAP7_75t_L g2700 ( 
.A1(n_2582),
.A2(n_2656),
.A3(n_2655),
.B1(n_2654),
.B2(n_2637),
.C1(n_2651),
.C2(n_2650),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_2641),
.A2(n_258),
.B1(n_255),
.B2(n_257),
.Y(n_2701)
);

OAI22xp5_ASAP7_75t_SL g2702 ( 
.A1(n_2644),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_2702)
);

NOR2x1_ASAP7_75t_L g2703 ( 
.A(n_2653),
.B(n_259),
.Y(n_2703)
);

OAI21xp33_ASAP7_75t_SL g2704 ( 
.A1(n_2603),
.A2(n_260),
.B(n_262),
.Y(n_2704)
);

XNOR2xp5_ASAP7_75t_L g2705 ( 
.A(n_2648),
.B(n_263),
.Y(n_2705)
);

OAI22xp33_ASAP7_75t_L g2706 ( 
.A1(n_2640),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_2706)
);

AOI211xp5_ASAP7_75t_L g2707 ( 
.A1(n_2593),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_2707)
);

OAI221xp5_ASAP7_75t_L g2708 ( 
.A1(n_2605),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.C(n_270),
.Y(n_2708)
);

OAI21xp5_ASAP7_75t_L g2709 ( 
.A1(n_2595),
.A2(n_2596),
.B(n_2615),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2630),
.Y(n_2710)
);

OAI22xp5_ASAP7_75t_L g2711 ( 
.A1(n_2583),
.A2(n_2602),
.B1(n_2589),
.B2(n_2626),
.Y(n_2711)
);

OAI21xp33_ASAP7_75t_L g2712 ( 
.A1(n_2591),
.A2(n_267),
.B(n_268),
.Y(n_2712)
);

OAI221xp5_ASAP7_75t_L g2713 ( 
.A1(n_2619),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.C(n_272),
.Y(n_2713)
);

OAI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2610),
.A2(n_271),
.B(n_272),
.Y(n_2714)
);

AOI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2616),
.A2(n_277),
.B1(n_273),
.B2(n_274),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2624),
.Y(n_2716)
);

OR2x2_ASAP7_75t_L g2717 ( 
.A(n_2620),
.B(n_273),
.Y(n_2717)
);

NOR4xp25_ASAP7_75t_L g2718 ( 
.A(n_2633),
.B(n_278),
.C(n_274),
.D(n_277),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2624),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2649),
.B(n_278),
.Y(n_2720)
);

A2O1A1Ixp33_ASAP7_75t_L g2721 ( 
.A1(n_2614),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_2721)
);

AOI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2661),
.A2(n_281),
.B(n_282),
.Y(n_2722)
);

AOI211xp5_ASAP7_75t_L g2723 ( 
.A1(n_2718),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_2723)
);

O2A1O1Ixp33_ASAP7_75t_L g2724 ( 
.A1(n_2665),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_2724)
);

AOI322xp5_ASAP7_75t_L g2725 ( 
.A1(n_2666),
.A2(n_285),
.A3(n_286),
.B1(n_287),
.B2(n_288),
.C1(n_289),
.C2(n_290),
.Y(n_2725)
);

NAND4xp25_ASAP7_75t_L g2726 ( 
.A(n_2692),
.B(n_291),
.C(n_286),
.D(n_289),
.Y(n_2726)
);

OAI221xp5_ASAP7_75t_SL g2727 ( 
.A1(n_2700),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.C(n_294),
.Y(n_2727)
);

NAND4xp25_ASAP7_75t_SL g2728 ( 
.A(n_2695),
.B(n_294),
.C(n_292),
.D(n_293),
.Y(n_2728)
);

AOI221x1_ASAP7_75t_L g2729 ( 
.A1(n_2663),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.C(n_298),
.Y(n_2729)
);

OAI221xp5_ASAP7_75t_L g2730 ( 
.A1(n_2712),
.A2(n_296),
.B1(n_299),
.B2(n_300),
.C(n_301),
.Y(n_2730)
);

AOI222xp33_ASAP7_75t_L g2731 ( 
.A1(n_2704),
.A2(n_2662),
.B1(n_2719),
.B2(n_2659),
.C1(n_2716),
.C2(n_2676),
.Y(n_2731)
);

AOI221x1_ASAP7_75t_L g2732 ( 
.A1(n_2675),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.C(n_302),
.Y(n_2732)
);

AOI221xp5_ASAP7_75t_L g2733 ( 
.A1(n_2685),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.C(n_306),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_SL g2734 ( 
.A(n_2706),
.B(n_303),
.Y(n_2734)
);

A2O1A1Ixp33_ASAP7_75t_L g2735 ( 
.A1(n_2697),
.A2(n_307),
.B(n_304),
.C(n_306),
.Y(n_2735)
);

AOI221xp5_ASAP7_75t_L g2736 ( 
.A1(n_2674),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.C(n_310),
.Y(n_2736)
);

NAND5xp2_ASAP7_75t_L g2737 ( 
.A(n_2668),
.B(n_308),
.C(n_309),
.D(n_310),
.E(n_311),
.Y(n_2737)
);

AOI221xp5_ASAP7_75t_L g2738 ( 
.A1(n_2673),
.A2(n_2688),
.B1(n_2711),
.B2(n_2681),
.C(n_2683),
.Y(n_2738)
);

OR2x2_ASAP7_75t_L g2739 ( 
.A(n_2672),
.B(n_311),
.Y(n_2739)
);

AOI22xp33_ASAP7_75t_L g2740 ( 
.A1(n_2691),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_2740)
);

O2A1O1Ixp5_ASAP7_75t_L g2741 ( 
.A1(n_2709),
.A2(n_315),
.B(n_313),
.C(n_314),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2720),
.Y(n_2742)
);

O2A1O1Ixp5_ASAP7_75t_L g2743 ( 
.A1(n_2717),
.A2(n_317),
.B(n_315),
.C(n_316),
.Y(n_2743)
);

AOI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2658),
.A2(n_319),
.B1(n_316),
.B2(n_318),
.Y(n_2744)
);

NAND3xp33_ASAP7_75t_SL g2745 ( 
.A(n_2687),
.B(n_2664),
.C(n_2667),
.Y(n_2745)
);

OAI21xp33_ASAP7_75t_L g2746 ( 
.A1(n_2668),
.A2(n_319),
.B(n_320),
.Y(n_2746)
);

INVx3_ASAP7_75t_L g2747 ( 
.A(n_2669),
.Y(n_2747)
);

NAND2xp33_ASAP7_75t_R g2748 ( 
.A(n_2693),
.B(n_513),
.Y(n_2748)
);

AOI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_2660),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_2749)
);

NAND3xp33_ASAP7_75t_L g2750 ( 
.A(n_2679),
.B(n_321),
.C(n_323),
.Y(n_2750)
);

NAND3x1_ASAP7_75t_L g2751 ( 
.A(n_2703),
.B(n_323),
.C(n_324),
.Y(n_2751)
);

AOI221xp5_ASAP7_75t_L g2752 ( 
.A1(n_2689),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.C(n_327),
.Y(n_2752)
);

NAND4xp75_ASAP7_75t_L g2753 ( 
.A(n_2699),
.B(n_327),
.C(n_325),
.D(n_326),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2671),
.B(n_329),
.Y(n_2754)
);

NOR2x1p5_ASAP7_75t_L g2755 ( 
.A(n_2710),
.B(n_329),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2696),
.B(n_331),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2705),
.Y(n_2757)
);

OAI221xp5_ASAP7_75t_L g2758 ( 
.A1(n_2714),
.A2(n_331),
.B1(n_332),
.B2(n_334),
.C(n_335),
.Y(n_2758)
);

AOI222xp33_ASAP7_75t_L g2759 ( 
.A1(n_2690),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.C1(n_336),
.C2(n_337),
.Y(n_2759)
);

AOI211xp5_ASAP7_75t_SL g2760 ( 
.A1(n_2684),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_2760)
);

INVx2_ASAP7_75t_SL g2761 ( 
.A(n_2670),
.Y(n_2761)
);

NAND3xp33_ASAP7_75t_L g2762 ( 
.A(n_2721),
.B(n_339),
.C(n_340),
.Y(n_2762)
);

AOI211x1_ASAP7_75t_SL g2763 ( 
.A1(n_2677),
.A2(n_341),
.B(n_339),
.C(n_340),
.Y(n_2763)
);

AOI22xp5_ASAP7_75t_L g2764 ( 
.A1(n_2680),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2702),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2657),
.B(n_342),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_SL g2767 ( 
.A(n_2715),
.B(n_343),
.Y(n_2767)
);

AOI22xp33_ASAP7_75t_L g2768 ( 
.A1(n_2686),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_2768)
);

AND4x2_ASAP7_75t_L g2769 ( 
.A(n_2713),
.B(n_349),
.C(n_347),
.D(n_348),
.Y(n_2769)
);

OAI211xp5_ASAP7_75t_SL g2770 ( 
.A1(n_2694),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2682),
.B(n_350),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2678),
.Y(n_2772)
);

OAI221xp5_ASAP7_75t_L g2773 ( 
.A1(n_2707),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.C(n_354),
.Y(n_2773)
);

AOI211xp5_ASAP7_75t_SL g2774 ( 
.A1(n_2708),
.A2(n_355),
.B(n_352),
.C(n_354),
.Y(n_2774)
);

NAND3xp33_ASAP7_75t_L g2775 ( 
.A(n_2727),
.B(n_2701),
.C(n_2698),
.Y(n_2775)
);

NAND4xp75_ASAP7_75t_L g2776 ( 
.A(n_2738),
.B(n_359),
.C(n_356),
.D(n_357),
.Y(n_2776)
);

AOI22xp5_ASAP7_75t_L g2777 ( 
.A1(n_2728),
.A2(n_2761),
.B1(n_2748),
.B2(n_2745),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2755),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2739),
.Y(n_2779)
);

NOR3xp33_ASAP7_75t_L g2780 ( 
.A(n_2747),
.B(n_513),
.C(n_357),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2769),
.Y(n_2781)
);

NOR2x1_ASAP7_75t_L g2782 ( 
.A(n_2753),
.B(n_359),
.Y(n_2782)
);

NOR2x1p5_ASAP7_75t_L g2783 ( 
.A(n_2756),
.B(n_360),
.Y(n_2783)
);

NOR3x1_ASAP7_75t_L g2784 ( 
.A(n_2730),
.B(n_512),
.C(n_361),
.Y(n_2784)
);

AO22x1_ASAP7_75t_L g2785 ( 
.A1(n_2765),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_2785)
);

INVxp67_ASAP7_75t_L g2786 ( 
.A(n_2737),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_L g2787 ( 
.A(n_2773),
.B(n_362),
.Y(n_2787)
);

NOR2x1p5_ASAP7_75t_L g2788 ( 
.A(n_2747),
.B(n_363),
.Y(n_2788)
);

NOR4xp75_ASAP7_75t_L g2789 ( 
.A(n_2751),
.B(n_364),
.C(n_365),
.D(n_366),
.Y(n_2789)
);

NOR3xp33_ASAP7_75t_L g2790 ( 
.A(n_2757),
.B(n_2754),
.C(n_2772),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2774),
.B(n_2740),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2743),
.Y(n_2792)
);

XNOR2xp5_ASAP7_75t_L g2793 ( 
.A(n_2763),
.B(n_2723),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2766),
.Y(n_2794)
);

NOR3xp33_ASAP7_75t_L g2795 ( 
.A(n_2742),
.B(n_511),
.C(n_364),
.Y(n_2795)
);

AO21x1_ASAP7_75t_L g2796 ( 
.A1(n_2722),
.A2(n_365),
.B(n_366),
.Y(n_2796)
);

NOR2x1p5_ASAP7_75t_L g2797 ( 
.A(n_2771),
.B(n_367),
.Y(n_2797)
);

NOR2x1_ASAP7_75t_SL g2798 ( 
.A(n_2750),
.B(n_2762),
.Y(n_2798)
);

NAND4xp75_ASAP7_75t_L g2799 ( 
.A(n_2729),
.B(n_367),
.C(n_369),
.D(n_370),
.Y(n_2799)
);

NOR3xp33_ASAP7_75t_SL g2800 ( 
.A(n_2734),
.B(n_370),
.C(n_371),
.Y(n_2800)
);

OAI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2758),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_2801)
);

INVxp67_ASAP7_75t_L g2802 ( 
.A(n_2726),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2746),
.B(n_373),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2741),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2764),
.Y(n_2805)
);

NAND3xp33_ASAP7_75t_SL g2806 ( 
.A(n_2731),
.B(n_375),
.C(n_376),
.Y(n_2806)
);

NOR2x1_ASAP7_75t_L g2807 ( 
.A(n_2770),
.B(n_375),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_SL g2808 ( 
.A(n_2733),
.B(n_377),
.Y(n_2808)
);

NOR3xp33_ASAP7_75t_L g2809 ( 
.A(n_2752),
.B(n_510),
.C(n_378),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2767),
.B(n_378),
.Y(n_2810)
);

NOR3xp33_ASAP7_75t_L g2811 ( 
.A(n_2736),
.B(n_379),
.C(n_380),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2735),
.Y(n_2812)
);

NAND4xp75_ASAP7_75t_L g2813 ( 
.A(n_2732),
.B(n_380),
.C(n_381),
.D(n_382),
.Y(n_2813)
);

NOR3xp33_ASAP7_75t_L g2814 ( 
.A(n_2724),
.B(n_2749),
.C(n_2744),
.Y(n_2814)
);

NOR2x1_ASAP7_75t_L g2815 ( 
.A(n_2760),
.B(n_382),
.Y(n_2815)
);

INVxp67_ASAP7_75t_SL g2816 ( 
.A(n_2759),
.Y(n_2816)
);

AOI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2808),
.A2(n_2768),
.B(n_2725),
.Y(n_2817)
);

AOI221xp5_ASAP7_75t_L g2818 ( 
.A1(n_2806),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.C(n_387),
.Y(n_2818)
);

NOR4xp25_ASAP7_75t_L g2819 ( 
.A(n_2781),
.B(n_383),
.C(n_384),
.D(n_385),
.Y(n_2819)
);

NAND3xp33_ASAP7_75t_L g2820 ( 
.A(n_2790),
.B(n_388),
.C(n_389),
.Y(n_2820)
);

AOI221xp5_ASAP7_75t_L g2821 ( 
.A1(n_2801),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.C(n_392),
.Y(n_2821)
);

NAND4xp75_ASAP7_75t_L g2822 ( 
.A(n_2782),
.B(n_390),
.C(n_391),
.D(n_392),
.Y(n_2822)
);

INVxp67_ASAP7_75t_SL g2823 ( 
.A(n_2788),
.Y(n_2823)
);

AOI211x1_ASAP7_75t_SL g2824 ( 
.A1(n_2775),
.A2(n_2805),
.B(n_2803),
.C(n_2793),
.Y(n_2824)
);

AOI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2816),
.A2(n_393),
.B(n_394),
.Y(n_2825)
);

NOR2x1_ASAP7_75t_L g2826 ( 
.A(n_2813),
.B(n_394),
.Y(n_2826)
);

NOR2xp67_ASAP7_75t_L g2827 ( 
.A(n_2786),
.B(n_395),
.Y(n_2827)
);

OAI221xp5_ASAP7_75t_L g2828 ( 
.A1(n_2777),
.A2(n_2811),
.B1(n_2809),
.B2(n_2800),
.C(n_2815),
.Y(n_2828)
);

AOI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2804),
.A2(n_395),
.B(n_396),
.Y(n_2829)
);

AOI22xp5_ASAP7_75t_L g2830 ( 
.A1(n_2810),
.A2(n_396),
.B1(n_397),
.B2(n_399),
.Y(n_2830)
);

NAND3xp33_ASAP7_75t_SL g2831 ( 
.A(n_2789),
.B(n_397),
.C(n_399),
.Y(n_2831)
);

NOR3xp33_ASAP7_75t_L g2832 ( 
.A(n_2792),
.B(n_400),
.C(n_401),
.Y(n_2832)
);

BUFx4f_ASAP7_75t_SL g2833 ( 
.A(n_2779),
.Y(n_2833)
);

NOR3xp33_ASAP7_75t_SL g2834 ( 
.A(n_2778),
.B(n_400),
.C(n_401),
.Y(n_2834)
);

NAND4xp25_ASAP7_75t_L g2835 ( 
.A(n_2784),
.B(n_402),
.C(n_404),
.D(n_405),
.Y(n_2835)
);

NOR3xp33_ASAP7_75t_L g2836 ( 
.A(n_2812),
.B(n_402),
.C(n_405),
.Y(n_2836)
);

NOR3xp33_ASAP7_75t_L g2837 ( 
.A(n_2802),
.B(n_406),
.C(n_407),
.Y(n_2837)
);

NOR2xp33_ASAP7_75t_L g2838 ( 
.A(n_2796),
.B(n_407),
.Y(n_2838)
);

NOR3xp33_ASAP7_75t_SL g2839 ( 
.A(n_2799),
.B(n_408),
.C(n_409),
.Y(n_2839)
);

NOR3xp33_ASAP7_75t_L g2840 ( 
.A(n_2794),
.B(n_2787),
.C(n_2791),
.Y(n_2840)
);

NOR2x1_ASAP7_75t_L g2841 ( 
.A(n_2776),
.B(n_2783),
.Y(n_2841)
);

AOI211x1_ASAP7_75t_SL g2842 ( 
.A1(n_2807),
.A2(n_408),
.B(n_409),
.C(n_410),
.Y(n_2842)
);

NAND4xp75_ASAP7_75t_L g2843 ( 
.A(n_2826),
.B(n_2841),
.C(n_2825),
.D(n_2827),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2822),
.Y(n_2844)
);

AOI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2831),
.A2(n_2814),
.B1(n_2797),
.B2(n_2780),
.Y(n_2845)
);

NAND4xp75_ASAP7_75t_L g2846 ( 
.A(n_2838),
.B(n_2798),
.C(n_2785),
.D(n_2795),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2834),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2842),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2839),
.B(n_2823),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2833),
.Y(n_2850)
);

NOR2x1_ASAP7_75t_L g2851 ( 
.A(n_2820),
.B(n_411),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2835),
.Y(n_2852)
);

NOR2x1p5_ASAP7_75t_L g2853 ( 
.A(n_2824),
.B(n_412),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2832),
.Y(n_2854)
);

AO22x2_ASAP7_75t_L g2855 ( 
.A1(n_2840),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_2855)
);

AND2x2_ASAP7_75t_SL g2856 ( 
.A(n_2818),
.B(n_2819),
.Y(n_2856)
);

INVxp67_ASAP7_75t_L g2857 ( 
.A(n_2829),
.Y(n_2857)
);

NAND2x1p5_ASAP7_75t_L g2858 ( 
.A(n_2830),
.B(n_413),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2836),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2828),
.Y(n_2860)
);

OR2x2_ASAP7_75t_L g2861 ( 
.A(n_2837),
.B(n_414),
.Y(n_2861)
);

NOR2x1_ASAP7_75t_L g2862 ( 
.A(n_2817),
.B(n_416),
.Y(n_2862)
);

NAND4xp75_ASAP7_75t_L g2863 ( 
.A(n_2821),
.B(n_416),
.C(n_417),
.D(n_418),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2833),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2822),
.Y(n_2865)
);

AND2x4_ASAP7_75t_L g2866 ( 
.A(n_2841),
.B(n_419),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2822),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2822),
.Y(n_2868)
);

INVx2_ASAP7_75t_SL g2869 ( 
.A(n_2826),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2822),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2822),
.Y(n_2871)
);

AND3x4_ASAP7_75t_L g2872 ( 
.A(n_2839),
.B(n_420),
.C(n_421),
.Y(n_2872)
);

NAND4xp75_ASAP7_75t_L g2873 ( 
.A(n_2826),
.B(n_420),
.C(n_421),
.D(n_422),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2822),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2822),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2822),
.Y(n_2876)
);

NOR2xp67_ASAP7_75t_SL g2877 ( 
.A(n_2843),
.B(n_2869),
.Y(n_2877)
);

AND2x4_ASAP7_75t_L g2878 ( 
.A(n_2844),
.B(n_422),
.Y(n_2878)
);

NAND2x1p5_ASAP7_75t_L g2879 ( 
.A(n_2862),
.B(n_423),
.Y(n_2879)
);

AND2x4_ASAP7_75t_L g2880 ( 
.A(n_2865),
.B(n_423),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2873),
.B(n_425),
.Y(n_2881)
);

OAI211xp5_ASAP7_75t_L g2882 ( 
.A1(n_2845),
.A2(n_426),
.B(n_427),
.C(n_428),
.Y(n_2882)
);

AOI211xp5_ASAP7_75t_L g2883 ( 
.A1(n_2861),
.A2(n_426),
.B(n_428),
.C(n_429),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2872),
.Y(n_2884)
);

NAND3xp33_ASAP7_75t_SL g2885 ( 
.A(n_2850),
.B(n_2868),
.C(n_2867),
.Y(n_2885)
);

AND2x4_ASAP7_75t_L g2886 ( 
.A(n_2870),
.B(n_429),
.Y(n_2886)
);

OR3x1_ASAP7_75t_L g2887 ( 
.A(n_2848),
.B(n_430),
.C(n_432),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2855),
.Y(n_2888)
);

AND4x1_ASAP7_75t_L g2889 ( 
.A(n_2849),
.B(n_430),
.C(n_432),
.D(n_433),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2856),
.B(n_433),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2853),
.B(n_434),
.Y(n_2891)
);

AND2x4_ASAP7_75t_L g2892 ( 
.A(n_2871),
.B(n_436),
.Y(n_2892)
);

NAND5xp2_ASAP7_75t_L g2893 ( 
.A(n_2858),
.B(n_436),
.C(n_437),
.D(n_438),
.E(n_439),
.Y(n_2893)
);

NOR2x1p5_ASAP7_75t_L g2894 ( 
.A(n_2846),
.B(n_439),
.Y(n_2894)
);

NOR3xp33_ASAP7_75t_L g2895 ( 
.A(n_2860),
.B(n_2857),
.C(n_2874),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2887),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2894),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2891),
.B(n_2866),
.Y(n_2898)
);

NAND5xp2_ASAP7_75t_L g2899 ( 
.A(n_2895),
.B(n_2879),
.C(n_2847),
.D(n_2875),
.E(n_2876),
.Y(n_2899)
);

NAND3xp33_ASAP7_75t_SL g2900 ( 
.A(n_2881),
.B(n_2852),
.C(n_2854),
.Y(n_2900)
);

AOI22xp33_ASAP7_75t_L g2901 ( 
.A1(n_2877),
.A2(n_2851),
.B1(n_2859),
.B2(n_2855),
.Y(n_2901)
);

NOR2x1_ASAP7_75t_L g2902 ( 
.A(n_2888),
.B(n_2863),
.Y(n_2902)
);

NOR2x1p5_ASAP7_75t_L g2903 ( 
.A(n_2885),
.B(n_2864),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2890),
.Y(n_2904)
);

AOI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2884),
.A2(n_440),
.B(n_441),
.Y(n_2905)
);

OR3x2_ASAP7_75t_L g2906 ( 
.A(n_2893),
.B(n_440),
.C(n_441),
.Y(n_2906)
);

NOR2x1_ASAP7_75t_L g2907 ( 
.A(n_2882),
.B(n_442),
.Y(n_2907)
);

NAND2x1p5_ASAP7_75t_L g2908 ( 
.A(n_2889),
.B(n_442),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_SL g2909 ( 
.A(n_2883),
.B(n_443),
.Y(n_2909)
);

OAI21xp33_ASAP7_75t_L g2910 ( 
.A1(n_2878),
.A2(n_443),
.B(n_444),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2908),
.Y(n_2911)
);

AOI22xp5_ASAP7_75t_L g2912 ( 
.A1(n_2906),
.A2(n_2892),
.B1(n_2886),
.B2(n_2880),
.Y(n_2912)
);

OAI221xp5_ASAP7_75t_L g2913 ( 
.A1(n_2901),
.A2(n_444),
.B1(n_445),
.B2(n_446),
.C(n_447),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2910),
.B(n_446),
.Y(n_2914)
);

HB1xp67_ASAP7_75t_L g2915 ( 
.A(n_2907),
.Y(n_2915)
);

OAI322xp33_ASAP7_75t_L g2916 ( 
.A1(n_2909),
.A2(n_447),
.A3(n_448),
.B1(n_449),
.B2(n_450),
.C1(n_451),
.C2(n_452),
.Y(n_2916)
);

AOI22xp33_ASAP7_75t_L g2917 ( 
.A1(n_2903),
.A2(n_451),
.B1(n_452),
.B2(n_453),
.Y(n_2917)
);

OA22x2_ASAP7_75t_L g2918 ( 
.A1(n_2896),
.A2(n_454),
.B1(n_455),
.B2(n_456),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2914),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2912),
.B(n_2902),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2918),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2915),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2911),
.Y(n_2923)
);

AO21x1_ASAP7_75t_L g2924 ( 
.A1(n_2922),
.A2(n_2898),
.B(n_2904),
.Y(n_2924)
);

OAI22xp5_ASAP7_75t_L g2925 ( 
.A1(n_2923),
.A2(n_2897),
.B1(n_2913),
.B2(n_2905),
.Y(n_2925)
);

OAI22x1_ASAP7_75t_L g2926 ( 
.A1(n_2921),
.A2(n_2899),
.B1(n_2900),
.B2(n_2916),
.Y(n_2926)
);

OAI22xp5_ASAP7_75t_L g2927 ( 
.A1(n_2920),
.A2(n_2917),
.B1(n_456),
.B2(n_457),
.Y(n_2927)
);

HB1xp67_ASAP7_75t_L g2928 ( 
.A(n_2919),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2927),
.B(n_454),
.Y(n_2929)
);

AOI21xp33_ASAP7_75t_SL g2930 ( 
.A1(n_2926),
.A2(n_457),
.B(n_458),
.Y(n_2930)
);

NAND4xp75_ASAP7_75t_L g2931 ( 
.A(n_2924),
.B(n_458),
.C(n_459),
.D(n_460),
.Y(n_2931)
);

OAI222xp33_ASAP7_75t_L g2932 ( 
.A1(n_2925),
.A2(n_459),
.B1(n_460),
.B2(n_461),
.C1(n_462),
.C2(n_463),
.Y(n_2932)
);

NOR3xp33_ASAP7_75t_SL g2933 ( 
.A(n_2928),
.B(n_461),
.C(n_462),
.Y(n_2933)
);

OAI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2927),
.A2(n_463),
.B1(n_465),
.B2(n_466),
.Y(n_2934)
);

AOI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_2934),
.A2(n_465),
.B1(n_467),
.B2(n_468),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2929),
.Y(n_2936)
);

AOI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2930),
.A2(n_468),
.B1(n_469),
.B2(n_470),
.Y(n_2937)
);

NAND3xp33_ASAP7_75t_L g2938 ( 
.A(n_2936),
.B(n_2933),
.C(n_2931),
.Y(n_2938)
);

NOR3xp33_ASAP7_75t_L g2939 ( 
.A(n_2935),
.B(n_2932),
.C(n_470),
.Y(n_2939)
);

OAI22xp5_ASAP7_75t_L g2940 ( 
.A1(n_2937),
.A2(n_469),
.B1(n_471),
.B2(n_472),
.Y(n_2940)
);

OAI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2938),
.A2(n_473),
.B1(n_474),
.B2(n_475),
.Y(n_2941)
);

OAI21x1_ASAP7_75t_L g2942 ( 
.A1(n_2940),
.A2(n_473),
.B(n_474),
.Y(n_2942)
);

OR2x6_ASAP7_75t_L g2943 ( 
.A(n_2942),
.B(n_2939),
.Y(n_2943)
);

OAI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2943),
.A2(n_2941),
.B(n_476),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_SL g2945 ( 
.A(n_2943),
.B(n_475),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2943),
.B(n_477),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2944),
.B(n_478),
.Y(n_2947)
);

AOI221xp5_ASAP7_75t_L g2948 ( 
.A1(n_2945),
.A2(n_510),
.B1(n_479),
.B2(n_480),
.C(n_481),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2947),
.Y(n_2949)
);

AOI22x1_ASAP7_75t_L g2950 ( 
.A1(n_2949),
.A2(n_2948),
.B1(n_2946),
.B2(n_480),
.Y(n_2950)
);

AOI221xp5_ASAP7_75t_L g2951 ( 
.A1(n_2950),
.A2(n_478),
.B1(n_479),
.B2(n_481),
.C(n_482),
.Y(n_2951)
);

AOI22xp33_ASAP7_75t_L g2952 ( 
.A1(n_2951),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_2952)
);

AOI211xp5_ASAP7_75t_L g2953 ( 
.A1(n_2952),
.A2(n_483),
.B(n_485),
.C(n_486),
.Y(n_2953)
);


endmodule