module real_jpeg_31074_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_578;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_611;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_634;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_0),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_0),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_0),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_0),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_1),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_1),
.A2(n_142),
.B1(n_190),
.B2(n_382),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_1),
.A2(n_190),
.B1(n_284),
.B2(n_465),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_1),
.A2(n_190),
.B1(n_533),
.B2(n_535),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_2),
.A2(n_171),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_2),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_2),
.A2(n_175),
.B1(n_244),
.B2(n_249),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_2),
.A2(n_175),
.B1(n_382),
.B2(n_387),
.Y(n_381)
);

OAI22x1_ASAP7_75t_SL g435 ( 
.A1(n_2),
.A2(n_175),
.B1(n_436),
.B2(n_438),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_4),
.A2(n_142),
.B1(n_146),
.B2(n_149),
.Y(n_141)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_4),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_4),
.A2(n_149),
.B1(n_227),
.B2(n_231),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_4),
.A2(n_149),
.B1(n_302),
.B2(n_306),
.Y(n_301)
);

AO22x1_ASAP7_75t_L g414 ( 
.A1(n_4),
.A2(n_149),
.B1(n_415),
.B2(n_419),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_5),
.A2(n_30),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_5),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_5),
.A2(n_67),
.B1(n_99),
.B2(n_104),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_5),
.A2(n_67),
.B1(n_217),
.B2(n_221),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_5),
.A2(n_67),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_6),
.A2(n_356),
.B1(n_359),
.B2(n_360),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_6),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_6),
.A2(n_359),
.B1(n_427),
.B2(n_429),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_6),
.A2(n_359),
.B1(n_549),
.B2(n_551),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_6),
.A2(n_359),
.B1(n_578),
.B2(n_579),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_7),
.A2(n_21),
.B(n_24),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_8),
.A2(n_371),
.B1(n_375),
.B2(n_376),
.Y(n_370)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_8),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_8),
.A2(n_375),
.B1(n_456),
.B2(n_459),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_8),
.A2(n_375),
.B1(n_566),
.B2(n_568),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_8),
.A2(n_375),
.B1(n_383),
.B2(n_617),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_9),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_9),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_9),
.A2(n_196),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_9),
.A2(n_196),
.B1(n_207),
.B2(n_518),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_9),
.A2(n_196),
.B1(n_601),
.B2(n_603),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_10),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_12),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_13),
.A2(n_349),
.B(n_351),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_13),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_13),
.Y(n_447)
);

OAI32xp33_ASAP7_75t_L g521 ( 
.A1(n_13),
.A2(n_184),
.A3(n_522),
.B1(n_525),
.B2(n_528),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_13),
.A2(n_90),
.B1(n_548),
.B2(n_554),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_13),
.B(n_159),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_13),
.A2(n_447),
.B1(n_630),
.B2(n_631),
.Y(n_629)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_14),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_14),
.Y(n_118)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_14),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_15),
.B(n_652),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_16),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_16),
.A2(n_81),
.B(n_85),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_16),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_16),
.A2(n_36),
.B1(n_206),
.B2(n_211),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_16),
.A2(n_36),
.B1(n_282),
.B2(n_284),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_17),
.A2(n_129),
.B1(n_133),
.B2(n_138),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_17),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_17),
.A2(n_138),
.B1(n_153),
.B2(n_156),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g269 ( 
.A1(n_17),
.A2(n_138),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_17),
.A2(n_105),
.B1(n_138),
.B2(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_18),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_18),
.Y(n_132)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_18),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_18),
.Y(n_145)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_19),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_19),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_71),
.B(n_651),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_68),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_27),
.B(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_27),
.B(n_334),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_27),
.B(n_68),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_37),
.B1(n_62),
.B2(n_63),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_28),
.A2(n_38),
.B1(n_62),
.B2(n_301),
.Y(n_329)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_32),
.Y(n_195)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_32),
.Y(n_200)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_32),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_32),
.Y(n_458)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_38),
.A2(n_62),
.B1(n_187),
.B2(n_192),
.Y(n_186)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_38),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_38),
.A2(n_62),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g347 ( 
.A1(n_38),
.A2(n_62),
.B1(n_348),
.B2(n_355),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_38),
.A2(n_62),
.B1(n_192),
.B2(n_455),
.Y(n_484)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_39),
.B(n_188),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_53),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_43),
.Y(n_305)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_43),
.Y(n_310)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_43),
.Y(n_461)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_46),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_46),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_48),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_48),
.Y(n_271)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_48),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22x1_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_56),
.B(n_182),
.Y(n_184)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_57),
.Y(n_158)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_57),
.Y(n_178)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_57),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_58),
.Y(n_374)
);

BUFx5_ASAP7_75t_L g379 ( 
.A(n_58),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_58),
.Y(n_406)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_60),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_61),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_61),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_61),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_61),
.Y(n_524)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_62),
.B(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_62),
.B(n_447),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_69),
.B(n_70),
.Y(n_68)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_66),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_70),
.A2(n_243),
.B(n_255),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_SL g268 ( 
.A(n_70),
.B(n_269),
.Y(n_268)
);

AOI22x1_ASAP7_75t_L g452 ( 
.A1(n_70),
.A2(n_275),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_336),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_333),
.B(n_335),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_320),
.B(n_332),
.Y(n_73)
);

AOI21x1_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_289),
.B(n_319),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_260),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_76),
.B(n_260),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_201),
.C(n_234),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_77),
.B(n_501),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_150),
.C(n_186),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_78),
.B(n_497),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_108),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_79),
.B(n_108),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_90),
.B(n_94),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_80),
.A2(n_474),
.B(n_476),
.Y(n_473)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_83),
.Y(n_441)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_84),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_84),
.Y(n_603)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_87),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_89),
.Y(n_413)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_89),
.Y(n_421)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_89),
.Y(n_538)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_90),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_90),
.A2(n_548),
.B1(n_565),
.B2(n_571),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_90),
.A2(n_600),
.B1(n_609),
.B2(n_611),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_92),
.Y(n_475)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_92),
.Y(n_557)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_93),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_95),
.A2(n_98),
.B(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_95),
.A2(n_239),
.B1(n_409),
.B2(n_414),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_95),
.A2(n_239),
.B1(n_598),
.B2(n_599),
.Y(n_597)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_101),
.Y(n_570)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_101),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_102),
.Y(n_437)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_102),
.Y(n_553)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_103),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_103),
.Y(n_562)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_128),
.B1(n_139),
.B2(n_141),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_109),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_109),
.A2(n_139),
.B1(n_141),
.B2(n_205),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_SL g277 ( 
.A1(n_109),
.A2(n_139),
.B(n_216),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_109),
.A2(n_139),
.B(n_216),
.Y(n_296)
);

OA22x2_ASAP7_75t_L g380 ( 
.A1(n_109),
.A2(n_139),
.B1(n_381),
.B2(n_388),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_109),
.A2(n_128),
.B1(n_139),
.B2(n_381),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_109),
.A2(n_139),
.B1(n_388),
.B2(n_516),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_109),
.A2(n_139),
.B1(n_615),
.B2(n_616),
.Y(n_614)
);

AO21x2_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_115),
.B(n_121),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_110),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_111),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_120),
.Y(n_529)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_124),
.Y(n_592)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_132),
.Y(n_618)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_137),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_139),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_139),
.B(n_447),
.Y(n_572)
);

BUFx4f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_144),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_145),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_145),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_151),
.B(n_186),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_159),
.B1(n_169),
.B2(n_179),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_152),
.A2(n_159),
.B1(n_179),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_159),
.A2(n_179),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_160),
.Y(n_288)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_170),
.A2(n_279),
.B1(n_287),
.B2(n_464),
.Y(n_485)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_173),
.Y(n_428)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_178),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_184),
.B(n_185),
.Y(n_179)
);

AO21x2_ASAP7_75t_L g279 ( 
.A1(n_180),
.A2(n_184),
.B(n_185),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_202),
.B(n_235),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_225),
.B(n_233),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_225),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_214),
.B1(n_215),
.B2(n_224),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_SL g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AO22x1_ASAP7_75t_SL g576 ( 
.A1(n_214),
.A2(n_224),
.B1(n_577),
.B2(n_582),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_214),
.A2(n_224),
.B1(n_517),
.B2(n_635),
.Y(n_634)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_220),
.Y(n_578)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_220),
.Y(n_585)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_223),
.Y(n_519)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_226),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVxp33_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_495),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_237),
.Y(n_495)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_242),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_239),
.A2(n_409),
.B1(n_435),
.B2(n_442),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_239),
.B(n_414),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_239),
.A2(n_435),
.B1(n_532),
.B2(n_539),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_257),
.B2(n_259),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_252),
.Y(n_399)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_254),
.Y(n_350)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_265),
.C(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_276),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_278),
.C(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_267),
.B(n_294),
.C(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_274),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

OAI22x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_287),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_279),
.A2(n_281),
.B1(n_287),
.B2(n_313),
.Y(n_312)
);

OA22x2_ASAP7_75t_L g363 ( 
.A1(n_279),
.A2(n_364),
.B1(n_369),
.B2(n_370),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_279),
.A2(n_369),
.B1(n_370),
.B2(n_426),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_279),
.A2(n_364),
.B1(n_369),
.B2(n_464),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_279),
.A2(n_287),
.B1(n_426),
.B2(n_629),
.Y(n_628)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_282),
.Y(n_368)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_284),
.Y(n_630)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g393 ( 
.A(n_286),
.Y(n_393)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_288),
.Y(n_369)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_292),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_297),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_298),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_311),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_312),
.C(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_313),
.Y(n_328)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

NOR2x1_ASAP7_75t_R g320 ( 
.A(n_321),
.B(n_330),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g332 ( 
.A(n_321),
.B(n_330),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_327),
.C(n_329),
.Y(n_334)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_333),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_342),
.Y(n_336)
);

NOR3xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.C(n_341),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_507),
.B(n_646),
.Y(n_342)
);

NAND4xp25_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_479),
.C(n_498),
.D(n_502),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_448),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_345),
.B(n_448),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_389),
.C(n_424),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_346),
.B(n_510),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_362),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_347),
.B(n_363),
.C(n_380),
.Y(n_477)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_350),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_350),
.Y(n_361)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_351),
.Y(n_407)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_380),
.Y(n_362)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx2_ASAP7_75t_SL g371 ( 
.A(n_372),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_373),
.Y(n_467)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_389),
.B(n_424),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_408),
.B1(n_422),
.B2(n_423),
.Y(n_389)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_390),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_390),
.B(n_423),
.Y(n_468)
);

OAI32xp33_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_394),
.A3(n_397),
.B1(n_400),
.B2(n_407),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_406),
.Y(n_633)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_408),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_421),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_433),
.C(n_446),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_425),
.B(n_513),
.Y(n_512)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_433),
.A2(n_434),
.B1(n_446),
.B2(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_446),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_447),
.B(n_529),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_447),
.B(n_554),
.Y(n_559)
);

OAI21xp33_ASAP7_75t_SL g582 ( 
.A1(n_447),
.A2(n_525),
.B(n_583),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_447),
.B(n_584),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_469),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_449),
.B(n_470),
.C(n_477),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_468),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_462),
.B2(n_463),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_462),
.C(n_468),
.Y(n_486)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_471),
.B1(n_477),
.B2(n_478),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_473),
.Y(n_482)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_477),
.Y(n_478)
);

A2O1A1O1Ixp25_ASAP7_75t_L g646 ( 
.A1(n_479),
.A2(n_498),
.B(n_647),
.C(n_649),
.D(n_650),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_488),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_480),
.B(n_488),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_486),
.C(n_487),
.Y(n_480)
);

XNOR2x1_ASAP7_75t_L g504 ( 
.A(n_481),
.B(n_505),
.Y(n_504)
);

XNOR2x1_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_482),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

INVxp33_ASAP7_75t_L g491 ( 
.A(n_484),
.Y(n_491)
);

INVxp33_ASAP7_75t_SL g492 ( 
.A(n_485),
.Y(n_492)
);

XNOR2x1_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_487),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_493),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_494),
.C(n_496),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.C(n_492),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_496),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_499),
.B(n_500),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_506),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_503),
.B(n_506),
.C(n_648),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_541),
.B(n_645),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_509),
.B(n_511),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_SL g645 ( 
.A(n_509),
.B(n_511),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_515),
.C(n_520),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g642 ( 
.A(n_512),
.B(n_643),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_515),
.B(n_520),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_530),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_521),
.A2(n_530),
.B1(n_531),
.B2(n_626),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_521),
.Y(n_626)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_532),
.Y(n_611)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

BUFx4f_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_542),
.A2(n_640),
.B(n_644),
.Y(n_541)
);

OAI31xp67_ASAP7_75t_L g542 ( 
.A1(n_543),
.A2(n_621),
.A3(n_638),
.B(n_639),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_544),
.A2(n_604),
.B(n_605),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_574),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_546),
.A2(n_563),
.B(n_573),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_547),
.B(n_558),
.Y(n_546)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx3_ASAP7_75t_SL g554 ( 
.A(n_555),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_556),
.Y(n_571)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_559),
.B(n_560),
.Y(n_558)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_562),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_572),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_564),
.B(n_572),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_565),
.Y(n_598)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_575),
.B(n_597),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_575),
.B(n_597),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_586),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_R g606 ( 
.A(n_576),
.B(n_586),
.Y(n_606)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_577),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_583),
.Y(n_593)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

AO22x1_ASAP7_75t_L g586 ( 
.A1(n_587),
.A2(n_593),
.B1(n_594),
.B2(n_596),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_SL g587 ( 
.A(n_588),
.B(n_590),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_606),
.B(n_607),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_606),
.B(n_607),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_608),
.B(n_612),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_608),
.B(n_619),
.C(n_623),
.Y(n_622)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_613),
.A2(n_614),
.B1(n_619),
.B2(n_620),
.Y(n_612)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_613),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_614),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_614),
.Y(n_623)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_616),
.Y(n_635)
);

INVx3_ASAP7_75t_SL g617 ( 
.A(n_618),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g621 ( 
.A(n_622),
.B(n_624),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_622),
.B(n_624),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_625),
.B(n_627),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_625),
.B(n_634),
.C(n_637),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_628),
.A2(n_634),
.B1(n_636),
.B2(n_637),
.Y(n_627)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_628),
.Y(n_637)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_634),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_L g640 ( 
.A(n_641),
.B(n_642),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_641),
.B(n_642),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_653),
.Y(n_652)
);


endmodule