module fake_ariane_3097_n_1483 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_49, n_20, n_283, n_50, n_187, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_251, n_116, n_39, n_155, n_127, n_1483);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1483;

wire n_913;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1432;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_967;
wire n_437;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_321;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1374;
wire n_1451;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_62),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_271),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_157),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_92),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_162),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_227),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_17),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_175),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_231),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_111),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_206),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_144),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_17),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_247),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_289),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_301),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_47),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_230),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_244),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_0),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_222),
.Y(n_339)
);

BUFx8_ASAP7_75t_SL g340 ( 
.A(n_40),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_98),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_304),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_243),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_199),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_114),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_193),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_53),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_182),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_239),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_63),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_9),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_268),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_57),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_249),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_32),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_172),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_45),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_307),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_233),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_87),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_276),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_260),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_35),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_94),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_171),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_81),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_38),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_133),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_68),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_12),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_278),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_55),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_134),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_168),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_190),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_286),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_136),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_43),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_254),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_209),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_77),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_131),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_53),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_218),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_163),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_170),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_149),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_143),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_99),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_270),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_265),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_140),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_228),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_28),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_1),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_223),
.Y(n_396)
);

BUFx5_ASAP7_75t_L g397 ( 
.A(n_89),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_177),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_267),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_314),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_145),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_298),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_236),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_291),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_108),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_27),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_303),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_160),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_202),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_189),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_152),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_255),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_141),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_96),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_128),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_155),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_232),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_185),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_253),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_285),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_186),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_203),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_115),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_40),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_138),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_122),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_293),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_237),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_12),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_312),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_56),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_112),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_14),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_225),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_272),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_3),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_302),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_238),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_80),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_224),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_205),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_61),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_44),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_72),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_113),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_28),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_273),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_33),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_97),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_288),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_287),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_33),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_79),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_24),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_250),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_315),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_76),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_251),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_116),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_86),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_48),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_216),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_119),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_217),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_73),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_248),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_308),
.Y(n_467)
);

BUFx2_ASAP7_75t_SL g468 ( 
.A(n_174),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_198),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_279),
.Y(n_470)
);

BUFx8_ASAP7_75t_SL g471 ( 
.A(n_69),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_283),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_256),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_226),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_38),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_37),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_32),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_212),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_15),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_313),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_88),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_246),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_180),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_290),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_169),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_29),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_24),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_297),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_16),
.Y(n_489)
);

BUFx5_ASAP7_75t_L g490 ( 
.A(n_183),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_240),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_280),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_252),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_148),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_196),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_60),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_213),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_21),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_153),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_49),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_204),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_221),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_85),
.Y(n_503)
);

BUFx10_ASAP7_75t_L g504 ( 
.A(n_215),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_95),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_261),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_176),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_48),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_46),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_263),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_292),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_127),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_309),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_284),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_10),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_19),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_306),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_78),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_50),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_241),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_74),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_27),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_229),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_135),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_156),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_275),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_15),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_158),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_269),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_47),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_117),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_173),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_7),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_310),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_62),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_120),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_340),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_433),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_471),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_433),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_516),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_448),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_372),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_349),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_372),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_516),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_350),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_351),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_383),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_479),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_479),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_431),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_358),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_323),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_366),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_475),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_479),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_439),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_458),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_479),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_493),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_532),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_492),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_360),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_477),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_486),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_378),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_487),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_316),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_522),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_527),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_420),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_322),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_378),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_330),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_420),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_500),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_455),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_455),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_335),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_338),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_533),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_347),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_500),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_353),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_478),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_395),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_478),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_504),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_395),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_429),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_331),
.B(n_0),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_355),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_504),
.Y(n_594)
);

INVxp33_ASAP7_75t_SL g595 ( 
.A(n_357),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_323),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_429),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_363),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_500),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_427),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g601 ( 
.A(n_500),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_364),
.Y(n_602)
);

NOR2xp67_ASAP7_75t_L g603 ( 
.A(n_367),
.B(n_1),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_427),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_513),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_370),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_394),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_384),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_474),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_466),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_406),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_424),
.Y(n_612)
);

INVxp33_ASAP7_75t_SL g613 ( 
.A(n_436),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_442),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_443),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_318),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_474),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_446),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_452),
.Y(n_619)
);

NOR2xp67_ASAP7_75t_L g620 ( 
.A(n_454),
.B(n_2),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_461),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_319),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_325),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_476),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_489),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_328),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_343),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_496),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_345),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_498),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_520),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_509),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_348),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_515),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_352),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_519),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_530),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_535),
.Y(n_638)
);

NOR2xp67_ASAP7_75t_L g639 ( 
.A(n_337),
.B(n_2),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_L g640 ( 
.A(n_337),
.B(n_3),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_317),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_344),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_508),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_361),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_362),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_320),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_321),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_520),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_536),
.B(n_4),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_369),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_324),
.Y(n_651)
);

CKINVDCx16_ASAP7_75t_R g652 ( 
.A(n_468),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_371),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_373),
.B(n_4),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_326),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_376),
.B(n_5),
.Y(n_656)
);

BUFx2_ASAP7_75t_SL g657 ( 
.A(n_389),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_382),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_385),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_386),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_396),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_403),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_404),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_407),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_415),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_430),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_327),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_444),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_450),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_457),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_459),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_462),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_332),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_333),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_464),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_356),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_334),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_336),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_472),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_473),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_480),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_491),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_341),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_342),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_499),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_346),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_507),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_512),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_518),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_523),
.B(n_5),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_525),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_528),
.B(n_6),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_354),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_529),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_534),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_551),
.Y(n_696)
);

CKINVDCx8_ASAP7_75t_R g697 ( 
.A(n_539),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_551),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_557),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_557),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_642),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_550),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_577),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_560),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_584),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_601),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_652),
.B(n_657),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_547),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_548),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_605),
.B(n_356),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_642),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_549),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_552),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_642),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_641),
.B(n_339),
.Y(n_715)
);

CKINVDCx8_ASAP7_75t_R g716 ( 
.A(n_544),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_642),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_556),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_646),
.B(n_453),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_577),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_612),
.B(n_329),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_565),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_599),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_611),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_599),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_611),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_566),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_568),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_554),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_631),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_554),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_570),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_571),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_540),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_541),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_546),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_616),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_631),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_662),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_587),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_647),
.B(n_469),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_621),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_651),
.B(n_365),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_622),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_623),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_626),
.Y(n_746)
);

BUFx8_ASAP7_75t_L g747 ( 
.A(n_688),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_627),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_590),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_655),
.B(n_365),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_662),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_608),
.B(n_380),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_591),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_575),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_629),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_610),
.B(n_380),
.Y(n_756)
);

AND2x6_ASAP7_75t_L g757 ( 
.A(n_633),
.B(n_344),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_635),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_644),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_645),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_650),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_597),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_538),
.B(n_377),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_653),
.B(n_344),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_658),
.Y(n_765)
);

BUFx8_ASAP7_75t_L g766 ( 
.A(n_602),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_659),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_674),
.B(n_387),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_663),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_664),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_677),
.B(n_387),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_665),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_621),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_666),
.Y(n_774)
);

INVx6_ASAP7_75t_L g775 ( 
.A(n_567),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_678),
.B(n_398),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_683),
.B(n_398),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_691),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_583),
.B(n_531),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_684),
.B(n_411),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_607),
.B(n_411),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_668),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_691),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_671),
.A2(n_465),
.B(n_451),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_672),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_675),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_679),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_638),
.A2(n_417),
.B1(n_465),
.B2(n_451),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_680),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_681),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_682),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_686),
.B(n_676),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_685),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_654),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_SL g795 ( 
.A1(n_542),
.A2(n_482),
.B1(n_521),
.B2(n_510),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_687),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_643),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_689),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_695),
.B(n_482),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_694),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_582),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_660),
.B(n_510),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_792),
.B(n_595),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_723),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_734),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_731),
.B(n_648),
.Y(n_806)
);

INVx5_ASAP7_75t_L g807 ( 
.A(n_757),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_735),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_731),
.B(n_648),
.Y(n_809)
);

BUFx12f_ASAP7_75t_L g810 ( 
.A(n_747),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_729),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_798),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_794),
.B(n_661),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_710),
.B(n_596),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_697),
.Y(n_815)
);

NOR2x1p5_ASAP7_75t_L g816 ( 
.A(n_707),
.B(n_537),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_736),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_723),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_723),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_801),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_737),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_775),
.B(n_603),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_721),
.B(n_569),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_737),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_725),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_725),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_755),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_755),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_743),
.B(n_613),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_725),
.Y(n_830)
);

NAND3x1_ASAP7_75t_L g831 ( 
.A(n_788),
.B(n_592),
.C(n_649),
.Y(n_831)
);

OAI21xp33_ASAP7_75t_L g832 ( 
.A1(n_758),
.A2(n_690),
.B(n_656),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_740),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_758),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_796),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_779),
.B(n_573),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_796),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_729),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_798),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_729),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_798),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_739),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_730),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_739),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_738),
.Y(n_845)
);

INVx5_ASAP7_75t_L g846 ( 
.A(n_757),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_750),
.B(n_669),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_701),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_754),
.B(n_580),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_763),
.B(n_581),
.Y(n_850)
);

INVx5_ASAP7_75t_L g851 ( 
.A(n_757),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_794),
.B(n_670),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_708),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_701),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_709),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_794),
.B(n_521),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_739),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_701),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_776),
.B(n_585),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_715),
.B(n_593),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_749),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_753),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_710),
.A2(n_692),
.B1(n_639),
.B2(n_640),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_751),
.Y(n_864)
);

INVxp33_ASAP7_75t_L g865 ( 
.A(n_724),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_751),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_712),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_781),
.B(n_598),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_713),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_751),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_762),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_716),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_781),
.B(n_606),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_797),
.B(n_553),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_718),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_711),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_722),
.Y(n_877)
);

BUFx4f_ASAP7_75t_L g878 ( 
.A(n_775),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_711),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_719),
.B(n_614),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_777),
.B(n_615),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_780),
.B(n_618),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_702),
.B(n_619),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_727),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_704),
.B(n_624),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_778),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_728),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_747),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_752),
.B(n_600),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_741),
.B(n_625),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_732),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_705),
.B(n_423),
.Y(n_892)
);

AND2x2_ASAP7_75t_SL g893 ( 
.A(n_726),
.B(n_628),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_773),
.B(n_559),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_742),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_706),
.B(n_397),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_778),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_778),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_711),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_744),
.B(n_397),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_696),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_766),
.Y(n_902)
);

AO21x2_ASAP7_75t_L g903 ( 
.A1(n_768),
.A2(n_620),
.B(n_630),
.Y(n_903)
);

AO22x2_ASAP7_75t_L g904 ( 
.A1(n_814),
.A2(n_795),
.B1(n_752),
.B2(n_756),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_847),
.B(n_859),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_821),
.Y(n_906)
);

AO22x2_ASAP7_75t_L g907 ( 
.A1(n_814),
.A2(n_889),
.B1(n_874),
.B2(n_894),
.Y(n_907)
);

AO22x2_ASAP7_75t_L g908 ( 
.A1(n_889),
.A2(n_756),
.B1(n_542),
.B2(n_558),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_847),
.A2(n_667),
.B1(n_673),
.B2(n_693),
.Y(n_909)
);

AO22x2_ASAP7_75t_L g910 ( 
.A1(n_823),
.A2(n_555),
.B1(n_643),
.B2(n_771),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_833),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_878),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_824),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_850),
.B(n_561),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_861),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_862),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_827),
.Y(n_917)
);

OAI221xp5_ASAP7_75t_L g918 ( 
.A1(n_863),
.A2(n_802),
.B1(n_799),
.B2(n_733),
.C(n_746),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_815),
.B(n_783),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_803),
.A2(n_667),
.B1(n_673),
.B2(n_638),
.Y(n_920)
);

BUFx8_ASAP7_75t_L g921 ( 
.A(n_810),
.Y(n_921)
);

OAI221xp5_ASAP7_75t_L g922 ( 
.A1(n_863),
.A2(n_759),
.B1(n_760),
.B2(n_748),
.C(n_745),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_859),
.B(n_761),
.Y(n_923)
);

AND2x6_ASAP7_75t_L g924 ( 
.A(n_868),
.B(n_873),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_806),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_836),
.B(n_562),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_871),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_828),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_803),
.A2(n_767),
.B1(n_769),
.B2(n_765),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_834),
.Y(n_930)
);

NOR2xp67_ASAP7_75t_L g931 ( 
.A(n_872),
.B(n_632),
.Y(n_931)
);

NAND2x1p5_ASAP7_75t_L g932 ( 
.A(n_878),
.B(n_783),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_901),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_849),
.B(n_634),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_835),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_882),
.B(n_770),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_829),
.B(n_563),
.Y(n_937)
);

AO22x2_ASAP7_75t_L g938 ( 
.A1(n_806),
.A2(n_609),
.B1(n_617),
.B2(n_604),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_837),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_805),
.Y(n_940)
);

OAI21xp33_ASAP7_75t_L g941 ( 
.A1(n_829),
.A2(n_637),
.B(n_636),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_895),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_902),
.B(n_572),
.Y(n_943)
);

OAI221xp5_ASAP7_75t_L g944 ( 
.A1(n_832),
.A2(n_782),
.B1(n_787),
.B2(n_786),
.C(n_774),
.Y(n_944)
);

NAND2xp33_ASAP7_75t_L g945 ( 
.A(n_856),
.B(n_793),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_808),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_817),
.Y(n_947)
);

BUFx8_ASAP7_75t_L g948 ( 
.A(n_809),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_853),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_882),
.B(n_783),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_813),
.B(n_772),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_809),
.B(n_576),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_843),
.Y(n_953)
);

AOI22x1_ASAP7_75t_L g954 ( 
.A1(n_855),
.A2(n_789),
.B1(n_790),
.B2(n_785),
.Y(n_954)
);

AO22x2_ASAP7_75t_L g955 ( 
.A1(n_831),
.A2(n_579),
.B1(n_586),
.B2(n_578),
.Y(n_955)
);

NAND2x1p5_ASAP7_75t_L g956 ( 
.A(n_870),
.B(n_791),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_822),
.B(n_588),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_867),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_869),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_845),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_813),
.B(n_800),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_852),
.B(n_564),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_883),
.B(n_885),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_842),
.B(n_699),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_888),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_812),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_883),
.B(n_885),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_893),
.B(n_589),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_875),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_852),
.B(n_594),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_877),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_884),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_887),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_865),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_890),
.B(n_543),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_891),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_812),
.B(n_757),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_839),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_900),
.Y(n_979)
);

OAI221xp5_ASAP7_75t_L g980 ( 
.A1(n_832),
.A2(n_700),
.B1(n_699),
.B2(n_703),
.C(n_698),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_841),
.B(n_764),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_820),
.Y(n_982)
);

AO22x2_ASAP7_75t_L g983 ( 
.A1(n_881),
.A2(n_766),
.B1(n_545),
.B2(n_574),
.Y(n_983)
);

AO22x2_ASAP7_75t_L g984 ( 
.A1(n_881),
.A2(n_545),
.B1(n_574),
.B2(n_543),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_890),
.B(n_359),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_900),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_896),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_892),
.B(n_764),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_896),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_822),
.B(n_784),
.Y(n_990)
);

AO22x2_ASAP7_75t_L g991 ( 
.A1(n_860),
.A2(n_880),
.B1(n_844),
.B2(n_842),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_892),
.B(n_764),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_857),
.Y(n_993)
);

OAI21xp33_ASAP7_75t_L g994 ( 
.A1(n_857),
.A2(n_700),
.B(n_368),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_864),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_864),
.Y(n_996)
);

AO22x2_ASAP7_75t_L g997 ( 
.A1(n_844),
.A2(n_720),
.B1(n_8),
.B2(n_6),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_856),
.Y(n_998)
);

OR2x6_ASAP7_75t_L g999 ( 
.A(n_816),
.B(n_886),
.Y(n_999)
);

NAND2x1p5_ASAP7_75t_L g1000 ( 
.A(n_886),
.B(n_344),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_866),
.B(n_374),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_866),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_804),
.Y(n_1003)
);

AO22x2_ASAP7_75t_L g1004 ( 
.A1(n_897),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_856),
.B(n_897),
.Y(n_1005)
);

NAND2xp33_ASAP7_75t_L g1006 ( 
.A(n_856),
.B(n_397),
.Y(n_1006)
);

AO22x2_ASAP7_75t_L g1007 ( 
.A1(n_898),
.A2(n_13),
.B1(n_10),
.B2(n_11),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_905),
.B(n_903),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_963),
.B(n_967),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_934),
.B(n_898),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_923),
.B(n_903),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_936),
.B(n_811),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_950),
.B(n_811),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_926),
.B(n_838),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_951),
.B(n_838),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_909),
.B(n_840),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_931),
.B(n_840),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_914),
.B(n_848),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_941),
.B(n_848),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_961),
.B(n_818),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_SL g1021 ( 
.A(n_912),
.B(n_848),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_920),
.B(n_854),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_929),
.B(n_854),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_982),
.B(n_985),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_937),
.B(n_899),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_962),
.B(n_899),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_970),
.B(n_899),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_SL g1028 ( 
.A(n_940),
.B(n_858),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_SL g1029 ( 
.A(n_946),
.B(n_947),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_925),
.B(n_858),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_SL g1031 ( 
.A(n_949),
.B(n_858),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_987),
.B(n_819),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_989),
.B(n_906),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_925),
.B(n_876),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_932),
.B(n_876),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_975),
.B(n_879),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_958),
.B(n_959),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_969),
.B(n_879),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_971),
.B(n_825),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_972),
.B(n_826),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_913),
.B(n_830),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_973),
.B(n_851),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_976),
.B(n_851),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_917),
.B(n_851),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_942),
.B(n_11),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_928),
.B(n_846),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_930),
.B(n_846),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_935),
.B(n_846),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_SL g1049 ( 
.A(n_939),
.B(n_375),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_960),
.B(n_807),
.Y(n_1050)
);

NAND2xp33_ASAP7_75t_SL g1051 ( 
.A(n_979),
.B(n_379),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_998),
.B(n_807),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_986),
.B(n_381),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_924),
.B(n_388),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_1001),
.B(n_390),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_919),
.B(n_391),
.Y(n_1056)
);

NAND2xp33_ASAP7_75t_SL g1057 ( 
.A(n_993),
.B(n_392),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_999),
.B(n_924),
.Y(n_1058)
);

NAND2xp33_ASAP7_75t_SL g1059 ( 
.A(n_995),
.B(n_393),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_918),
.B(n_399),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_968),
.B(n_13),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_953),
.B(n_400),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_996),
.B(n_14),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_957),
.B(n_974),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_966),
.B(n_401),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_911),
.B(n_915),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_978),
.B(n_402),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_965),
.B(n_405),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_952),
.B(n_16),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_948),
.B(n_408),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_1002),
.B(n_409),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_1005),
.B(n_410),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_956),
.B(n_412),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_994),
.B(n_413),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_964),
.B(n_414),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_999),
.B(n_916),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_943),
.B(n_416),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_954),
.B(n_418),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_927),
.B(n_419),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_988),
.B(n_421),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_SL g1081 ( 
.A(n_977),
.B(n_422),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_907),
.B(n_18),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_992),
.B(n_425),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1003),
.B(n_426),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_1000),
.B(n_428),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_933),
.B(n_432),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_SL g1087 ( 
.A(n_1004),
.B(n_434),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_981),
.B(n_435),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_SL g1089 ( 
.A(n_1004),
.B(n_1007),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_L g1090 ( 
.A(n_1009),
.B(n_944),
.C(n_922),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1033),
.A2(n_1007),
.B1(n_991),
.B2(n_997),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1008),
.A2(n_980),
.B(n_990),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1024),
.B(n_904),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1032),
.A2(n_990),
.B(n_945),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1011),
.B(n_904),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1037),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1012),
.A2(n_1006),
.B(n_991),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1041),
.A2(n_1015),
.B(n_1039),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_1064),
.Y(n_1099)
);

INVxp67_ASAP7_75t_SL g1100 ( 
.A(n_1023),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_1058),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_SL g1102 ( 
.A(n_1076),
.B(n_921),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1060),
.A2(n_997),
.B1(n_907),
.B2(n_910),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1076),
.B(n_910),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_1016),
.B(n_938),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_SL g1106 ( 
.A1(n_1054),
.A2(n_20),
.B(n_21),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1053),
.A2(n_955),
.B1(n_984),
.B2(n_983),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1069),
.B(n_938),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1066),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1013),
.A2(n_490),
.B(n_397),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1020),
.Y(n_1111)
);

AOI221xp5_ASAP7_75t_L g1112 ( 
.A1(n_1089),
.A2(n_984),
.B1(n_955),
.B2(n_983),
.C(n_908),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_1082),
.Y(n_1113)
);

AO32x2_ASAP7_75t_L g1114 ( 
.A1(n_1087),
.A2(n_908),
.A3(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_1045),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1010),
.B(n_20),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1061),
.B(n_22),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1077),
.B(n_23),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_SL g1119 ( 
.A1(n_1025),
.A2(n_526),
.B(n_438),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1029),
.A2(n_437),
.B(n_441),
.C(n_440),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1080),
.A2(n_447),
.B(n_445),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1022),
.B(n_1018),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1078),
.A2(n_490),
.B(n_397),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1038),
.A2(n_490),
.B(n_397),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1070),
.B(n_25),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1014),
.B(n_26),
.Y(n_1126)
);

AOI31xp67_ASAP7_75t_L g1127 ( 
.A1(n_1019),
.A2(n_490),
.A3(n_717),
.B(n_714),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1040),
.A2(n_1026),
.B(n_1083),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1027),
.A2(n_1088),
.B(n_1035),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1063),
.A2(n_490),
.A3(n_717),
.B(n_714),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1055),
.A2(n_456),
.B(n_449),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_1068),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1030),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1063),
.A2(n_495),
.B(n_463),
.C(n_467),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1051),
.A2(n_470),
.B(n_460),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_1021),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_SL g1137 ( 
.A(n_1062),
.B(n_481),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1049),
.A2(n_502),
.B(n_484),
.C(n_485),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1074),
.A2(n_488),
.B(n_483),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1072),
.A2(n_497),
.B(n_494),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1034),
.Y(n_1141)
);

BUFx8_ASAP7_75t_L g1142 ( 
.A(n_1057),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1028),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_1059),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1031),
.A2(n_1075),
.B(n_1081),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1036),
.A2(n_490),
.B(n_71),
.Y(n_1146)
);

AOI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1044),
.A2(n_717),
.B(n_714),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1017),
.Y(n_1148)
);

AO31x2_ASAP7_75t_L g1149 ( 
.A1(n_1084),
.A2(n_526),
.A3(n_187),
.B(n_188),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1050),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1071),
.A2(n_26),
.B(n_29),
.C(n_30),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1073),
.B(n_501),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1065),
.A2(n_505),
.B(n_503),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1042),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1079),
.A2(n_511),
.B(n_506),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1043),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1056),
.B(n_30),
.Y(n_1157)
);

NOR3xp33_ASAP7_75t_L g1158 ( 
.A(n_1067),
.B(n_517),
.C(n_514),
.Y(n_1158)
);

OAI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1117),
.A2(n_1086),
.B1(n_1085),
.B2(n_1047),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1109),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1096),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1111),
.B(n_1052),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1133),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1150),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_SL g1165 ( 
.A1(n_1134),
.A2(n_1048),
.B(n_1046),
.C(n_35),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1141),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1124),
.A2(n_75),
.B(n_70),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1110),
.A2(n_83),
.B(n_82),
.Y(n_1168)
);

BUFx2_ASAP7_75t_R g1169 ( 
.A(n_1101),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1112),
.A2(n_526),
.B1(n_524),
.B2(n_36),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_SL g1171 ( 
.A(n_1102),
.B(n_31),
.Y(n_1171)
);

CKINVDCx8_ASAP7_75t_R g1172 ( 
.A(n_1144),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_1136),
.B(n_84),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1132),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1090),
.A2(n_31),
.B(n_34),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1122),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1113),
.B(n_34),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1092),
.A2(n_36),
.B(n_37),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1126),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1104),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_L g1181 ( 
.A1(n_1097),
.A2(n_39),
.B(n_41),
.C(n_42),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1123),
.A2(n_91),
.B(n_90),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1146),
.A2(n_100),
.B(n_93),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1113),
.B(n_43),
.Y(n_1184)
);

OAI221xp5_ASAP7_75t_L g1185 ( 
.A1(n_1090),
.A2(n_1107),
.B1(n_1091),
.B2(n_1103),
.C(n_1137),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1147),
.A2(n_1128),
.B(n_1129),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1154),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1100),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1094),
.A2(n_102),
.B(n_101),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1156),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1116),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1115),
.B(n_44),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1104),
.A2(n_1108),
.B1(n_1105),
.B2(n_1095),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1148),
.Y(n_1194)
);

AOI21xp33_ASAP7_75t_L g1195 ( 
.A1(n_1093),
.A2(n_45),
.B(n_46),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1098),
.B(n_49),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1142),
.Y(n_1197)
);

AOI221xp5_ASAP7_75t_L g1198 ( 
.A1(n_1125),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.C(n_54),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1157),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_1199)
);

AOI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1145),
.A2(n_200),
.B(n_305),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1116),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1106),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1151),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1118),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1142),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_L g1206 ( 
.A(n_1137),
.B(n_55),
.C(n_56),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1099),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1114),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1136),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1143),
.A2(n_57),
.B(n_58),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_L g1211 ( 
.A(n_1152),
.B(n_58),
.C(n_59),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1114),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1114),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1136),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1143),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1130),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1120),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1149),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1158),
.B(n_103),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1127),
.A2(n_207),
.B(n_299),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1119),
.A2(n_201),
.B(n_296),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1155),
.A2(n_66),
.B(n_67),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1139),
.A2(n_104),
.B(n_105),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1138),
.A2(n_1121),
.B(n_1140),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1149),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1218),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1216),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_SL g1228 ( 
.A(n_1172),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1186),
.A2(n_1167),
.B(n_1168),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1208),
.B(n_1130),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1189),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1205),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1225),
.Y(n_1233)
);

BUFx2_ASAP7_75t_SL g1234 ( 
.A(n_1209),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1161),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1185),
.A2(n_1135),
.B1(n_1131),
.B2(n_1153),
.Y(n_1236)
);

INVx11_ASAP7_75t_L g1237 ( 
.A(n_1169),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1200),
.A2(n_1183),
.B(n_1220),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1212),
.B(n_106),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1166),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1202),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1176),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1190),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1185),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1179),
.B(n_118),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1196),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_1209),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1191),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1220),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1196),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1213),
.B(n_121),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1188),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1182),
.A2(n_123),
.B(n_124),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1194),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1207),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1160),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1163),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1164),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1187),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1162),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1182),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_SL g1262 ( 
.A1(n_1222),
.A2(n_125),
.B(n_126),
.C(n_129),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1178),
.A2(n_130),
.B(n_132),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1193),
.B(n_137),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1192),
.B(n_311),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1201),
.B(n_139),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1184),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1162),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1181),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1174),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1223),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1214),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1197),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1173),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1181),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1175),
.B(n_142),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1204),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1173),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1184),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1184),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1203),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1177),
.B(n_146),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1210),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1210),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1221),
.A2(n_147),
.B(n_150),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1219),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1215),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1219),
.Y(n_1288)
);

NAND2xp33_ASAP7_75t_R g1289 ( 
.A(n_1273),
.B(n_1267),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_R g1290 ( 
.A(n_1232),
.B(n_1171),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1286),
.B(n_1159),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1260),
.B(n_1198),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1255),
.B(n_1206),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1255),
.B(n_1211),
.Y(n_1294)
);

NAND2xp33_ASAP7_75t_R g1295 ( 
.A(n_1267),
.B(n_1171),
.Y(n_1295)
);

OR2x6_ASAP7_75t_L g1296 ( 
.A(n_1286),
.B(n_1215),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1255),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_R g1298 ( 
.A(n_1228),
.B(n_1169),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1288),
.B(n_1199),
.Y(n_1299)
);

NAND2xp33_ASAP7_75t_R g1300 ( 
.A(n_1282),
.B(n_1224),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_R g1301 ( 
.A(n_1270),
.B(n_1180),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_R g1302 ( 
.A(n_1270),
.B(n_151),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1277),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1240),
.B(n_1199),
.Y(n_1304)
);

XNOR2xp5_ASAP7_75t_L g1305 ( 
.A(n_1237),
.B(n_1198),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1237),
.Y(n_1306)
);

NAND2xp33_ASAP7_75t_R g1307 ( 
.A(n_1282),
.B(n_1224),
.Y(n_1307)
);

NAND2xp33_ASAP7_75t_R g1308 ( 
.A(n_1274),
.B(n_154),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1242),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1279),
.B(n_1280),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1243),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1234),
.B(n_1217),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1260),
.B(n_1195),
.Y(n_1313)
);

XNOR2xp5_ASAP7_75t_L g1314 ( 
.A(n_1279),
.B(n_1170),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1272),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1278),
.B(n_1165),
.Y(n_1316)
);

BUFx10_ASAP7_75t_L g1317 ( 
.A(n_1272),
.Y(n_1317)
);

NAND2xp33_ASAP7_75t_R g1318 ( 
.A(n_1278),
.B(n_159),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_R g1319 ( 
.A(n_1278),
.B(n_161),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1247),
.B(n_164),
.Y(n_1320)
);

NAND2xp33_ASAP7_75t_R g1321 ( 
.A(n_1245),
.B(n_165),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1234),
.B(n_166),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1247),
.B(n_167),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1268),
.B(n_178),
.Y(n_1324)
);

XNOR2xp5_ASAP7_75t_L g1325 ( 
.A(n_1248),
.B(n_179),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1235),
.Y(n_1326)
);

XNOR2xp5_ASAP7_75t_L g1327 ( 
.A(n_1254),
.B(n_181),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1247),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_R g1329 ( 
.A(n_1265),
.B(n_184),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1247),
.B(n_191),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_R g1331 ( 
.A(n_1246),
.B(n_192),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1235),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1250),
.B(n_194),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1256),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_R g1335 ( 
.A(n_1250),
.B(n_1287),
.Y(n_1335)
);

BUFx12f_ASAP7_75t_L g1336 ( 
.A(n_1264),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1252),
.B(n_195),
.Y(n_1337)
);

NAND2xp33_ASAP7_75t_R g1338 ( 
.A(n_1276),
.B(n_197),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1291),
.B(n_1283),
.Y(n_1339)
);

INVx5_ASAP7_75t_L g1340 ( 
.A(n_1312),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1303),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1310),
.B(n_1230),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1311),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1297),
.B(n_1241),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1309),
.B(n_1241),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1326),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1335),
.B(n_1281),
.Y(n_1347)
);

NOR2x1_ASAP7_75t_L g1348 ( 
.A(n_1315),
.B(n_1281),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1305),
.A2(n_1287),
.B(n_1263),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1317),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1332),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1328),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1334),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1296),
.B(n_1284),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1304),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1313),
.B(n_1226),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1312),
.A2(n_1244),
.B1(n_1236),
.B2(n_1251),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1299),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1292),
.B(n_1226),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1294),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1294),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1293),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1333),
.B(n_1233),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1337),
.B(n_1239),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1316),
.B(n_1269),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1324),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1325),
.B(n_1269),
.Y(n_1367)
);

OAI221xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1314),
.A2(n_1251),
.B1(n_1264),
.B2(n_1275),
.C(n_1266),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1336),
.B(n_1275),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1322),
.B(n_1261),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1322),
.B(n_1231),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1300),
.B(n_1227),
.Y(n_1372)
);

NAND3xp33_ASAP7_75t_L g1373 ( 
.A(n_1349),
.B(n_1307),
.C(n_1338),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1340),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1339),
.B(n_1231),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1357),
.A2(n_1321),
.B1(n_1295),
.B2(n_1318),
.Y(n_1376)
);

AOI221xp5_ASAP7_75t_L g1377 ( 
.A1(n_1368),
.A2(n_1290),
.B1(n_1301),
.B2(n_1302),
.C(n_1331),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1344),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1346),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1367),
.A2(n_1327),
.B1(n_1330),
.B2(n_1323),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1365),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1340),
.B(n_1298),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1355),
.B(n_1261),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1351),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1347),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1343),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1367),
.A2(n_1257),
.B1(n_1259),
.B2(n_1258),
.Y(n_1387)
);

OAI211xp5_ASAP7_75t_L g1388 ( 
.A1(n_1341),
.A2(n_1329),
.B(n_1262),
.C(n_1319),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1343),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1345),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1342),
.B(n_1306),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1351),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1356),
.B(n_1259),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1369),
.B(n_1289),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1345),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1394),
.B(n_1340),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1381),
.B(n_1363),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1385),
.B(n_1350),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1381),
.B(n_1363),
.Y(n_1399)
);

INVxp33_ASAP7_75t_L g1400 ( 
.A(n_1373),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1386),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1389),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1390),
.B(n_1369),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_SL g1404 ( 
.A1(n_1382),
.A2(n_1371),
.B(n_1347),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1383),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1393),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1395),
.B(n_1354),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1378),
.B(n_1352),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1391),
.B(n_1350),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1383),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1379),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1403),
.B(n_1380),
.Y(n_1412)
);

OAI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1400),
.A2(n_1376),
.B1(n_1377),
.B2(n_1340),
.Y(n_1413)
);

NAND2xp33_ASAP7_75t_SL g1414 ( 
.A(n_1403),
.B(n_1361),
.Y(n_1414)
);

INVxp33_ASAP7_75t_SL g1415 ( 
.A(n_1409),
.Y(n_1415)
);

OAI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1400),
.A2(n_1377),
.B1(n_1388),
.B2(n_1387),
.C(n_1366),
.Y(n_1416)
);

AO221x2_ASAP7_75t_L g1417 ( 
.A1(n_1407),
.A2(n_1360),
.B1(n_1362),
.B2(n_1364),
.C(n_1358),
.Y(n_1417)
);

NOR2x1_ASAP7_75t_L g1418 ( 
.A(n_1404),
.B(n_1348),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1410),
.B(n_1359),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1406),
.B(n_1361),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1397),
.B(n_1339),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1409),
.Y(n_1422)
);

NOR2x1_ASAP7_75t_L g1423 ( 
.A(n_1398),
.B(n_1375),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1399),
.B(n_1339),
.Y(n_1424)
);

OAI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1396),
.A2(n_1366),
.B1(n_1308),
.B2(n_1372),
.C(n_1353),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1396),
.B(n_1374),
.Y(n_1426)
);

NOR2x1_ASAP7_75t_L g1427 ( 
.A(n_1418),
.B(n_1422),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1419),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1412),
.Y(n_1429)
);

INVx4_ASAP7_75t_L g1430 ( 
.A(n_1420),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1415),
.B(n_1401),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1413),
.A2(n_1405),
.B(n_1402),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_SL g1433 ( 
.A1(n_1416),
.A2(n_1405),
.B(n_1352),
.C(n_1271),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1421),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1417),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1424),
.Y(n_1436)
);

NOR2x1_ASAP7_75t_L g1437 ( 
.A(n_1423),
.B(n_1426),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1414),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1425),
.Y(n_1439)
);

NOR3xp33_ASAP7_75t_L g1440 ( 
.A(n_1427),
.B(n_1370),
.C(n_1371),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1430),
.B(n_1408),
.Y(n_1441)
);

NOR2x1_ASAP7_75t_L g1442 ( 
.A(n_1429),
.B(n_1320),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1431),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1428),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1443),
.B(n_1438),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1441),
.B(n_1435),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1444),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1442),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1440),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1446),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1445),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1448),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1447),
.B(n_1439),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1451),
.B(n_1449),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1450),
.B(n_1437),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1453),
.A2(n_1433),
.B(n_1432),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1452),
.B(n_1434),
.Y(n_1457)
);

NOR2x1_ASAP7_75t_L g1458 ( 
.A(n_1450),
.B(n_1436),
.Y(n_1458)
);

OA22x2_ASAP7_75t_L g1459 ( 
.A1(n_1455),
.A2(n_1434),
.B1(n_1374),
.B2(n_1411),
.Y(n_1459)
);

OAI211xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1458),
.A2(n_1249),
.B(n_1271),
.C(n_1231),
.Y(n_1460)
);

AOI221xp5_ASAP7_75t_L g1461 ( 
.A1(n_1456),
.A2(n_1261),
.B1(n_1249),
.B2(n_1392),
.C(n_1384),
.Y(n_1461)
);

NOR2x1_ASAP7_75t_L g1462 ( 
.A(n_1460),
.B(n_1454),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1461),
.Y(n_1463)
);

NOR4xp75_ASAP7_75t_L g1464 ( 
.A(n_1459),
.B(n_1457),
.C(n_1271),
.D(n_1249),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1462),
.B(n_1261),
.Y(n_1465)
);

NAND2xp33_ASAP7_75t_SL g1466 ( 
.A(n_1463),
.B(n_1249),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_R g1467 ( 
.A(n_1464),
.B(n_208),
.Y(n_1467)
);

NAND4xp75_ASAP7_75t_L g1468 ( 
.A(n_1465),
.B(n_1253),
.C(n_1285),
.D(n_214),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1466),
.Y(n_1469)
);

NAND4xp75_ASAP7_75t_L g1470 ( 
.A(n_1467),
.B(n_210),
.C(n_211),
.D(n_219),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1469),
.A2(n_1238),
.B1(n_1229),
.B2(n_235),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1470),
.B(n_1229),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1468),
.Y(n_1473)
);

AO22x2_ASAP7_75t_L g1474 ( 
.A1(n_1472),
.A2(n_220),
.B1(n_234),
.B2(n_242),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1473),
.B(n_245),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1471),
.Y(n_1476)
);

NAND2xp33_ASAP7_75t_R g1477 ( 
.A(n_1473),
.B(n_295),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1474),
.A2(n_1476),
.B1(n_1475),
.B2(n_1477),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1478),
.B(n_257),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_L g1480 ( 
.A(n_1479),
.B(n_258),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1480),
.Y(n_1481)
);

AOI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1481),
.A2(n_259),
.B1(n_262),
.B2(n_264),
.C(n_266),
.Y(n_1482)
);

AOI211xp5_ASAP7_75t_L g1483 ( 
.A1(n_1482),
.A2(n_277),
.B(n_281),
.C(n_282),
.Y(n_1483)
);


endmodule