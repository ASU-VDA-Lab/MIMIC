module fake_jpeg_16058_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_5),
.B(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_54),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_58),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_64),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_50),
.B1(n_51),
.B2(n_46),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_47),
.B1(n_45),
.B2(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_0),
.Y(n_73)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_72),
.Y(n_79)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_47),
.C(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_1),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_82),
.B1(n_71),
.B2(n_3),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_1),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_64),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_85),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_44),
.B1(n_40),
.B2(n_4),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_2),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_71),
.B1(n_25),
.B2(n_26),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_2),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_95),
.B(n_78),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_3),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_95),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_4),
.C(n_5),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_99),
.B(n_101),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_28),
.B(n_38),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_6),
.B(n_7),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_102),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_106),
.A2(n_100),
.B1(n_8),
.B2(n_11),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_109),
.Y(n_112)
);

AO32x1_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_100),
.A3(n_97),
.B1(n_89),
.B2(n_7),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_107),
.A3(n_13),
.B1(n_15),
.B2(n_21),
.C1(n_24),
.C2(n_27),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_113),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_116),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_112),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_118),
.B(n_29),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_10),
.B(n_30),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_36),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_37),
.Y(n_125)
);


endmodule