module fake_jpeg_1211_n_181 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_181);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_82),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_43),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

OA21x2_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_44),
.B(n_64),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_90),
.B1(n_98),
.B2(n_95),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_91),
.Y(n_109)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_48),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_95),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_44),
.B(n_53),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_97),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_56),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_107),
.Y(n_130)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_102),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_54),
.Y(n_123)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_60),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_115),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_60),
.B1(n_59),
.B2(n_61),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_59),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_1),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_1),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_124),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_123),
.A2(n_128),
.B(n_12),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_54),
.B1(n_4),
.B2(n_5),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_129),
.B1(n_132),
.B2(n_137),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_102),
.B1(n_114),
.B2(n_11),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_6),
.B(n_7),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_27),
.B1(n_37),
.B2(n_36),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_21),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_24),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_9),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_103),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_120),
.B(n_12),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_148),
.B(n_154),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_149),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_13),
.B1(n_14),
.B2(n_18),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_150),
.B(n_25),
.C(n_29),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_126),
.B(n_127),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_134),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_41),
.B(n_22),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_150),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_136),
.C(n_129),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.C(n_144),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_30),
.C(n_31),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_152),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_164),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_159),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_165),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_167),
.Y(n_171)
);

OAI22x1_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_151),
.B1(n_148),
.B2(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_155),
.C(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_173),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_164),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_170),
.B1(n_161),
.B2(n_172),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_172),
.Y(n_179)
);

NAND4xp25_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_151),
.C(n_157),
.D(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_34),
.Y(n_181)
);


endmodule