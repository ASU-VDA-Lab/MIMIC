module fake_jpeg_12911_n_88 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_3),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_5),
.B(n_10),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_46),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_30),
.B1(n_29),
.B2(n_33),
.Y(n_50)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_1),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_64),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_16),
.B(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_41),
.B1(n_44),
.B2(n_42),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_62),
.B1(n_63),
.B2(n_7),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_31),
.C(n_28),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_3),
.C(n_7),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_35),
.B1(n_32),
.B2(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_35),
.B1(n_32),
.B2(n_4),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_2),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_32),
.B(n_6),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_76),
.C(n_69),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_57),
.B(n_58),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_69),
.B1(n_73),
.B2(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_8),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_79),
.B(n_74),
.C(n_67),
.D(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_77),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_81),
.C(n_14),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_13),
.Y(n_85)
);

OAI31xp33_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_15),
.A3(n_18),
.B(n_20),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_22),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_27),
.Y(n_88)
);


endmodule