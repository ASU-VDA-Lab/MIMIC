module fake_jpeg_11073_n_496 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_496);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_496;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_51),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_52),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_88),
.Y(n_111)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_57),
.B(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_16),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_15),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_71),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_15),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_82),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_43),
.B(n_14),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_19),
.B(n_14),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_40),
.B(n_1),
.Y(n_88)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_91),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_93),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_97),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_19),
.B(n_2),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_96),
.Y(n_126)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_41),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_40),
.B1(n_48),
.B2(n_22),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_99),
.A2(n_137),
.B1(n_140),
.B2(n_143),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_34),
.B1(n_41),
.B2(n_21),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_101),
.A2(n_129),
.B1(n_147),
.B2(n_38),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_56),
.A2(n_48),
.B1(n_25),
.B2(n_21),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_119),
.B1(n_122),
.B2(n_133),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_53),
.A2(n_40),
.B1(n_48),
.B2(n_25),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_68),
.B(n_24),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_121),
.B(n_46),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_63),
.A2(n_48),
.B1(n_21),
.B2(n_26),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_51),
.A2(n_41),
.B1(n_26),
.B2(n_25),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_65),
.A2(n_26),
.B1(n_45),
.B2(n_30),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_49),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_30),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_59),
.A2(n_49),
.B1(n_47),
.B2(n_28),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_69),
.A2(n_75),
.B1(n_76),
.B2(n_72),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_73),
.A2(n_47),
.B1(n_28),
.B2(n_29),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_78),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_62),
.B(n_39),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_97),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_74),
.A2(n_39),
.B1(n_24),
.B2(n_29),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_30),
.B1(n_153),
.B2(n_112),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_70),
.B(n_46),
.C(n_45),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_55),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_188),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_99),
.A2(n_54),
.B1(n_64),
.B2(n_96),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_155),
.Y(n_242)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_158),
.Y(n_253)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_159),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_160),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_161),
.B(n_170),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_162),
.A2(n_139),
.B1(n_144),
.B2(n_100),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_163),
.B(n_173),
.Y(n_212)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_166),
.B(n_192),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_117),
.A2(n_50),
.B1(n_66),
.B2(n_60),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_167),
.A2(n_190),
.B(n_205),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_94),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_180),
.C(n_182),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_169),
.A2(n_171),
.B1(n_194),
.B2(n_202),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_111),
.A2(n_93),
.B1(n_92),
.B2(n_91),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_98),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_119),
.A2(n_90),
.B1(n_81),
.B2(n_79),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_175),
.A2(n_146),
.B1(n_131),
.B2(n_134),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_2),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_3),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_109),
.B(n_141),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_104),
.B(n_77),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_181),
.B(n_183),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_108),
.A2(n_89),
.B(n_38),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_185),
.Y(n_246)
);

BUFx2_ASAP7_75t_SL g186 ( 
.A(n_151),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_117),
.B(n_67),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_189),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_114),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_125),
.B(n_85),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_132),
.A2(n_35),
.B1(n_23),
.B2(n_5),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_109),
.B(n_3),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_191),
.B(n_197),
.Y(n_244)
);

NAND2xp67_ASAP7_75t_SL g192 ( 
.A(n_148),
.B(n_35),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_102),
.B(n_3),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_201),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_128),
.A2(n_23),
.B1(n_4),
.B2(n_5),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_196),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_102),
.B(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_200),
.Y(n_243)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_138),
.A2(n_23),
.B1(n_4),
.B2(n_6),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_204),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_114),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_126),
.B(n_3),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

AO22x1_ASAP7_75t_L g207 ( 
.A1(n_132),
.A2(n_23),
.B1(n_4),
.B2(n_6),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_130),
.B(n_113),
.C(n_8),
.Y(n_226)
);

AOI32xp33_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_126),
.A3(n_130),
.B1(n_113),
.B2(n_114),
.Y(n_208)
);

AOI31xp33_ASAP7_75t_SL g261 ( 
.A1(n_208),
.A2(n_167),
.A3(n_192),
.B(n_190),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_154),
.A2(n_120),
.B1(n_149),
.B2(n_103),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_216),
.A2(n_221),
.B1(n_230),
.B2(n_240),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_172),
.A2(n_149),
.B1(n_120),
.B2(n_103),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_223),
.B(n_163),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_226),
.A2(n_193),
.B(n_185),
.C(n_200),
.Y(n_294)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_228),
.Y(n_292)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_172),
.A2(n_127),
.B1(n_131),
.B2(n_134),
.Y(n_230)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_235),
.A2(n_198),
.B1(n_174),
.B2(n_165),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_239),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_162),
.A2(n_127),
.B1(n_146),
.B2(n_134),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_199),
.A2(n_144),
.B1(n_100),
.B2(n_105),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_241),
.A2(n_185),
.B1(n_207),
.B2(n_196),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_170),
.B(n_146),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_249),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_166),
.B(n_4),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_166),
.B(n_7),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_161),
.Y(n_268)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_160),
.A2(n_105),
.B1(n_23),
.B2(n_10),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_255),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_257),
.B(n_264),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_199),
.B(n_203),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_259),
.A2(n_265),
.B(n_290),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_261),
.B(n_294),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_176),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_262),
.B(n_271),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_214),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_217),
.A2(n_160),
.B(n_182),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_238),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_268),
.B(n_274),
.Y(n_338)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_242),
.A2(n_169),
.B1(n_179),
.B2(n_155),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_270),
.A2(n_280),
.B1(n_295),
.B2(n_230),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_183),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_213),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_272),
.B(n_279),
.Y(n_313)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_227),
.B(n_188),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_158),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_283),
.C(n_293),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_213),
.B(n_168),
.C(n_180),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_250),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_205),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_288),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_209),
.B(n_168),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_242),
.A2(n_179),
.B1(n_155),
.B2(n_171),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_282),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_223),
.B(n_204),
.Y(n_283)
);

AO21x2_ASAP7_75t_L g284 ( 
.A1(n_240),
.A2(n_156),
.B(n_155),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_284),
.A2(n_287),
.B1(n_299),
.B2(n_256),
.Y(n_325)
);

AOI22x1_ASAP7_75t_SL g285 ( 
.A1(n_221),
.A2(n_202),
.B1(n_194),
.B2(n_207),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g332 ( 
.A1(n_285),
.A2(n_297),
.B(n_237),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_232),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_296),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_234),
.B(n_205),
.Y(n_288)
);

INVx13_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

INVx13_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_232),
.B(n_180),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_201),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_222),
.B(n_184),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_226),
.A2(n_193),
.B(n_164),
.C(n_159),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_234),
.B(n_157),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_231),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_222),
.B(n_8),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_219),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_236),
.B(n_249),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_247),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_288),
.C(n_301),
.Y(n_351)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_307),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_225),
.Y(n_308)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_308),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_328),
.B1(n_331),
.B2(n_284),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_310),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_259),
.A2(n_265),
.B(n_254),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_314),
.A2(n_326),
.B(n_298),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_225),
.Y(n_316)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_284),
.A2(n_211),
.B1(n_291),
.B2(n_270),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_317),
.A2(n_320),
.B1(n_325),
.B2(n_332),
.Y(n_346)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_318),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_284),
.A2(n_211),
.B1(n_235),
.B2(n_254),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_255),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_321),
.A2(n_332),
.B(n_334),
.Y(n_366)
);

AND2x2_ASAP7_75t_SL g324 ( 
.A(n_277),
.B(n_286),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_324),
.A2(n_335),
.B(n_278),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_294),
.A2(n_234),
.B(n_233),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_280),
.A2(n_256),
.B1(n_224),
.B2(n_220),
.Y(n_328)
);

OAI32xp33_ASAP7_75t_L g329 ( 
.A1(n_260),
.A2(n_247),
.A3(n_237),
.B1(n_251),
.B2(n_218),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_295),
.Y(n_344)
);

XNOR2x1_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_341),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_297),
.A2(n_252),
.B1(n_210),
.B2(n_228),
.Y(n_331)
);

AND2x6_ASAP7_75t_L g334 ( 
.A(n_272),
.B(n_229),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_268),
.B(n_218),
.Y(n_335)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_269),
.Y(n_339)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_339),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_260),
.B(n_231),
.Y(n_340)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_340),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_329),
.Y(n_342)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

XNOR2x1_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_341),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_345),
.A2(n_347),
.B1(n_363),
.B2(n_372),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_346),
.A2(n_360),
.B1(n_361),
.B2(n_347),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_309),
.A2(n_328),
.B1(n_284),
.B2(n_317),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_313),
.B(n_279),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_349),
.C(n_350),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_290),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_303),
.B(n_290),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_368),
.C(n_371),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_352),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_330),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_353),
.B(n_356),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_315),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_357),
.A2(n_331),
.B(n_321),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_322),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_332),
.A2(n_258),
.B1(n_284),
.B2(n_285),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_360),
.A2(n_361),
.B1(n_346),
.B2(n_357),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_258),
.B1(n_261),
.B2(n_291),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_319),
.A2(n_275),
.B1(n_299),
.B2(n_273),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_314),
.A2(n_305),
.B(n_326),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_364),
.A2(n_306),
.B(n_335),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_324),
.B(n_298),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_315),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_369),
.B(n_333),
.Y(n_401)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_302),
.Y(n_370)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_282),
.C(n_281),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_319),
.A2(n_293),
.B1(n_257),
.B2(n_292),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_364),
.A2(n_305),
.B(n_334),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_375),
.A2(n_383),
.B(n_388),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_376),
.A2(n_385),
.B1(n_397),
.B2(n_311),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_377),
.B(n_378),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_365),
.Y(n_380)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_380),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_350),
.B(n_322),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_384),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_367),
.Y(n_389)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_372),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_390),
.B(n_402),
.Y(n_412)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_391),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_349),
.B(n_340),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_336),
.Y(n_425)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_393),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_337),
.C(n_339),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_399),
.C(n_362),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_358),
.A2(n_333),
.B1(n_336),
.B2(n_311),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_355),
.B(n_333),
.Y(n_398)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_398),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_351),
.B(n_371),
.C(n_374),
.Y(n_399)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_401),
.Y(n_424)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_419),
.Y(n_443)
);

NOR3xp33_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_312),
.C(n_323),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_423),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_398),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_389),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_409),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_394),
.A2(n_333),
.B1(n_343),
.B2(n_363),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_410),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_399),
.C(n_379),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_418),
.C(n_414),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_394),
.A2(n_344),
.B1(n_366),
.B2(n_302),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_415),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_387),
.B(n_379),
.C(n_395),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_374),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_377),
.B(n_392),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_425),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_421),
.A2(n_402),
.B1(n_393),
.B2(n_391),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_375),
.B(n_366),
.Y(n_423)
);

FAx1_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_383),
.CI(n_397),
.CON(n_426),
.SN(n_426)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_439),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_413),
.A2(n_382),
.B(n_388),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_427),
.A2(n_263),
.B(n_266),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_429),
.B(n_436),
.Y(n_458)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_418),
.C(n_404),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_435),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_424),
.B(n_381),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_378),
.C(n_385),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_437),
.Y(n_448)
);

FAx1_ASAP7_75t_SL g438 ( 
.A(n_416),
.B(n_380),
.CI(n_327),
.CON(n_438),
.SN(n_438)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_441),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_423),
.A2(n_396),
.B1(n_359),
.B2(n_373),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_444),
.Y(n_455)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_407),
.B(n_327),
.Y(n_444)
);

AOI322xp5_ASAP7_75t_SL g445 ( 
.A1(n_428),
.A2(n_421),
.A3(n_416),
.B1(n_406),
.B2(n_422),
.C1(n_289),
.C2(n_419),
.Y(n_445)
);

BUFx24_ASAP7_75t_SL g470 ( 
.A(n_445),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_420),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_447),
.B(n_450),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_425),
.C(n_417),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_443),
.B(n_408),
.C(n_263),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_454),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_453),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_436),
.C(n_442),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_266),
.C(n_310),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_440),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_318),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_459),
.B(n_439),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_465),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_432),
.Y(n_462)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_462),
.Y(n_474)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_448),
.Y(n_464)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_464),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_457),
.A2(n_431),
.B1(n_444),
.B2(n_433),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_468),
.Y(n_480)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_446),
.Y(n_467)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_467),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_450),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_430),
.Y(n_469)
);

AOI322xp5_ASAP7_75t_L g479 ( 
.A1(n_469),
.A2(n_456),
.A3(n_438),
.B1(n_455),
.B2(n_459),
.C1(n_289),
.C2(n_373),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_449),
.B(n_426),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_472),
.A2(n_426),
.B(n_463),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_481),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_463),
.A2(n_449),
.B1(n_454),
.B2(n_455),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_478),
.B(n_479),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_472),
.A2(n_438),
.B(n_276),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_480),
.A2(n_471),
.B(n_470),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_484),
.A2(n_486),
.B(n_487),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_462),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_485),
.A2(n_477),
.B1(n_481),
.B2(n_475),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_461),
.C(n_251),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_478),
.C(n_476),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_489),
.B(n_485),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_210),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_490),
.B(n_491),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_483),
.A2(n_13),
.B(n_11),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_488),
.Y(n_494)
);

AO21x1_ASAP7_75t_L g495 ( 
.A1(n_494),
.A2(n_492),
.B(n_11),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_495),
.A2(n_12),
.B(n_400),
.Y(n_496)
);


endmodule