module fake_jpeg_29479_n_398 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_398);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_398;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_61),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_65),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_23),
.B(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_79),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_30),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_0),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

CKINVDCx9p33_ASAP7_75t_R g81 ( 
.A(n_33),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_81),
.Y(n_111)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_47),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_118),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_32),
.B1(n_42),
.B2(n_34),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_95),
.A2(n_100),
.B1(n_125),
.B2(n_32),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_44),
.B1(n_40),
.B2(n_39),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_64),
.B(n_50),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_123),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx5_ASAP7_75t_SL g161 ( 
.A(n_106),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_31),
.Y(n_118)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_58),
.B(n_50),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_47),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_52),
.A2(n_37),
.B1(n_34),
.B2(n_35),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_129),
.Y(n_165)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_92),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_139),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_94),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_45),
.B(n_48),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_148),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_149),
.Y(n_170)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

CKINVDCx6p67_ASAP7_75t_R g183 ( 
.A(n_146),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_126),
.A2(n_32),
.B1(n_67),
.B2(n_86),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_147),
.A2(n_153),
.B1(n_159),
.B2(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_154),
.Y(n_189)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_62),
.B1(n_84),
.B2(n_77),
.Y(n_155)
);

AO22x2_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_128),
.B1(n_63),
.B2(n_66),
.Y(n_178)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_102),
.B(n_109),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_160),
.B(n_168),
.Y(n_175)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_162),
.Y(n_172)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_163),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_108),
.A2(n_31),
.B1(n_32),
.B2(n_48),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_111),
.B(n_106),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_167),
.Y(n_187)
);

INVx6_ASAP7_75t_SL g168 ( 
.A(n_111),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_107),
.C(n_109),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_174),
.B(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_107),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_185),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_131),
.B1(n_121),
.B2(n_119),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_41),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_93),
.C(n_98),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_99),
.C(n_114),
.Y(n_185)
);

CKINVDCx12_ASAP7_75t_R g190 ( 
.A(n_161),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_190),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_137),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_196),
.A2(n_187),
.B1(n_172),
.B2(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_199),
.A2(n_207),
.B(n_208),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_179),
.B1(n_178),
.B2(n_183),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_95),
.B1(n_185),
.B2(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_155),
.B1(n_100),
.B2(n_147),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_205),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_171),
.B(n_51),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_165),
.B(n_139),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_206),
.A2(n_207),
.B(n_199),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_188),
.A2(n_161),
.B1(n_144),
.B2(n_167),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_188),
.A2(n_162),
.B1(n_156),
.B2(n_165),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_212),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_131),
.B1(n_116),
.B2(n_146),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_211),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_45),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_230),
.B1(n_203),
.B2(n_206),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_174),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_220),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_221),
.A2(n_208),
.B(n_202),
.Y(n_239)
);

AO22x1_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_203),
.B1(n_196),
.B2(n_178),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_226),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_186),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_193),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_199),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_187),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_195),
.A2(n_183),
.B1(n_172),
.B2(n_184),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_195),
.B1(n_182),
.B2(n_204),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_181),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_24),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_199),
.B(n_183),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_235),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_202),
.C(n_198),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_43),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_238),
.A2(n_246),
.B1(n_221),
.B2(n_225),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_247),
.B(n_248),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_213),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_242),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_194),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_181),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_249),
.C(n_253),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_244),
.A2(n_215),
.B1(n_214),
.B2(n_235),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_205),
.B1(n_209),
.B2(n_201),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_184),
.B(n_197),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_223),
.B(n_225),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_186),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_134),
.B1(n_182),
.B2(n_101),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_230),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_145),
.C(n_114),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_227),
.Y(n_259)
);

OAI32xp33_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_173),
.A3(n_24),
.B1(n_28),
.B2(n_43),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_258),
.A2(n_266),
.B1(n_250),
.B2(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_270),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_225),
.B1(n_221),
.B2(n_224),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_263),
.A2(n_264),
.B1(n_267),
.B2(n_269),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_238),
.A2(n_214),
.B1(n_217),
.B2(n_219),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_217),
.B1(n_219),
.B2(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_222),
.B1(n_182),
.B2(n_166),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_159),
.B1(n_150),
.B2(n_135),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_130),
.B1(n_119),
.B2(n_59),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_173),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_173),
.Y(n_272)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_236),
.Y(n_278)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_282),
.Y(n_299)
);

BUFx12_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_279),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_280),
.A2(n_292),
.B1(n_296),
.B2(n_132),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_237),
.C(n_246),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_40),
.C(n_39),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_253),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_286),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_265),
.A2(n_250),
.B(n_252),
.C(n_255),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_283),
.A2(n_297),
.B(n_41),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_252),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_256),
.B(n_267),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_261),
.A2(n_130),
.B1(n_25),
.B2(n_35),
.Y(n_296)
);

BUFx12f_ASAP7_75t_SL g297 ( 
.A(n_265),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_258),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_298),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_310),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_274),
.B1(n_262),
.B2(n_271),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_301),
.A2(n_303),
.B1(n_283),
.B2(n_279),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_68),
.B1(n_74),
.B2(n_69),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_309),
.C(n_320),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_305),
.A2(n_283),
.B1(n_279),
.B2(n_25),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_0),
.B(n_1),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_307),
.Y(n_325)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_173),
.C(n_25),
.Y(n_309)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_278),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_2),
.Y(n_313)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_3),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_315),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_4),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_317),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_291),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_318),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_284),
.A2(n_5),
.B(n_6),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_6),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_277),
.B(n_288),
.Y(n_320)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_337),
.Y(n_343)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_312),
.A2(n_321),
.B1(n_300),
.B2(n_306),
.Y(n_328)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_328),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_312),
.B1(n_311),
.B2(n_301),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_307),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_315),
.A2(n_283),
.B1(n_40),
.B2(n_44),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_334),
.B(n_336),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_303),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_317),
.A2(n_44),
.B1(n_40),
.B2(n_37),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_302),
.B(n_44),
.C(n_28),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_338),
.B(n_302),
.C(n_304),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_349),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_341),
.B(n_342),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_326),
.B(n_310),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_324),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_309),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_345),
.B(n_348),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_299),
.C(n_319),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_308),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_28),
.C(n_43),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_323),
.C(n_348),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_354),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_328),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_330),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_356),
.B(n_359),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_347),
.Y(n_357)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_358),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_335),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_360),
.B(n_362),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_334),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_346),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_363),
.B(n_325),
.Y(n_370)
);

A2O1A1Ixp33_ASAP7_75t_SL g365 ( 
.A1(n_362),
.A2(n_325),
.B(n_337),
.C(n_344),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_365),
.B(n_366),
.Y(n_378)
);

NOR2x1_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_332),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_355),
.C(n_354),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_371),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_370),
.B(n_374),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_357),
.A2(n_88),
.B1(n_28),
.B2(n_8),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g374 ( 
.A1(n_359),
.A2(n_6),
.B(n_7),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_373),
.B(n_28),
.C(n_43),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_375),
.A2(n_381),
.B(n_372),
.Y(n_384)
);

MAJx2_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_7),
.C(n_8),
.Y(n_379)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_8),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_382),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_28),
.C(n_43),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_9),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_377),
.C(n_369),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_383),
.B(n_388),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_387),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_378),
.Y(n_387)
);

OAI21x1_ASAP7_75t_L g388 ( 
.A1(n_376),
.A2(n_365),
.B(n_12),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_386),
.A2(n_10),
.B(n_12),
.Y(n_390)
);

MAJx2_ASAP7_75t_L g392 ( 
.A(n_390),
.B(n_385),
.C(n_13),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_392),
.A2(n_393),
.B(n_389),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_391),
.A2(n_12),
.B(n_13),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_394),
.A2(n_13),
.B(n_14),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_395),
.A2(n_14),
.B(n_16),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_396),
.B(n_16),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_397),
.B(n_17),
.Y(n_398)
);


endmodule