module real_aes_18316_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_850, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_850;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g841 ( .A(n_0), .B(n_842), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_1), .A2(n_33), .B1(n_134), .B2(n_157), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_2), .A2(n_9), .B1(n_176), .B2(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g842 ( .A(n_3), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_4), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_5), .A2(n_10), .B1(n_193), .B2(n_196), .Y(n_192) );
OR2x2_ASAP7_75t_L g115 ( .A(n_6), .B(n_29), .Y(n_115) );
BUFx2_ASAP7_75t_L g847 ( .A(n_6), .Y(n_847) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_7), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_8), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_11), .B(n_137), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_12), .A2(n_98), .B1(n_176), .B2(n_177), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_13), .A2(n_30), .B1(n_142), .B2(n_209), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g109 ( .A1(n_14), .A2(n_17), .B1(n_110), .B2(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_14), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_15), .B(n_137), .Y(n_136) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_16), .A2(n_45), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g111 ( .A(n_17), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_18), .B(n_501), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_19), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_20), .A2(n_37), .B1(n_162), .B2(n_163), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_21), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_22), .A2(n_43), .B1(n_163), .B2(n_176), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_23), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_24), .B(n_142), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_25), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_26), .B(n_194), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_27), .B(n_151), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_28), .Y(n_616) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_29), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_31), .A2(n_81), .B1(n_134), .B2(n_232), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_32), .A2(n_36), .B1(n_133), .B2(n_134), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_34), .A2(n_48), .B1(n_176), .B2(n_180), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_35), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_38), .B(n_137), .Y(n_484) );
INVx2_ASAP7_75t_L g806 ( .A(n_39), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_40), .A2(n_51), .B1(n_821), .B2(n_822), .Y(n_820) );
INVx1_ASAP7_75t_L g822 ( .A(n_40), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_41), .B(n_138), .Y(n_496) );
BUFx3_ASAP7_75t_L g114 ( .A(n_42), .Y(n_114) );
INVx1_ASAP7_75t_L g830 ( .A(n_42), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_44), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g544 ( .A(n_46), .B(n_504), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_47), .B(n_210), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_49), .B(n_194), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_50), .B(n_162), .Y(n_620) );
INVx1_ASAP7_75t_L g821 ( .A(n_51), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_52), .A2(n_68), .B1(n_162), .B2(n_180), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_53), .A2(n_71), .B1(n_133), .B2(n_134), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_54), .B(n_529), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_55), .A2(n_235), .B(n_485), .C(n_538), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_56), .A2(n_94), .B1(n_176), .B2(n_196), .Y(n_222) );
INVx1_ASAP7_75t_L g129 ( .A(n_57), .Y(n_129) );
AND2x4_ASAP7_75t_L g148 ( .A(n_58), .B(n_149), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_59), .A2(n_60), .B1(n_163), .B2(n_213), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_61), .B(n_151), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_62), .B(n_504), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_63), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_64), .B(n_163), .Y(n_489) );
INVx1_ASAP7_75t_L g149 ( .A(n_65), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_66), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_67), .B(n_151), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_69), .B(n_134), .Y(n_524) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_70), .B(n_138), .C(n_157), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_72), .B(n_134), .Y(n_551) );
INVx2_ASAP7_75t_L g139 ( .A(n_73), .Y(n_139) );
CKINVDCx14_ASAP7_75t_R g471 ( .A(n_74), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_74), .A2(n_471), .B1(n_820), .B2(n_823), .Y(n_819) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_75), .B(n_199), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_76), .B(n_137), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_77), .B(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_78), .A2(n_95), .B1(n_163), .B2(n_235), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_79), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_80), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_82), .A2(n_89), .B1(n_194), .B2(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g834 ( .A(n_83), .B(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_84), .B(n_137), .Y(n_617) );
NAND2xp33_ASAP7_75t_SL g569 ( .A(n_85), .B(n_143), .Y(n_569) );
OAI32xp33_ASAP7_75t_L g102 ( .A1(n_86), .A2(n_103), .A3(n_810), .B1(n_836), .B2(n_848), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_87), .B(n_178), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_88), .B(n_151), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_90), .Y(n_203) );
INVx1_ASAP7_75t_L g467 ( .A(n_91), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_91), .B(n_829), .Y(n_828) );
NAND2xp33_ASAP7_75t_L g144 ( .A(n_92), .B(n_137), .Y(n_144) );
NAND2xp33_ASAP7_75t_L g552 ( .A(n_93), .B(n_143), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_96), .B(n_504), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_97), .B(n_143), .C(n_199), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_99), .B(n_800), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_100), .B(n_134), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_101), .B(n_194), .Y(n_527) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI22x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_801), .B1(n_807), .B2(n_808), .Y(n_104) );
OAI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_468), .B(n_799), .Y(n_105) );
NAND2xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_116), .Y(n_106) );
NOR2xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_112), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR3xp33_ASAP7_75t_L g807 ( .A(n_109), .B(n_112), .C(n_803), .Y(n_807) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g800 ( .A(n_113), .B(n_466), .Y(n_800) );
NOR2x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx1_ASAP7_75t_L g831 ( .A(n_115), .Y(n_831) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_116), .Y(n_809) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_117), .B(n_463), .Y(n_116) );
NAND2x1p5_ASAP7_75t_L g117 ( .A(n_118), .B(n_407), .Y(n_117) );
NOR3x1_ASAP7_75t_L g118 ( .A(n_119), .B(n_325), .C(n_362), .Y(n_118) );
NAND4xp75_ASAP7_75t_L g119 ( .A(n_120), .B(n_245), .C(n_279), .D(n_309), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI32xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_167), .A3(n_217), .B1(n_226), .B2(n_240), .Y(n_121) );
OR2x2_ASAP7_75t_L g226 ( .A(n_122), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_123), .A2(n_437), .B(n_439), .Y(n_436) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_152), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_124), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g308 ( .A(n_124), .B(n_254), .Y(n_308) );
AND2x2_ASAP7_75t_L g403 ( .A(n_124), .B(n_219), .Y(n_403) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g252 ( .A(n_125), .Y(n_252) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_130), .B(n_150), .Y(n_125) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_126), .A2(n_130), .B(n_150), .Y(n_285) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
INVx4_ASAP7_75t_L g151 ( .A(n_127), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_127), .B(n_166), .Y(n_165) );
BUFx3_ASAP7_75t_L g214 ( .A(n_127), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_127), .B(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_127), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g480 ( .A(n_127), .Y(n_480) );
AND2x4_ASAP7_75t_SL g559 ( .A(n_127), .B(n_490), .Y(n_559) );
INVx1_ASAP7_75t_SL g562 ( .A(n_127), .Y(n_562) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g184 ( .A(n_128), .Y(n_184) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_140), .B(n_146), .Y(n_130) );
O2A1O1Ixp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_136), .C(n_138), .Y(n_131) );
INVx4_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g180 ( .A(n_134), .Y(n_180) );
INVx1_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
OAI22xp33_ASAP7_75t_L g541 ( .A1(n_134), .A2(n_163), .B1(n_542), .B2(n_543), .Y(n_541) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_135), .Y(n_137) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_135), .Y(n_157) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
INVx1_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g195 ( .A(n_135), .Y(n_195) );
INVx1_ASAP7_75t_L g210 ( .A(n_135), .Y(n_210) );
INVx1_ASAP7_75t_L g213 ( .A(n_135), .Y(n_213) );
INVx2_ASAP7_75t_L g233 ( .A(n_135), .Y(n_233) );
INVx1_ASAP7_75t_L g235 ( .A(n_135), .Y(n_235) );
INVx3_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
INVx1_ASAP7_75t_L g501 ( .A(n_137), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_137), .A2(n_565), .B(n_566), .Y(n_564) );
INVx6_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_138), .A2(n_488), .B(n_489), .Y(n_487) );
O2A1O1Ixp5_ASAP7_75t_L g615 ( .A1(n_138), .A2(n_177), .B(n_616), .C(n_617), .Y(n_615) );
BUFx8_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g160 ( .A(n_139), .Y(n_160) );
INVx1_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
INVx1_ASAP7_75t_L g486 ( .A(n_139), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_144), .B(n_145), .Y(n_140) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g162 ( .A(n_143), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g155 ( .A1(n_145), .A2(n_156), .B1(n_158), .B2(n_161), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g174 ( .A1(n_145), .A2(n_158), .B1(n_175), .B2(n_179), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_145), .A2(n_192), .B1(n_197), .B2(n_198), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_145), .A2(n_158), .B1(n_208), .B2(n_211), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_145), .A2(n_198), .B1(n_222), .B2(n_223), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_145), .A2(n_231), .B1(n_234), .B2(n_236), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_145), .A2(n_158), .B1(n_270), .B2(n_271), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_145), .A2(n_158), .B1(n_507), .B2(n_509), .Y(n_506) );
INVx2_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_SL g237 ( .A(n_147), .Y(n_237) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx10_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
BUFx10_ASAP7_75t_L g490 ( .A(n_148), .Y(n_490) );
INVx2_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
INVx2_ASAP7_75t_L g276 ( .A(n_152), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_152), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_153), .Y(n_263) );
INVx1_ASAP7_75t_L g307 ( .A(n_153), .Y(n_307) );
AND2x2_ASAP7_75t_L g351 ( .A(n_153), .B(n_285), .Y(n_351) );
OR2x2_ASAP7_75t_L g405 ( .A(n_153), .B(n_229), .Y(n_405) );
AO31x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .A3(n_164), .B(n_165), .Y(n_153) );
INVx2_ASAP7_75t_L g173 ( .A(n_154), .Y(n_173) );
AO31x2_ASAP7_75t_L g190 ( .A1(n_154), .A2(n_191), .A3(n_200), .B(n_202), .Y(n_190) );
AO31x2_ASAP7_75t_L g206 ( .A1(n_154), .A2(n_207), .A3(n_214), .B(n_215), .Y(n_206) );
AO31x2_ASAP7_75t_L g505 ( .A1(n_154), .A2(n_183), .A3(n_506), .B(n_510), .Y(n_505) );
INVx2_ASAP7_75t_L g529 ( .A(n_157), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_158), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g530 ( .A(n_159), .Y(n_530) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g556 ( .A(n_160), .Y(n_556) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_163), .A2(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g508 ( .A(n_163), .Y(n_508) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_168), .A2(n_331), .B1(n_423), .B2(n_425), .Y(n_422) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_188), .Y(n_168) );
INVx4_ASAP7_75t_L g248 ( .A(n_169), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_169), .A2(n_228), .B1(n_260), .B2(n_262), .Y(n_259) );
OR2x2_ASAP7_75t_L g265 ( .A(n_169), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g384 ( .A(n_169), .B(n_283), .Y(n_384) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g304 ( .A(n_170), .B(n_189), .Y(n_304) );
AND2x2_ASAP7_75t_L g395 ( .A(n_170), .B(n_267), .Y(n_395) );
AND2x2_ASAP7_75t_L g450 ( .A(n_170), .B(n_206), .Y(n_450) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g244 ( .A(n_171), .Y(n_244) );
AND2x4_ASAP7_75t_L g371 ( .A(n_171), .B(n_267), .Y(n_371) );
AO31x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_174), .A3(n_181), .B(n_185), .Y(n_171) );
AO31x2_ASAP7_75t_L g220 ( .A1(n_172), .A2(n_200), .A3(n_221), .B(n_224), .Y(n_220) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp67_ASAP7_75t_SL g535 ( .A(n_173), .B(n_182), .Y(n_535) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_181), .A2(n_237), .A3(n_269), .B(n_272), .Y(n_268) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_SL g202 ( .A(n_183), .B(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_183), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g187 ( .A(n_184), .Y(n_187) );
INVx2_ASAP7_75t_L g201 ( .A(n_184), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_187), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g504 ( .A(n_187), .Y(n_504) );
INVx2_ASAP7_75t_L g531 ( .A(n_187), .Y(n_531) );
NAND2x1_ASAP7_75t_L g247 ( .A(n_188), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_188), .B(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_204), .Y(n_188) );
INVx2_ASAP7_75t_L g242 ( .A(n_189), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_189), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g290 ( .A(n_189), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_189), .B(n_292), .Y(n_317) );
AND2x2_ASAP7_75t_L g320 ( .A(n_189), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g380 ( .A(n_189), .Y(n_380) );
INVx4_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_190), .B(n_205), .Y(n_258) );
BUFx2_ASAP7_75t_L g296 ( .A(n_190), .Y(n_296) );
AND2x2_ASAP7_75t_L g345 ( .A(n_190), .B(n_206), .Y(n_345) );
AND2x2_ASAP7_75t_L g387 ( .A(n_190), .B(n_268), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_190), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g236 ( .A(n_199), .Y(n_236) );
INVx1_ASAP7_75t_L g502 ( .A(n_199), .Y(n_502) );
BUFx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_201), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_206), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g298 ( .A(n_206), .B(n_268), .Y(n_298) );
INVx1_ASAP7_75t_L g321 ( .A(n_206), .Y(n_321) );
INVx2_ASAP7_75t_L g341 ( .A(n_206), .Y(n_341) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_206), .Y(n_386) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AO31x2_ASAP7_75t_L g229 ( .A1(n_214), .A2(n_230), .A3(n_237), .B(n_238), .Y(n_229) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g305 ( .A(n_218), .B(n_306), .Y(n_305) );
NOR2x1p5_ASAP7_75t_L g411 ( .A(n_218), .B(n_405), .Y(n_411) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x4_ASAP7_75t_L g228 ( .A(n_219), .B(n_229), .Y(n_228) );
INVx3_ASAP7_75t_L g261 ( .A(n_219), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_219), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_219), .B(n_337), .Y(n_336) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g253 ( .A(n_220), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g311 ( .A(n_220), .B(n_229), .Y(n_311) );
BUFx2_ASAP7_75t_L g424 ( .A(n_220), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_226), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g462 ( .A(n_226), .Y(n_462) );
INVx2_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g398 ( .A(n_228), .Y(n_398) );
AND2x4_ASAP7_75t_L g421 ( .A(n_228), .B(n_351), .Y(n_421) );
AND2x2_ASAP7_75t_L g445 ( .A(n_228), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
BUFx2_ASAP7_75t_L g278 ( .A(n_229), .Y(n_278) );
INVx1_ASAP7_75t_L g334 ( .A(n_229), .Y(n_334) );
OR2x2_ASAP7_75t_L g456 ( .A(n_229), .B(n_313), .Y(n_456) );
INVx2_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_233), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g557 ( .A(n_235), .Y(n_557) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g302 ( .A(n_242), .Y(n_302) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_243), .Y(n_319) );
INVx1_ASAP7_75t_L g323 ( .A(n_243), .Y(n_323) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g264 ( .A(n_244), .Y(n_264) );
OR2x2_ASAP7_75t_L g301 ( .A(n_244), .B(n_293), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_249), .B(n_255), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_250), .A2(n_344), .B1(n_346), .B2(n_349), .Y(n_343) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
OR2x2_ASAP7_75t_L g389 ( .A(n_252), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g397 ( .A(n_252), .Y(n_397) );
AND2x2_ASAP7_75t_L g410 ( .A(n_252), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g372 ( .A(n_253), .B(n_351), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_259), .B1(n_265), .B2(n_274), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g324 ( .A(n_258), .Y(n_324) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g282 ( .A(n_261), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g350 ( .A(n_261), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g359 ( .A(n_261), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_261), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_262), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g347 ( .A(n_264), .B(n_348), .Y(n_347) );
INVx3_ASAP7_75t_L g361 ( .A(n_264), .Y(n_361) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g293 ( .A(n_268), .Y(n_293) );
AND2x4_ASAP7_75t_L g340 ( .A(n_268), .B(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_268), .Y(n_356) );
INVx1_ASAP7_75t_L g420 ( .A(n_268), .Y(n_420) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
AND2x4_ASAP7_75t_L g312 ( .A(n_276), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
INVx1_ASAP7_75t_L g287 ( .A(n_278), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_288), .B1(n_299), .B2(n_305), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g281 ( .A(n_282), .B(n_286), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_284), .Y(n_337) );
INVx1_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_289), .B(n_294), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_290), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g442 ( .A(n_291), .Y(n_442) );
INVx1_ASAP7_75t_L g461 ( .A(n_291), .Y(n_461) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2x1_ASAP7_75t_L g438 ( .A(n_295), .B(n_361), .Y(n_438) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g454 ( .A(n_296), .Y(n_454) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
INVx2_ASAP7_75t_L g392 ( .A(n_300), .Y(n_392) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx2_ASAP7_75t_L g381 ( .A(n_301), .Y(n_381) );
AND2x4_ASAP7_75t_L g383 ( .A(n_302), .B(n_340), .Y(n_383) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_306), .A2(n_452), .B1(n_455), .B2(n_457), .Y(n_451) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx2_ASAP7_75t_L g376 ( .A(n_307), .Y(n_376) );
INVx1_ASAP7_75t_L g330 ( .A(n_308), .Y(n_330) );
AND2x4_ASAP7_75t_L g423 ( .A(n_308), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g431 ( .A(n_308), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_314), .Y(n_309) );
AND2x4_ASAP7_75t_SL g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_SL g374 ( .A(n_311), .Y(n_374) );
INVx2_ASAP7_75t_L g390 ( .A(n_311), .Y(n_390) );
INVx1_ASAP7_75t_L g417 ( .A(n_312), .Y(n_417) );
AND2x2_ASAP7_75t_L g448 ( .A(n_312), .B(n_359), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .C(n_322), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_319), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g360 ( .A(n_320), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_320), .B(n_395), .Y(n_428) );
INVx1_ASAP7_75t_L g348 ( .A(n_321), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_323), .B(n_387), .Y(n_413) );
INVx1_ASAP7_75t_L g368 ( .A(n_324), .Y(n_368) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_342), .C(n_352), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_331), .B(n_338), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g446 ( .A(n_329), .Y(n_446) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_335), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI32xp33_ASAP7_75t_L g382 ( .A1(n_333), .A2(n_383), .A3(n_384), .B1(n_385), .B2(n_388), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_333), .B(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g366 ( .A(n_340), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g401 ( .A(n_340), .B(n_361), .Y(n_401) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_345), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g406 ( .A(n_345), .B(n_355), .Y(n_406) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g434 ( .A(n_348), .Y(n_434) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_350), .A2(n_353), .B1(n_357), .B2(n_360), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_351), .B(n_359), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_353), .A2(n_411), .B1(n_448), .B2(n_449), .Y(n_447) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g449 ( .A(n_355), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_357), .A2(n_400), .B1(n_402), .B2(n_406), .Y(n_399) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g441 ( .A(n_361), .Y(n_441) );
NAND4xp25_ASAP7_75t_L g362 ( .A(n_363), .B(n_382), .C(n_391), .D(n_399), .Y(n_362) );
O2A1O1Ixp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_369), .B(n_372), .C(n_373), .Y(n_363) );
NOR2x1_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g427 ( .A(n_371), .B(n_386), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_371), .B(n_454), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_378), .A2(n_416), .B1(n_418), .B2(n_421), .Y(n_415) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI21xp5_ASAP7_75t_L g444 ( .A1(n_383), .A2(n_388), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI21xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_396), .Y(n_391) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_R g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_406), .A2(n_423), .B1(n_460), .B2(n_462), .Y(n_459) );
NOR3x1_ASAP7_75t_L g407 ( .A(n_408), .B(n_429), .C(n_443), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_422), .Y(n_408) );
AOI21xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g435 ( .A(n_410), .Y(n_435) );
INVx2_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
INVx1_ASAP7_75t_L g432 ( .A(n_424), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_426), .A2(n_430), .B1(n_433), .B2(n_435), .C(n_436), .Y(n_429) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
NAND4xp25_ASAP7_75t_SL g443 ( .A(n_444), .B(n_447), .C(n_451), .D(n_459), .Y(n_443) );
AND2x2_ASAP7_75t_L g457 ( .A(n_450), .B(n_458), .Y(n_457) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx4_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx12f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g798 ( .A(n_467), .Y(n_798) );
INVx1_ASAP7_75t_L g813 ( .A(n_468), .Y(n_813) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_795), .Y(n_469) );
XNOR2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
BUFx2_ASAP7_75t_L g817 ( .A(n_472), .Y(n_817) );
NAND2x1p5_ASAP7_75t_SL g472 ( .A(n_473), .B(n_729), .Y(n_472) );
NOR2x1_ASAP7_75t_L g473 ( .A(n_474), .B(n_665), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g474 ( .A(n_475), .B(n_587), .C(n_626), .D(n_655), .Y(n_474) );
O2A1O1Ixp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_512), .B(n_519), .C(n_571), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_492), .Y(n_476) );
INVx2_ASAP7_75t_L g515 ( .A(n_477), .Y(n_515) );
AND2x2_ASAP7_75t_L g653 ( .A(n_477), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_477), .B(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_477), .B(n_573), .Y(n_748) );
OR2x2_ASAP7_75t_L g784 ( .A(n_477), .B(n_700), .Y(n_784) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g681 ( .A(n_478), .B(n_493), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g707 ( .A(n_478), .B(n_517), .Y(n_707) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g642 ( .A(n_479), .Y(n_642) );
OAI21x1_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_491), .Y(n_479) );
OAI21x1_ASAP7_75t_L g493 ( .A1(n_480), .A2(n_494), .B(n_503), .Y(n_493) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_480), .A2(n_481), .B(n_491), .Y(n_575) );
OA21x2_ASAP7_75t_L g610 ( .A1(n_480), .A2(n_494), .B(n_503), .Y(n_610) );
OAI21x1_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_487), .B(n_490), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_485), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_485), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_485), .A2(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_485), .A2(n_568), .B(n_569), .Y(n_567) );
BUFx4f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI21x1_ASAP7_75t_L g494 ( .A1(n_490), .A2(n_495), .B(n_498), .Y(n_494) );
OAI21x1_ASAP7_75t_L g522 ( .A1(n_490), .A2(n_523), .B(n_526), .Y(n_522) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_490), .A2(n_564), .B(n_567), .Y(n_563) );
OAI21x1_ASAP7_75t_L g614 ( .A1(n_490), .A2(n_615), .B(n_618), .Y(n_614) );
AND2x2_ASAP7_75t_L g581 ( .A(n_492), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_492), .B(n_611), .Y(n_625) );
AND2x2_ASAP7_75t_L g633 ( .A(n_492), .B(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_492), .Y(n_656) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_505), .Y(n_492) );
INVx1_ASAP7_75t_L g517 ( .A(n_493), .Y(n_517) );
INVx1_ASAP7_75t_L g573 ( .A(n_493), .Y(n_573) );
AND2x2_ASAP7_75t_L g643 ( .A(n_493), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g704 ( .A(n_493), .B(n_612), .Y(n_704) );
AOI21x1_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B(n_502), .Y(n_498) );
INVx1_ASAP7_75t_L g518 ( .A(n_505), .Y(n_518) );
AND2x2_ASAP7_75t_L g574 ( .A(n_505), .B(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_505), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_505), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g687 ( .A(n_505), .B(n_642), .Y(n_687) );
OR2x2_ASAP7_75t_L g700 ( .A(n_505), .B(n_610), .Y(n_700) );
OR2x2_ASAP7_75t_L g710 ( .A(n_505), .B(n_575), .Y(n_710) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_515), .B(n_726), .Y(n_772) );
INVx1_ASAP7_75t_L g628 ( .A(n_516), .Y(n_628) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AND2x2_ASAP7_75t_L g712 ( .A(n_518), .B(n_575), .Y(n_712) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_545), .Y(n_519) );
AND2x2_ASAP7_75t_L g585 ( .A(n_520), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g647 ( .A(n_520), .Y(n_647) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_533), .Y(n_520) );
BUFx2_ASAP7_75t_L g754 ( .A(n_521), .Y(n_754) );
OAI21xp33_ASAP7_75t_SL g521 ( .A1(n_522), .A2(n_531), .B(n_532), .Y(n_521) );
OAI21x1_ASAP7_75t_L g595 ( .A1(n_522), .A2(n_531), .B(n_532), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_530), .Y(n_526) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_531), .A2(n_614), .B(n_621), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g644 ( .A1(n_531), .A2(n_614), .B(n_621), .Y(n_644) );
AND2x2_ASAP7_75t_L g593 ( .A(n_533), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g579 ( .A(n_534), .B(n_561), .Y(n_579) );
INVx2_ASAP7_75t_L g605 ( .A(n_534), .Y(n_605) );
AOI21x1_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B(n_544), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
AND2x2_ASAP7_75t_L g751 ( .A(n_545), .B(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_560), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g578 ( .A(n_547), .Y(n_578) );
BUFx2_ASAP7_75t_L g586 ( .A(n_547), .Y(n_586) );
OR2x2_ASAP7_75t_L g590 ( .A(n_547), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g650 ( .A(n_547), .B(n_594), .Y(n_650) );
AND2x4_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
OAI21x1_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_553), .B(n_559), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_556), .B1(n_557), .B2(n_558), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_555), .A2(n_619), .B(n_620), .Y(n_618) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g637 ( .A(n_560), .Y(n_637) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_560), .Y(n_651) );
INVx2_ASAP7_75t_L g676 ( .A(n_560), .Y(n_676) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g591 ( .A(n_561), .Y(n_591) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B(n_570), .Y(n_561) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B1(n_580), .B2(n_584), .Y(n_571) );
INVx1_ASAP7_75t_L g661 ( .A(n_572), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx2_ASAP7_75t_L g672 ( .A(n_573), .Y(n_672) );
AND2x2_ASAP7_75t_L g689 ( .A(n_574), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_574), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g583 ( .A(n_575), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_576), .B(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_577), .B(n_593), .Y(n_684) );
AND2x2_ASAP7_75t_L g692 ( .A(n_577), .B(n_658), .Y(n_692) );
AND2x2_ASAP7_75t_L g768 ( .A(n_577), .B(n_715), .Y(n_768) );
BUFx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g603 ( .A(n_578), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g624 ( .A(n_578), .B(n_594), .Y(n_624) );
OR2x2_ASAP7_75t_L g636 ( .A(n_578), .B(n_637), .Y(n_636) );
NAND2x1_ASAP7_75t_L g670 ( .A(n_578), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g675 ( .A(n_578), .Y(n_675) );
INVx2_ASAP7_75t_L g669 ( .A(n_579), .Y(n_669) );
AND2x2_ASAP7_75t_L g695 ( .A(n_579), .B(n_659), .Y(n_695) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_582), .Y(n_631) );
INVx1_ASAP7_75t_L g698 ( .A(n_582), .Y(n_698) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g682 ( .A(n_583), .B(n_612), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g693 ( .A1(n_584), .A2(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_L g755 ( .A(n_586), .B(n_695), .Y(n_755) );
INVx1_ASAP7_75t_L g791 ( .A(n_586), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_596), .B(n_600), .Y(n_587) );
AOI322xp5_ASAP7_75t_L g739 ( .A1(n_588), .A2(n_635), .A3(n_740), .B1(n_741), .B2(n_742), .C1(n_743), .C2(n_746), .Y(n_739) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g727 ( .A(n_590), .B(n_592), .C(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g606 ( .A(n_591), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g735 ( .A(n_591), .B(n_736), .Y(n_735) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_591), .Y(n_787) );
OR2x2_ASAP7_75t_L g683 ( .A(n_592), .B(n_636), .Y(n_683) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g671 ( .A(n_594), .Y(n_671) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g607 ( .A(n_595), .Y(n_607) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVxp67_ASAP7_75t_SL g732 ( .A(n_597), .Y(n_732) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g703 ( .A(n_598), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g766 ( .A(n_599), .B(n_726), .Y(n_766) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_608), .B(n_622), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_602), .B(n_780), .Y(n_779) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .Y(n_602) );
AND2x2_ASAP7_75t_L g658 ( .A(n_604), .B(n_659), .Y(n_658) );
AND3x2_ASAP7_75t_L g702 ( .A(n_604), .B(n_606), .C(n_675), .Y(n_702) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g664 ( .A(n_605), .Y(n_664) );
AND2x2_ASAP7_75t_L g715 ( .A(n_605), .B(n_676), .Y(n_715) );
INVx2_ASAP7_75t_L g738 ( .A(n_605), .Y(n_738) );
AND2x2_ASAP7_75t_L g742 ( .A(n_606), .B(n_738), .Y(n_742) );
INVx2_ASAP7_75t_L g659 ( .A(n_607), .Y(n_659) );
OR2x2_ASAP7_75t_L g793 ( .A(n_607), .B(n_676), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_608), .B(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g745 ( .A(n_609), .Y(n_745) );
AND2x2_ASAP7_75t_L g654 ( .A(n_610), .B(n_644), .Y(n_654) );
AND2x2_ASAP7_75t_L g690 ( .A(n_610), .B(n_612), .Y(n_690) );
AND2x2_ASAP7_75t_L g686 ( .A(n_611), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_611), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g758 ( .A(n_611), .Y(n_758) );
BUFx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g629 ( .A(n_612), .Y(n_629) );
INVxp67_ASAP7_75t_SL g634 ( .A(n_612), .Y(n_634) );
INVxp67_ASAP7_75t_SL g680 ( .A(n_612), .Y(n_680) );
INVx1_ASAP7_75t_L g726 ( .A(n_612), .Y(n_726) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_635), .B(n_638), .Y(n_626) );
OAI31xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .A3(n_630), .B(n_632), .Y(n_627) );
INVx1_ASAP7_75t_L g709 ( .A(n_629), .Y(n_709) );
OAI32xp33_ASAP7_75t_L g667 ( .A1(n_630), .A2(n_639), .A3(n_668), .B1(n_672), .B2(n_673), .Y(n_667) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g660 ( .A(n_636), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_645), .B1(n_648), .B2(n_652), .Y(n_638) );
OAI22xp33_ASAP7_75t_SL g723 ( .A1(n_639), .A2(n_684), .B1(n_724), .B2(n_725), .Y(n_723) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx2_ASAP7_75t_L g781 ( .A(n_641), .Y(n_781) );
BUFx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g736 ( .A(n_644), .Y(n_736) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
AND2x2_ASAP7_75t_L g662 ( .A(n_650), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g737 ( .A(n_650), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g788 ( .A(n_650), .Y(n_788) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g728 ( .A(n_654), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_661), .B2(n_662), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_657), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
AND2x2_ASAP7_75t_L g714 ( .A(n_659), .B(n_675), .Y(n_714) );
AOI211xp5_ASAP7_75t_L g719 ( .A1(n_662), .A2(n_720), .B(n_723), .C(n_727), .Y(n_719) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_664), .Y(n_777) );
INVx1_ASAP7_75t_L g794 ( .A(n_664), .Y(n_794) );
NAND4xp25_ASAP7_75t_L g665 ( .A(n_666), .B(n_688), .C(n_701), .D(n_719), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_677), .Y(n_666) );
OR2x6_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_671), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g776 ( .A(n_674), .B(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_677) );
NOR2xp33_ASAP7_75t_SL g678 ( .A(n_679), .B(n_682), .Y(n_678) );
BUFx2_ASAP7_75t_L g691 ( .A(n_679), .Y(n_691) );
AND2x4_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_685), .B(n_771), .Y(n_770) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g740 ( .A(n_687), .B(n_726), .Y(n_740) );
O2A1O1Ixp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_692), .C(n_693), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_690), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g750 ( .A(n_697), .B(n_751), .Y(n_750) );
AND2x4_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_705), .B2(n_713), .C(n_716), .Y(n_701) );
AND2x2_ASAP7_75t_L g780 ( .A(n_704), .B(n_781), .Y(n_780) );
NAND3xp33_ASAP7_75t_SL g705 ( .A(n_706), .B(n_708), .C(n_711), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_709), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_709), .B(n_745), .Y(n_775) );
INVx1_ASAP7_75t_L g718 ( .A(n_710), .Y(n_718) );
INVx1_ASAP7_75t_L g722 ( .A(n_710), .Y(n_722) );
AND2x2_ASAP7_75t_L g763 ( .A(n_712), .B(n_752), .Y(n_763) );
NAND2xp33_ASAP7_75t_SL g764 ( .A(n_712), .B(n_734), .Y(n_764) );
AND2x4_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g724 ( .A(n_715), .Y(n_724) );
NOR3x1_ASAP7_75t_L g729 ( .A(n_730), .B(n_759), .C(n_778), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_739), .C(n_749), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g752 ( .A(n_736), .Y(n_752) );
INVx2_ASAP7_75t_L g741 ( .A(n_738), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_740), .A2(n_783), .B1(n_790), .B2(n_850), .Y(n_789) );
O2A1O1Ixp5_ASAP7_75t_L g761 ( .A1(n_741), .A2(n_753), .B(n_762), .C(n_764), .Y(n_761) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AO21x1_ASAP7_75t_L g765 ( .A1(n_744), .A2(n_766), .B(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g757 ( .A(n_748), .B(n_758), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_753), .B1(n_755), .B2(n_756), .Y(n_749) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND4xp75_ASAP7_75t_L g759 ( .A(n_760), .B(n_765), .C(n_769), .D(n_773), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND3xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_782), .C(n_789), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_785), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVxp67_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
AND2x4_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
NOR2x1p5_ASAP7_75t_SL g792 ( .A(n_793), .B(n_794), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_798), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_803), .A2(n_815), .B(n_834), .Y(n_814) );
CKINVDCx11_ASAP7_75t_R g803 ( .A(n_804), .Y(n_803) );
BUFx6f_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx3_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g812 ( .A(n_807), .Y(n_812) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OA21x2_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_813), .B(n_814), .Y(n_811) );
OAI22xp5_ASAP7_75t_SL g815 ( .A1(n_816), .A2(n_817), .B1(n_818), .B2(n_832), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_824), .Y(n_818) );
INVx1_ASAP7_75t_L g833 ( .A(n_819), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_820), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_824), .B(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
BUFx2_ASAP7_75t_L g835 ( .A(n_827), .Y(n_835) );
AND2x6_ASAP7_75t_SL g827 ( .A(n_828), .B(n_831), .Y(n_827) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_830), .Y(n_839) );
INVx3_ASAP7_75t_SL g848 ( .A(n_836), .Y(n_848) );
OR2x6_ASAP7_75t_L g836 ( .A(n_837), .B(n_843), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NOR2x1p5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NOR2x1p5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
endmodule