module real_aes_441_n_239 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_239);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_239;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_397;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_623;
wire n_249;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_0), .A2(n_209), .B1(n_381), .B2(n_422), .Y(n_435) );
AO222x2_ASAP7_75t_SL g669 ( .A1(n_1), .A2(n_30), .B1(n_145), .B2(n_416), .C1(n_506), .C2(n_670), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_2), .A2(n_222), .B1(n_318), .B2(n_322), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_3), .A2(n_126), .B1(n_380), .B2(n_381), .Y(n_453) );
AO22x2_ASAP7_75t_L g267 ( .A1(n_4), .A2(n_166), .B1(n_257), .B2(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g650 ( .A(n_4), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_5), .A2(n_25), .B1(n_277), .B2(n_501), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_6), .A2(n_117), .B1(n_377), .B2(n_378), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_7), .A2(n_694), .B1(n_695), .B2(n_696), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_7), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_8), .A2(n_206), .B1(n_318), .B2(n_322), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_9), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_10), .A2(n_56), .B1(n_508), .B2(n_510), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_11), .A2(n_93), .B1(n_300), .B2(n_506), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_12), .A2(n_59), .B1(n_394), .B2(n_395), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_13), .A2(n_152), .B1(n_308), .B2(n_443), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_14), .A2(n_171), .B1(n_354), .B2(n_355), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_15), .A2(n_78), .B1(n_278), .B2(n_418), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_16), .A2(n_86), .B1(n_392), .B2(n_395), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_17), .A2(n_36), .B1(n_481), .B2(n_635), .Y(n_634) );
AO22x2_ASAP7_75t_L g264 ( .A1(n_18), .A2(n_58), .B1(n_257), .B2(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_18), .B(n_649), .Y(n_648) );
XOR2xp5_ASAP7_75t_SL g622 ( .A(n_19), .B(n_623), .Y(n_622) );
XOR2x2_ASAP7_75t_L g639 ( .A(n_19), .B(n_624), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_20), .A2(n_43), .B1(n_391), .B2(n_392), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_21), .A2(n_155), .B1(n_304), .B2(n_307), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_22), .A2(n_40), .B1(n_283), .B2(n_287), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_23), .A2(n_128), .B1(n_413), .B2(n_440), .Y(n_439) );
AO222x2_ASAP7_75t_SL g472 ( .A1(n_24), .A2(n_143), .B1(n_229), .B2(n_251), .C1(n_344), .C2(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_26), .A2(n_55), .B1(n_307), .B2(n_357), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_27), .A2(n_131), .B1(n_523), .B2(n_607), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_28), .A2(n_47), .B1(n_271), .B2(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_29), .A2(n_76), .B1(n_443), .B2(n_444), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_31), .A2(n_185), .B1(n_354), .B2(n_355), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_32), .A2(n_237), .B1(n_392), .B2(n_395), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_33), .A2(n_230), .B1(n_484), .B2(n_607), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_34), .A2(n_217), .B1(n_318), .B2(n_322), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_35), .A2(n_150), .B1(n_346), .B2(n_347), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_37), .A2(n_170), .B1(n_395), .B2(n_413), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_38), .A2(n_227), .B1(n_327), .B2(n_331), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_39), .A2(n_179), .B1(n_349), .B2(n_504), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_41), .A2(n_140), .B1(n_613), .B2(n_614), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_42), .A2(n_95), .B1(n_359), .B2(n_360), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_44), .B(n_375), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_45), .A2(n_178), .B1(n_563), .B2(n_564), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_46), .A2(n_233), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_48), .A2(n_79), .B1(n_270), .B2(n_277), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_49), .A2(n_188), .B1(n_471), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_50), .A2(n_187), .B1(n_389), .B2(n_394), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_51), .A2(n_142), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_52), .A2(n_62), .B1(n_324), .B2(n_480), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_53), .A2(n_183), .B1(n_333), .B2(n_392), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_54), .A2(n_91), .B1(n_508), .B2(n_510), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_57), .A2(n_107), .B1(n_380), .B2(n_381), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_60), .A2(n_138), .B1(n_509), .B2(n_537), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_61), .A2(n_90), .B1(n_477), .B2(n_478), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_63), .A2(n_223), .B1(n_383), .B2(n_384), .Y(n_382) );
XNOR2x2_ASAP7_75t_L g574 ( .A(n_64), .B(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_65), .A2(n_176), .B1(n_294), .B2(n_535), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_66), .B(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_67), .A2(n_151), .B1(n_389), .B2(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_68), .A2(n_204), .B1(n_440), .B2(n_541), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_69), .A2(n_119), .B1(n_604), .B2(n_605), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_70), .A2(n_96), .B1(n_349), .B2(n_350), .Y(n_348) );
INVx3_ASAP7_75t_L g257 ( .A(n_71), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_72), .A2(n_235), .B1(n_418), .B2(n_468), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_73), .A2(n_146), .B1(n_271), .B2(n_350), .Y(n_533) );
AO22x2_ASAP7_75t_L g530 ( .A1(n_74), .A2(n_531), .B1(n_545), .B2(n_546), .Y(n_530) );
INVx1_ASAP7_75t_L g545 ( .A(n_74), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_75), .A2(n_213), .B1(n_487), .B2(n_488), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_77), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_80), .A2(n_97), .B1(n_347), .B2(n_613), .Y(n_631) );
XOR2x2_ASAP7_75t_L g448 ( .A(n_81), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_82), .B(n_512), .Y(n_511) );
OA22x2_ASAP7_75t_L g597 ( .A1(n_83), .A2(n_598), .B1(n_599), .B2(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_83), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_84), .A2(n_186), .B1(n_383), .B2(n_384), .Y(n_452) );
AO22x1_ASAP7_75t_L g577 ( .A1(n_85), .A2(n_139), .B1(n_468), .B2(n_578), .Y(n_577) );
INVx1_ASAP7_75t_SL g258 ( .A(n_87), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_87), .B(n_116), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_88), .A2(n_111), .B1(n_604), .B2(n_605), .Y(n_603) );
AOI222xp33_ASAP7_75t_L g637 ( .A1(n_89), .A2(n_100), .B1(n_212), .B2(n_342), .C1(n_508), .C2(n_510), .Y(n_637) );
INVx2_ASAP7_75t_L g658 ( .A(n_92), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_94), .A2(n_203), .B1(n_284), .B2(n_344), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_98), .A2(n_189), .B1(n_304), .B2(n_594), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_99), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_101), .A2(n_114), .B1(n_391), .B2(n_408), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_102), .A2(n_122), .B1(n_501), .B2(n_503), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_103), .A2(n_113), .B1(n_395), .B2(n_519), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_104), .A2(n_193), .B1(n_307), .B2(n_357), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_105), .A2(n_238), .B1(n_443), .B2(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_106), .A2(n_124), .B1(n_523), .B2(n_525), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_108), .A2(n_220), .B1(n_377), .B2(n_378), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_109), .B(n_250), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_110), .A2(n_199), .B1(n_318), .B2(n_687), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_112), .A2(n_205), .B1(n_388), .B2(n_389), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_115), .B(n_375), .Y(n_374) );
AO22x2_ASAP7_75t_L g260 ( .A1(n_116), .A2(n_174), .B1(n_257), .B2(n_261), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_118), .A2(n_172), .B1(n_284), .B2(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_120), .A2(n_226), .B1(n_347), .B2(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_121), .B(n_416), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_123), .A2(n_148), .B1(n_346), .B2(n_535), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_125), .A2(n_197), .B1(n_383), .B2(n_384), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_127), .A2(n_141), .B1(n_480), .B2(n_481), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_129), .B(n_416), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_130), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_132), .A2(n_214), .B1(n_311), .B2(n_314), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_133), .Y(n_431) );
INVx1_ASAP7_75t_L g259 ( .A(n_134), .Y(n_259) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_135), .A2(n_182), .B1(n_355), .B2(n_410), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_136), .A2(n_158), .B1(n_508), .B2(n_510), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_137), .A2(n_156), .B1(n_440), .B2(n_541), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_144), .A2(n_163), .B1(n_354), .B2(n_355), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_147), .A2(n_232), .B1(n_410), .B2(n_411), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_149), .A2(n_231), .B1(n_377), .B2(n_378), .Y(n_434) );
AO22x2_ASAP7_75t_L g464 ( .A1(n_153), .A2(n_465), .B1(n_489), .B2(n_490), .Y(n_464) );
INVx1_ASAP7_75t_L g490 ( .A(n_153), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_154), .A2(n_198), .B1(n_517), .B2(n_520), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_157), .A2(n_218), .B1(n_617), .B2(n_619), .Y(n_616) );
XNOR2x1_ASAP7_75t_L g371 ( .A(n_159), .B(n_372), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_160), .A2(n_177), .B1(n_314), .B2(n_363), .Y(n_362) );
AO22x1_ASAP7_75t_L g579 ( .A1(n_161), .A2(n_225), .B1(n_537), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_162), .A2(n_190), .B1(n_487), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_164), .A2(n_180), .B1(n_487), .B2(n_488), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_165), .A2(n_194), .B1(n_566), .B2(n_567), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_167), .A2(n_211), .B1(n_294), .B2(n_298), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_168), .A2(n_224), .B1(n_481), .B2(n_563), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_169), .A2(n_208), .B1(n_587), .B2(n_588), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_173), .B(n_512), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_175), .A2(n_184), .B1(n_485), .B2(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_181), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g664 ( .A(n_191), .Y(n_664) );
AO21x2_ASAP7_75t_L g666 ( .A1(n_191), .A2(n_667), .B(n_688), .Y(n_666) );
XOR2x2_ASAP7_75t_L g497 ( .A(n_192), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g645 ( .A(n_195), .Y(n_645) );
AND2x4_ASAP7_75t_L g660 ( .A(n_195), .B(n_646), .Y(n_660) );
AO21x1_ASAP7_75t_L g662 ( .A1(n_195), .A2(n_656), .B(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_196), .A2(n_228), .B1(n_284), .B2(n_344), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_200), .A2(n_210), .B1(n_359), .B2(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g646 ( .A(n_201), .Y(n_646) );
AND2x2_ASAP7_75t_R g698 ( .A(n_201), .B(n_645), .Y(n_698) );
AO21x1_ASAP7_75t_SL g652 ( .A1(n_202), .A2(n_653), .B(n_661), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_207), .A2(n_246), .B1(n_247), .B2(n_334), .Y(n_245) );
INVx1_ASAP7_75t_L g334 ( .A(n_207), .Y(n_334) );
INVxp67_ASAP7_75t_L g657 ( .A(n_215), .Y(n_657) );
XNOR2x1_ASAP7_75t_L g338 ( .A(n_216), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g446 ( .A(n_219), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_221), .A2(n_236), .B1(n_422), .B2(n_423), .Y(n_421) );
OA22x2_ASAP7_75t_L g401 ( .A1(n_234), .A2(n_402), .B1(n_403), .B2(n_424), .Y(n_401) );
INVx1_ASAP7_75t_L g424 ( .A(n_234), .Y(n_424) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_492), .B(n_641), .C(n_652), .Y(n_239) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_240), .A2(n_492), .B(n_642), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B1(n_365), .B2(n_366), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_335), .B1(n_336), .B2(n_364), .Y(n_242) );
INVx1_ASAP7_75t_L g364 ( .A(n_243), .Y(n_364) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
BUFx2_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_302), .Y(n_247) );
NAND4xp25_ASAP7_75t_SL g248 ( .A(n_249), .B(n_269), .C(n_282), .D(n_293), .Y(n_248) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx4_ASAP7_75t_SL g342 ( .A(n_252), .Y(n_342) );
INVx3_ASAP7_75t_L g416 ( .A(n_252), .Y(n_416) );
INVx3_ASAP7_75t_SL g514 ( .A(n_252), .Y(n_514) );
INVx4_ASAP7_75t_SL g584 ( .A(n_252), .Y(n_584) );
INVx6_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_262), .Y(n_253) );
AND2x4_ASAP7_75t_L g279 ( .A(n_254), .B(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g300 ( .A(n_254), .B(n_301), .Y(n_300) );
AND2x4_ASAP7_75t_L g375 ( .A(n_254), .B(n_262), .Y(n_375) );
AND2x2_ASAP7_75t_L g378 ( .A(n_254), .B(n_280), .Y(n_378) );
AND2x2_ASAP7_75t_L g381 ( .A(n_254), .B(n_301), .Y(n_381) );
AND2x2_ASAP7_75t_L g423 ( .A(n_254), .B(n_301), .Y(n_423) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_260), .Y(n_254) );
AND2x2_ASAP7_75t_L g275 ( .A(n_255), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_255), .Y(n_292) );
INVx2_ASAP7_75t_L g297 ( .A(n_255), .Y(n_297) );
OAI22x1_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B1(n_258), .B2(n_259), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g261 ( .A(n_257), .Y(n_261) );
INVx2_ASAP7_75t_L g265 ( .A(n_257), .Y(n_265) );
INVx1_ASAP7_75t_L g268 ( .A(n_257), .Y(n_268) );
INVx2_ASAP7_75t_L g276 ( .A(n_260), .Y(n_276) );
AND2x2_ASAP7_75t_L g296 ( .A(n_260), .B(n_297), .Y(n_296) );
BUFx2_ASAP7_75t_L g325 ( .A(n_260), .Y(n_325) );
AND2x4_ASAP7_75t_L g306 ( .A(n_262), .B(n_275), .Y(n_306) );
AND2x4_ASAP7_75t_L g313 ( .A(n_262), .B(n_309), .Y(n_313) );
AND2x2_ASAP7_75t_L g330 ( .A(n_262), .B(n_296), .Y(n_330) );
AND2x2_ASAP7_75t_L g388 ( .A(n_262), .B(n_275), .Y(n_388) );
AND2x6_ASAP7_75t_L g392 ( .A(n_262), .B(n_296), .Y(n_392) );
AND2x2_ASAP7_75t_L g394 ( .A(n_262), .B(n_309), .Y(n_394) );
AND2x2_ASAP7_75t_L g408 ( .A(n_262), .B(n_275), .Y(n_408) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g274 ( .A(n_264), .Y(n_274) );
AND2x4_ASAP7_75t_L g286 ( .A(n_264), .B(n_266), .Y(n_286) );
AND2x2_ASAP7_75t_L g291 ( .A(n_264), .B(n_267), .Y(n_291) );
INVxp67_ASAP7_75t_L g301 ( .A(n_266), .Y(n_301) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g273 ( .A(n_267), .B(n_274), .Y(n_273) );
BUFx6f_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_272), .Y(n_349) );
INVx3_ASAP7_75t_L g419 ( .A(n_272), .Y(n_419) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
AND2x4_ASAP7_75t_L g316 ( .A(n_273), .B(n_309), .Y(n_316) );
AND2x2_ASAP7_75t_L g321 ( .A(n_273), .B(n_296), .Y(n_321) );
AND2x2_ASAP7_75t_L g354 ( .A(n_273), .B(n_296), .Y(n_354) );
AND2x4_ASAP7_75t_L g377 ( .A(n_273), .B(n_275), .Y(n_377) );
AND2x6_ASAP7_75t_L g395 ( .A(n_273), .B(n_309), .Y(n_395) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_274), .Y(n_281) );
AND2x2_ASAP7_75t_L g285 ( .A(n_275), .B(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g383 ( .A(n_275), .B(n_286), .Y(n_383) );
AND2x4_ASAP7_75t_L g309 ( .A(n_276), .B(n_297), .Y(n_309) );
BUFx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
BUFx6f_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g351 ( .A(n_279), .Y(n_351) );
INVx2_ASAP7_75t_L g469 ( .A(n_279), .Y(n_469) );
BUFx3_ASAP7_75t_L g504 ( .A(n_279), .Y(n_504) );
BUFx4f_ASAP7_75t_L g630 ( .A(n_279), .Y(n_630) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g474 ( .A(n_285), .Y(n_474) );
BUFx3_ASAP7_75t_L g509 ( .A(n_285), .Y(n_509) );
AND2x4_ASAP7_75t_L g295 ( .A(n_286), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g333 ( .A(n_286), .B(n_309), .Y(n_333) );
AND2x2_ASAP7_75t_L g380 ( .A(n_286), .B(n_296), .Y(n_380) );
AND2x2_ASAP7_75t_L g391 ( .A(n_286), .B(n_309), .Y(n_391) );
AND2x2_ASAP7_75t_L g422 ( .A(n_286), .B(n_296), .Y(n_422) );
BUFx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g344 ( .A(n_289), .Y(n_344) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx12f_ASAP7_75t_L g537 ( .A(n_290), .Y(n_537) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x4_ASAP7_75t_L g308 ( .A(n_291), .B(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g324 ( .A(n_291), .B(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g355 ( .A(n_291), .B(n_325), .Y(n_355) );
AND2x2_ASAP7_75t_SL g384 ( .A(n_291), .B(n_292), .Y(n_384) );
AND2x4_ASAP7_75t_L g389 ( .A(n_291), .B(n_309), .Y(n_389) );
BUFx2_ASAP7_75t_L g506 ( .A(n_294), .Y(n_506) );
BUFx4f_ASAP7_75t_SL g613 ( .A(n_294), .Y(n_613) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_L g346 ( .A(n_295), .Y(n_346) );
BUFx3_ASAP7_75t_L g471 ( .A(n_295), .Y(n_471) );
INVx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_SL g347 ( .A(n_299), .Y(n_347) );
INVx2_ASAP7_75t_L g535 ( .A(n_299), .Y(n_535) );
INVx2_ASAP7_75t_L g614 ( .A(n_299), .Y(n_614) );
INVx2_ASAP7_75t_L g670 ( .A(n_299), .Y(n_670) );
INVx6_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND4xp25_ASAP7_75t_L g302 ( .A(n_303), .B(n_310), .C(n_317), .D(n_326), .Y(n_302) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g477 ( .A(n_305), .Y(n_477) );
INVx1_ASAP7_75t_SL g528 ( .A(n_305), .Y(n_528) );
INVx2_ASAP7_75t_L g604 ( .A(n_305), .Y(n_604) );
INVx6_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g357 ( .A(n_306), .Y(n_357) );
BUFx3_ASAP7_75t_L g443 ( .A(n_306), .Y(n_443) );
BUFx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx3_ASAP7_75t_L g444 ( .A(n_308), .Y(n_444) );
BUFx2_ASAP7_75t_SL g485 ( .A(n_308), .Y(n_485) );
INVx2_ASAP7_75t_L g595 ( .A(n_308), .Y(n_595) );
BUFx2_ASAP7_75t_SL g605 ( .A(n_308), .Y(n_605) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_311), .Y(n_484) );
INVx2_ASAP7_75t_L g524 ( .A(n_311), .Y(n_524) );
INVx4_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx3_ASAP7_75t_L g363 ( .A(n_312), .Y(n_363) );
INVx3_ASAP7_75t_SL g413 ( .A(n_312), .Y(n_413) );
INVx2_ASAP7_75t_L g541 ( .A(n_312), .Y(n_541) );
INVx2_ASAP7_75t_SL g590 ( .A(n_312), .Y(n_590) );
INVx8_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_SL g488 ( .A(n_315), .Y(n_488) );
INVx2_ASAP7_75t_L g520 ( .A(n_315), .Y(n_520) );
INVx2_ASAP7_75t_L g567 ( .A(n_315), .Y(n_567) );
INVx2_ASAP7_75t_L g588 ( .A(n_315), .Y(n_588) );
INVx2_ASAP7_75t_L g609 ( .A(n_315), .Y(n_609) );
INVx2_ASAP7_75t_SL g685 ( .A(n_315), .Y(n_685) );
INVx8_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g563 ( .A(n_320), .Y(n_563) );
INVx2_ASAP7_75t_L g636 ( .A(n_320), .Y(n_636) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx3_ASAP7_75t_L g410 ( .A(n_321), .Y(n_410) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_321), .Y(n_480) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx3_ASAP7_75t_L g481 ( .A(n_323), .Y(n_481) );
INVx2_ASAP7_75t_L g564 ( .A(n_323), .Y(n_564) );
INVx2_ASAP7_75t_L g687 ( .A(n_323), .Y(n_687) );
INVx5_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
BUFx2_ASAP7_75t_L g411 ( .A(n_324), .Y(n_411) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx3_ASAP7_75t_L g359 ( .A(n_329), .Y(n_359) );
INVx2_ASAP7_75t_SL g487 ( .A(n_329), .Y(n_487) );
INVx2_ASAP7_75t_L g587 ( .A(n_329), .Y(n_587) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx2_ASAP7_75t_L g519 ( .A(n_330), .Y(n_519) );
BUFx2_ASAP7_75t_L g566 ( .A(n_330), .Y(n_566) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g361 ( .A(n_333), .Y(n_361) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_333), .Y(n_440) );
BUFx3_ASAP7_75t_L g591 ( .A(n_333), .Y(n_591) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_352), .Y(n_339) );
NAND4xp25_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .C(n_345), .D(n_348), .Y(n_340) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_344), .Y(n_510) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NAND4xp25_ASAP7_75t_L g352 ( .A(n_353), .B(n_356), .C(n_358), .D(n_362), .Y(n_352) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g478 ( .A(n_361), .Y(n_478) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
XNOR2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_396), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_385), .Y(n_372) );
NAND4xp25_ASAP7_75t_SL g373 ( .A(n_374), .B(n_376), .C(n_379), .D(n_382), .Y(n_373) );
INVx2_ASAP7_75t_SL g430 ( .A(n_375), .Y(n_430) );
NAND4xp25_ASAP7_75t_SL g385 ( .A(n_386), .B(n_387), .C(n_390), .D(n_393), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B1(n_463), .B2(n_491), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_425), .B1(n_461), .B2(n_462), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g462 ( .A(n_401), .Y(n_462) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR2xp67_ASAP7_75t_L g403 ( .A(n_404), .B(n_414), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_409), .C(n_412), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .C(n_420), .D(n_421), .Y(n_414) );
INVx2_ASAP7_75t_SL g618 ( .A(n_418), .Y(n_618) );
INVx4_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g502 ( .A(n_419), .Y(n_502) );
INVx2_ASAP7_75t_L g578 ( .A(n_419), .Y(n_578) );
INVx2_ASAP7_75t_L g461 ( .A(n_425), .Y(n_461) );
OA22x2_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_447), .B1(n_448), .B2(n_460), .Y(n_425) );
INVx1_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
XOR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_446), .Y(n_426) );
NAND2x1_ASAP7_75t_L g427 ( .A(n_428), .B(n_436), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_433), .Y(n_428) );
OAI21xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_431), .B(n_432), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_441), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx2_ASAP7_75t_L g526 ( .A(n_440), .Y(n_526) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_440), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_445), .Y(n_441) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_444), .Y(n_682) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_455), .Y(n_449) );
NAND4xp25_ASAP7_75t_SL g450 ( .A(n_451), .B(n_452), .C(n_453), .D(n_454), .Y(n_450) );
NAND4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .C(n_458), .D(n_459), .Y(n_455) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_SL g491 ( .A(n_464), .Y(n_491) );
INVx1_ASAP7_75t_SL g489 ( .A(n_465), .Y(n_489) );
NOR4xp75_ASAP7_75t_L g465 ( .A(n_466), .B(n_472), .C(n_475), .D(n_482), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .Y(n_466) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g620 ( .A(n_469), .Y(n_620) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g580 ( .A(n_474), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_479), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_486), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_622), .B1(n_638), .B2(n_640), .Y(n_492) );
INVx1_ASAP7_75t_L g640 ( .A(n_493), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_548), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_497), .B1(n_529), .B2(n_547), .Y(n_495) );
INVx4_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NOR2x1_ASAP7_75t_L g498 ( .A(n_499), .B(n_515), .Y(n_498) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_500), .B(n_505), .C(n_507), .D(n_511), .Y(n_499) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx6f_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
BUFx6f_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI21xp33_ASAP7_75t_SL g554 ( .A1(n_513), .A2(n_555), .B(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND4xp25_ASAP7_75t_L g515 ( .A(n_516), .B(n_521), .C(n_522), .D(n_527), .Y(n_515) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_SL g547 ( .A(n_529), .Y(n_547) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g546 ( .A(n_531), .Y(n_546) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_532), .B(n_539), .Y(n_531) );
NAND4xp25_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .C(n_536), .D(n_538), .Y(n_532) );
NAND4xp25_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .C(n_543), .D(n_544), .Y(n_539) );
INVx1_ASAP7_75t_L g676 ( .A(n_541), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_596), .B1(n_597), .B2(n_621), .Y(n_548) );
INVx1_ASAP7_75t_L g621 ( .A(n_549), .Y(n_621) );
OAI22xp5_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_551), .B1(n_572), .B2(n_573), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
XNOR2x1_ASAP7_75t_L g551 ( .A(n_552), .B(n_571), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_560), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_568), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_585), .Y(n_575) );
NOR3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .C(n_581), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AND4x1_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .C(n_592), .D(n_593), .Y(n_585) );
BUFx2_ASAP7_75t_L g679 ( .A(n_591), .Y(n_679) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_601), .B(n_610), .Y(n_600) );
NAND4xp25_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .C(n_606), .D(n_608), .Y(n_601) );
NAND4xp25_ASAP7_75t_SL g610 ( .A(n_611), .B(n_612), .C(n_615), .D(n_616), .Y(n_610) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx3_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND4xp75_ASAP7_75t_SL g624 ( .A(n_625), .B(n_628), .C(n_632), .D(n_637), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_647), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_644), .B(n_648), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g663 ( .A(n_646), .Y(n_663) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_659), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI222xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_664), .B1(n_665), .B2(n_690), .C1(n_693), .C2(n_697), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_664), .B(n_683), .Y(n_689) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_667), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_674), .C(n_683), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
NOR4xp25_ASAP7_75t_L g688 ( .A(n_669), .B(n_671), .C(n_675), .D(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
OAI221xp5_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_677), .B1(n_678), .B2(n_680), .C(n_681), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
CKINVDCx6p67_ASAP7_75t_R g691 ( .A(n_692), .Y(n_691) );
CKINVDCx16_ASAP7_75t_R g695 ( .A(n_694), .Y(n_695) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
endmodule