module real_jpeg_26229_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_148;
wire n_19;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_4),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_4),
.A2(n_42),
.B1(n_51),
.B2(n_52),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_4),
.A2(n_42),
.B1(n_67),
.B2(n_68),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_5),
.A2(n_51),
.B1(n_52),
.B2(n_66),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_6),
.B(n_36),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_6),
.B(n_52),
.C(n_54),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_6),
.A2(n_37),
.B1(n_40),
.B2(n_114),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_6),
.B(n_109),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_114),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_6),
.B(n_67),
.C(n_80),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_6),
.A2(n_69),
.B(n_222),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_85),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_7),
.A2(n_37),
.B1(n_40),
.B2(n_85),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_37),
.B1(n_40),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_9),
.A2(n_49),
.B1(n_67),
.B2(n_68),
.Y(n_172)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_11),
.A2(n_27),
.B1(n_37),
.B2(n_40),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_11),
.A2(n_27),
.B1(n_51),
.B2(n_52),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_11),
.A2(n_27),
.B1(n_67),
.B2(n_68),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_14),
.A2(n_37),
.B1(n_40),
.B2(n_58),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_14),
.A2(n_32),
.B1(n_45),
.B2(n_58),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_14),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_14),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_67),
.B1(n_68),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_15),
.A2(n_51),
.B1(n_52),
.B2(n_72),
.Y(n_130)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_16),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_148),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_146),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_125),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_20),
.B(n_125),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.C(n_99),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_21),
.A2(n_22),
.B1(n_86),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_62),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_46),
.B2(n_47),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_25),
.B(n_46),
.C(n_62),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_36),
.B2(n_41),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_26),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_28),
.B(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_30),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_30),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_30),
.A2(n_143),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_33),
.A2(n_37),
.B(n_113),
.C(n_115),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_SL g115 ( 
.A(n_34),
.B(n_40),
.C(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_35),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_35),
.B(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_37),
.B(n_187),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_41),
.Y(n_140)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B(n_56),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_48),
.A2(n_50),
.B1(n_60),
.B2(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_50),
.A2(n_56),
.B(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_52),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_52),
.B(n_230),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_57),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_59),
.A2(n_107),
.B1(n_109),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_60),
.A2(n_108),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_76),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_63),
.B(n_76),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_65),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_119)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_70),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_68),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_68),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_71),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_69),
.A2(n_75),
.B(n_88),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_69),
.A2(n_122),
.B1(n_124),
.B2(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_69),
.B(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_69),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_70),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_73),
.B(n_114),
.Y(n_247)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_75),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_77),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_77),
.A2(n_210),
.B(n_228),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_78),
.A2(n_95),
.B1(n_96),
.B2(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_78),
.B(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_78),
.A2(n_96),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_82),
.A2(n_83),
.B(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_82),
.A2(n_159),
.B(n_195),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_82),
.B(n_114),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_86),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_93),
.B1(n_97),
.B2(n_98),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_98),
.Y(n_134)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_92),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_96),
.B(n_160),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_99),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.C(n_110),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_100),
.B(n_105),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_110),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_119),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_111),
.A2(n_112),
.B1(n_119),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_113),
.A2(n_114),
.B(n_116),
.Y(n_162)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_120),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_124),
.A2(n_235),
.B(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_145),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_133),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_144),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B(n_142),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_179),
.B(n_266),
.C(n_271),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_173),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_163),
.C(n_166),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_151),
.A2(n_152),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_161),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_157),
.C(n_161),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_156),
.Y(n_168)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_166),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_174),
.B(n_177),
.C(n_178),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_259),
.B(n_265),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_211),
.B(n_258),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_200),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_184),
.B(n_200),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_193),
.C(n_197),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_185),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_188),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_193),
.A2(n_197),
.B1(n_198),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_201),
.B(n_207),
.C(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_252),
.B(n_257),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_231),
.B(n_251),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_225),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_225),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_219),
.C(n_220),
.Y(n_256)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_229),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_240),
.B(n_250),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_238),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_245),
.B(n_249),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_264),
.Y(n_265)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);


endmodule