module fake_jpeg_18792_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_60),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_52),
.B1(n_51),
.B2(n_63),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_72),
.B1(n_75),
.B2(n_54),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_69),
.A2(n_49),
.B1(n_50),
.B2(n_55),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_58),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_90),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_72),
.B1(n_42),
.B2(n_62),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_55),
.C(n_56),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_60),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_54),
.B(n_50),
.Y(n_94)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_104),
.B1(n_4),
.B2(n_5),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_25),
.Y(n_114)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_48),
.B1(n_45),
.B2(n_20),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_106),
.B1(n_6),
.B2(n_9),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_112),
.B1(n_116),
.B2(n_96),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_24),
.B(n_36),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_5),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.C(n_115),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_6),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_117),
.B(n_118),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_108),
.C(n_95),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_114),
.C(n_112),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_121),
.B1(n_100),
.B2(n_102),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_110),
.B(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_13),
.B(n_17),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_26),
.B(n_27),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_29),
.Y(n_130)
);


endmodule