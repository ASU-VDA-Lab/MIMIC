module fake_netlist_5_521_n_1939 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1939);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1939;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_368;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_31),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_115),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_168),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_38),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_72),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_25),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_25),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_80),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_69),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_30),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_96),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_58),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_57),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_165),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_51),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_93),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_92),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_61),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_90),
.Y(n_215)
);

BUFx8_ASAP7_75t_SL g216 ( 
.A(n_75),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_2),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_91),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_37),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_26),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_106),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_58),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_31),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_42),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_89),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_137),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_21),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_10),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_177),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_152),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_119),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_41),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_143),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_56),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_79),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_87),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_99),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_77),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_68),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_150),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_38),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_24),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_68),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_9),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_30),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_105),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_190),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_76),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_85),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_174),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_135),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_130),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_2),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_98),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_24),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_95),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_81),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_126),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_66),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_46),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_188),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_14),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_180),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_49),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_70),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_45),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_55),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_104),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_167),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_108),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_153),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_4),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_83),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_88),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_163),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_84),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_29),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_82),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_145),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_39),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_112),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_110),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_175),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_29),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_184),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_186),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_170),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_1),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_161),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_181),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_154),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_120),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_14),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_9),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_26),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_111),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_5),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_169),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_179),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_71),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_5),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_28),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_49),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_125),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_185),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_61),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_187),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_101),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_62),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_133),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_97),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_162),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_8),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_171),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_123),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_141),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_47),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_10),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_157),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_8),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_109),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_74),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_27),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_35),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_182),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_172),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_13),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_134),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_183),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_86),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_102),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_140),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_67),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_148),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_17),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_78),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_131),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_191),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_21),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_189),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_48),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_27),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_3),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_128),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_107),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_94),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_7),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_6),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_33),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_103),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_151),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_53),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_17),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_54),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_54),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_158),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_1),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_12),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_11),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_28),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_62),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_178),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_11),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_44),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_138),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_116),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_19),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_63),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_46),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_40),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_65),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_6),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_132),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_16),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_32),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_44),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_36),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_52),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_65),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_15),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_40),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_59),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_160),
.Y(n_386)
);

BUFx10_ASAP7_75t_L g387 ( 
.A(n_73),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_166),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_144),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_139),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_32),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_298),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_326),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_208),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_364),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_336),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_336),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_336),
.Y(n_401)
);

INVxp33_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_336),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_201),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_287),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_287),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_385),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_238),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_192),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_192),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_192),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_363),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_192),
.Y(n_416)
);

INVxp33_ASAP7_75t_SL g417 ( 
.A(n_203),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_192),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_256),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_239),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_249),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_256),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_256),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_256),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_256),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_246),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_230),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_229),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_382),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_250),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_237),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_246),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_310),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_323),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_323),
.Y(n_435)
);

INVxp33_ASAP7_75t_SL g436 ( 
.A(n_203),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_242),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_367),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_254),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_367),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_367),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_244),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_273),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_197),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_225),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_226),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_245),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_247),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_248),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_265),
.Y(n_452)
);

BUFx6f_ASAP7_75t_SL g453 ( 
.A(n_234),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_275),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_290),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_280),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_276),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_233),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_262),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_291),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_301),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_300),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_331),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_305),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_306),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_233),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_327),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_216),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_207),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_263),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_330),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_344),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_388),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_346),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_356),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_358),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_378),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_381),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_272),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_195),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_267),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_269),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_232),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_272),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_198),
.Y(n_486)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_207),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_270),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_236),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_307),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_240),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_241),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_307),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_198),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_296),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_251),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_227),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_297),
.Y(n_498)
);

INVxp33_ASAP7_75t_SL g499 ( 
.A(n_214),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_328),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_396),
.A2(n_309),
.B1(n_312),
.B2(n_304),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_469),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_380),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_438),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_429),
.A2(n_321),
.B1(n_338),
.B2(n_316),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_484),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_397),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_412),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_424),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_412),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_489),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_413),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_392),
.A2(n_243),
.B(n_200),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_424),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_408),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_328),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_491),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_415),
.B(n_341),
.Y(n_522)
);

NOR2x1_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_341),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_414),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_416),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_444),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_416),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_496),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_405),
.Y(n_529)
);

AND2x2_ASAP7_75t_R g530 ( 
.A(n_394),
.B(n_210),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_418),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_485),
.B(n_380),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_L g533 ( 
.A(n_393),
.B(n_214),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_440),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_419),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_408),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_473),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_458),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_393),
.B(n_234),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_419),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_415),
.B(n_194),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_411),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_455),
.B(n_194),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_422),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_423),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_423),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_425),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_425),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_441),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_442),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_427),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_395),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_399),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_439),
.B(n_200),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_406),
.B(n_243),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_417),
.A2(n_222),
.B1(n_362),
.B2(n_220),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_407),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_409),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_395),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_420),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_428),
.B(n_349),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_410),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_R g565 ( 
.A(n_468),
.B(n_427),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_400),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_401),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_426),
.B(n_227),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_431),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_398),
.B(n_403),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_404),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_398),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_421),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_433),
.B(n_221),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_458),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_466),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_466),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_432),
.B(n_255),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_430),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_434),
.B(n_255),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_445),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_435),
.B(n_258),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_446),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_486),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_556),
.B(n_417),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_570),
.B(n_431),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_570),
.B(n_437),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_538),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_520),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_538),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_545),
.A2(n_258),
.B1(n_377),
.B2(n_320),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_504),
.B(n_494),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_554),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_R g595 ( 
.A(n_507),
.B(n_457),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_563),
.B(n_481),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_554),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_520),
.Y(n_598)
);

NOR2x1p5_ASAP7_75t_L g599 ( 
.A(n_507),
.B(n_437),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_575),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_575),
.Y(n_601)
);

AOI21x1_ASAP7_75t_L g602 ( 
.A1(n_572),
.A2(n_311),
.B(n_299),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_570),
.B(n_443),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_518),
.Y(n_604)
);

OAI22xp33_ASAP7_75t_L g605 ( 
.A1(n_501),
.A2(n_402),
.B1(n_235),
.B2(n_361),
.Y(n_605)
);

AO22x2_ASAP7_75t_L g606 ( 
.A1(n_503),
.A2(n_377),
.B1(n_320),
.B2(n_311),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_531),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_504),
.B(n_494),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_518),
.B(n_443),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_572),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_531),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_558),
.B(n_461),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_512),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_534),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_518),
.A2(n_469),
.B1(n_487),
.B2(n_436),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_L g616 ( 
.A1(n_506),
.A2(n_569),
.B1(n_574),
.B2(n_500),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_534),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_552),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_552),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_510),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_557),
.A2(n_487),
.B1(n_499),
.B2(n_436),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_536),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_536),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_512),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_561),
.Y(n_625)
);

AND3x2_ASAP7_75t_L g626 ( 
.A(n_508),
.B(n_315),
.C(n_299),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_561),
.B(n_449),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_561),
.B(n_449),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_521),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_555),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_536),
.Y(n_631)
);

CKINVDCx6p67_ASAP7_75t_R g632 ( 
.A(n_529),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_508),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_523),
.B(n_450),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_569),
.B(n_450),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_575),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_566),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_576),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_517),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_522),
.Y(n_640)
);

INVxp33_ASAP7_75t_SL g641 ( 
.A(n_502),
.Y(n_641)
);

AOI21x1_ASAP7_75t_L g642 ( 
.A1(n_555),
.A2(n_386),
.B(n_315),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_576),
.Y(n_643)
);

INVx8_ASAP7_75t_L g644 ( 
.A(n_543),
.Y(n_644)
);

BUFx6f_ASAP7_75t_SL g645 ( 
.A(n_543),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_576),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_566),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_540),
.B(n_499),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_557),
.A2(n_386),
.B1(n_448),
.B2(n_447),
.Y(n_649)
);

AND2x2_ASAP7_75t_SL g650 ( 
.A(n_553),
.B(n_205),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_567),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_577),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_566),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_567),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_577),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_539),
.B(n_459),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_532),
.B(n_497),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_553),
.B(n_459),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_517),
.B(n_470),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_566),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_532),
.B(n_470),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_577),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_537),
.B(n_482),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_539),
.B(n_482),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_533),
.B(n_488),
.C(n_483),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_584),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_510),
.Y(n_667)
);

INVxp33_ASAP7_75t_SL g668 ( 
.A(n_565),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_522),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_544),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_R g672 ( 
.A(n_521),
.B(n_463),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_510),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_510),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_559),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_537),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_510),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_566),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_528),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_560),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_564),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_516),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_528),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_543),
.B(n_205),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_522),
.B(n_483),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_509),
.Y(n_686)
);

AOI21x1_ASAP7_75t_L g687 ( 
.A1(n_578),
.A2(n_581),
.B(n_511),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_568),
.B(n_488),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_571),
.B(n_495),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_509),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_511),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_568),
.B(n_451),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_516),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_513),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_557),
.B(n_495),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_516),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_516),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_513),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_562),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_514),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_516),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_526),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_571),
.B(n_498),
.Y(n_703)
);

INVxp33_ASAP7_75t_SL g704 ( 
.A(n_573),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_514),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_519),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_571),
.B(n_498),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_571),
.B(n_252),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_519),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_526),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_571),
.B(n_253),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_583),
.B(n_234),
.Y(n_712)
);

AO21x2_ASAP7_75t_L g713 ( 
.A1(n_515),
.A2(n_204),
.B(n_196),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_583),
.A2(n_515),
.B1(n_585),
.B2(n_454),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_585),
.B(n_387),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_505),
.B(n_452),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_524),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_526),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_541),
.Y(n_719)
);

INVx4_ASAP7_75t_SL g720 ( 
.A(n_526),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_535),
.A2(n_453),
.B1(n_193),
.B2(n_199),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_573),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_585),
.A2(n_467),
.B1(n_479),
.B2(n_478),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_524),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_525),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_526),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_541),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_525),
.Y(n_728)
);

INVxp33_ASAP7_75t_SL g729 ( 
.A(n_582),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_527),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_527),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_542),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_579),
.B(n_456),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_542),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_579),
.B(n_453),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_547),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_547),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_640),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_604),
.B(n_548),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_640),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_650),
.B(n_604),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_650),
.B(n_205),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_600),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_670),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_669),
.B(n_548),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_600),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_616),
.B(n_205),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_586),
.B(n_582),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_688),
.B(n_609),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_587),
.A2(n_271),
.B1(n_293),
.B2(n_288),
.Y(n_750)
);

INVxp33_ASAP7_75t_L g751 ( 
.A(n_595),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_669),
.B(n_549),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_594),
.B(n_597),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_670),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_688),
.B(n_460),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_594),
.B(n_549),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_656),
.B(n_193),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_601),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_675),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_597),
.B(n_541),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_610),
.B(n_541),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_633),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_610),
.B(n_541),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_664),
.B(n_627),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_593),
.B(n_546),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_628),
.B(n_588),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_593),
.B(n_546),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_608),
.B(n_546),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_603),
.A2(n_462),
.B(n_464),
.C(n_465),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_648),
.A2(n_302),
.B1(n_257),
.B2(n_259),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_608),
.B(n_546),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_675),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_635),
.B(n_199),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_686),
.B(n_546),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_689),
.B(n_205),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_655),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_655),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_722),
.B(n_530),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_703),
.B(n_707),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_690),
.B(n_550),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_644),
.Y(n_781)
);

INVx8_ASAP7_75t_L g782 ( 
.A(n_644),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_661),
.A2(n_308),
.B1(n_289),
.B2(n_292),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_635),
.B(n_202),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_680),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_690),
.B(n_550),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_596),
.B(n_202),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_691),
.B(n_694),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_691),
.B(n_550),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_633),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_615),
.B(n_195),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_681),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_694),
.B(n_550),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_698),
.B(n_585),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_698),
.B(n_585),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_692),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_685),
.B(n_206),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_636),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_625),
.B(n_348),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_657),
.B(n_195),
.Y(n_800)
);

OR2x6_ASAP7_75t_SL g801 ( 
.A(n_589),
.B(n_591),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_708),
.A2(n_551),
.B(n_219),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_700),
.B(n_551),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_733),
.Y(n_804)
);

INVx6_ASAP7_75t_L g805 ( 
.A(n_644),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_644),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_692),
.Y(n_807)
);

AOI22x1_ASAP7_75t_SL g808 ( 
.A1(n_613),
.A2(n_580),
.B1(n_217),
.B2(n_384),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_695),
.B(n_666),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_733),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_705),
.B(n_706),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_665),
.B(n_206),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_692),
.B(n_712),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_706),
.B(n_551),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_634),
.A2(n_645),
.B1(n_692),
.B2(n_658),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_605),
.B(n_209),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_625),
.B(n_348),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_709),
.B(n_212),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_716),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_638),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_714),
.B(n_348),
.Y(n_821)
);

BUFx8_ASAP7_75t_L g822 ( 
.A(n_722),
.Y(n_822)
);

AND2x4_ASAP7_75t_SL g823 ( 
.A(n_632),
.B(n_387),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_622),
.B(n_348),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_709),
.B(n_717),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_717),
.B(n_209),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_724),
.B(n_224),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_622),
.B(n_348),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_724),
.B(n_211),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_623),
.B(n_368),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_623),
.B(n_368),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_725),
.B(n_211),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_657),
.B(n_471),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_728),
.B(n_228),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_716),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_L g836 ( 
.A(n_684),
.B(n_233),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_737),
.B(n_213),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_730),
.B(n_260),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_606),
.A2(n_368),
.B1(n_233),
.B2(n_261),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_621),
.A2(n_278),
.B1(n_274),
.B2(n_266),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_730),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_731),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_731),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_631),
.B(n_368),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_735),
.B(n_472),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_631),
.B(n_233),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_659),
.B(n_663),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_732),
.B(n_264),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_L g849 ( 
.A(n_639),
.B(n_676),
.C(n_591),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_732),
.B(n_734),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_734),
.B(n_286),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_643),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_620),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_687),
.B(n_213),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_620),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_736),
.B(n_313),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_620),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_630),
.B(n_233),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_736),
.B(n_314),
.Y(n_859)
);

AOI22x1_ASAP7_75t_L g860 ( 
.A1(n_606),
.A2(n_369),
.B1(n_325),
.B2(n_333),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_646),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_626),
.B(n_474),
.Y(n_862)
);

BUFx12f_ASAP7_75t_SL g863 ( 
.A(n_668),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_630),
.B(n_334),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_599),
.B(n_721),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_592),
.A2(n_475),
.B(n_477),
.C(n_476),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_606),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_651),
.B(n_335),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_L g869 ( 
.A(n_649),
.B(n_215),
.C(n_347),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_672),
.B(n_231),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_646),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_651),
.B(n_654),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_613),
.B(n_624),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_645),
.A2(n_711),
.B1(n_606),
.B2(n_715),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_654),
.B(n_339),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_719),
.B(n_353),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_618),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_624),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_719),
.B(n_354),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_687),
.B(n_233),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_629),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_652),
.B(n_376),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_662),
.B(n_389),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_619),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_645),
.A2(n_215),
.B1(n_218),
.B2(n_390),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_662),
.B(n_268),
.Y(n_886)
);

INVx5_ASAP7_75t_L g887 ( 
.A(n_781),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_764),
.B(n_607),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_764),
.B(n_607),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_766),
.B(n_611),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_766),
.B(n_611),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_779),
.B(n_614),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_841),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_833),
.B(n_671),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_749),
.A2(n_619),
.B(n_667),
.C(n_726),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_842),
.Y(n_896)
);

NAND2x1p5_ASAP7_75t_L g897 ( 
.A(n_781),
.B(n_637),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_843),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_754),
.Y(n_899)
);

NAND3xp33_ASAP7_75t_SL g900 ( 
.A(n_816),
.B(n_679),
.C(n_629),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_877),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_863),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_777),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_884),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_754),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_753),
.B(n_617),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_754),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_788),
.B(n_617),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_754),
.B(n_641),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_833),
.B(n_699),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_850),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_811),
.B(n_713),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_800),
.B(n_679),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_825),
.B(n_765),
.Y(n_914)
);

NAND3xp33_ASAP7_75t_SL g915 ( 
.A(n_816),
.B(n_683),
.C(n_589),
.Y(n_915)
);

NOR2x2_ASAP7_75t_L g916 ( 
.A(n_778),
.B(n_612),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_767),
.B(n_713),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_755),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_747),
.A2(n_713),
.B1(n_684),
.B2(n_598),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_777),
.Y(n_920)
);

BUFx8_ASAP7_75t_L g921 ( 
.A(n_878),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_768),
.B(n_590),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_872),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_822),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_757),
.B(n_641),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_748),
.B(n_704),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_SL g927 ( 
.A1(n_791),
.A2(n_729),
.B1(n_704),
.B2(n_453),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_771),
.B(n_741),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_819),
.B(n_683),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_798),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_790),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_759),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_762),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_835),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_757),
.A2(n_729),
.B1(n_684),
.B2(n_660),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_738),
.Y(n_936)
);

INVxp33_ASAP7_75t_L g937 ( 
.A(n_873),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_740),
.B(n_667),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_772),
.B(n_674),
.Y(n_939)
);

INVx5_ASAP7_75t_L g940 ( 
.A(n_781),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_847),
.B(n_612),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_820),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_781),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_847),
.A2(n_684),
.B1(n_660),
.B2(n_637),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_785),
.B(n_674),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_796),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_821),
.A2(n_660),
.B(n_637),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_744),
.B(n_682),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_SL g949 ( 
.A(n_865),
.B(n_218),
.Y(n_949)
);

INVx5_ASAP7_75t_L g950 ( 
.A(n_806),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_809),
.A2(n_684),
.B1(n_726),
.B2(n_718),
.Y(n_951)
);

NAND3xp33_ASAP7_75t_L g952 ( 
.A(n_773),
.B(n_723),
.C(n_284),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_792),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_738),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_804),
.B(n_682),
.Y(n_955)
);

BUFx4f_ASAP7_75t_L g956 ( 
.A(n_881),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_862),
.Y(n_957)
);

BUFx8_ASAP7_75t_L g958 ( 
.A(n_870),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_743),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_823),
.Y(n_960)
);

CKINVDCx6p67_ASAP7_75t_R g961 ( 
.A(n_801),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_806),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_809),
.B(n_223),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_747),
.A2(n_684),
.B1(n_718),
.B2(n_710),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_822),
.Y(n_965)
);

BUFx8_ASAP7_75t_L g966 ( 
.A(n_862),
.Y(n_966)
);

BUFx12f_ASAP7_75t_SL g967 ( 
.A(n_778),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_746),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_806),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_806),
.B(n_223),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_796),
.B(n_696),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_758),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_853),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_845),
.B(n_284),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_807),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_L g976 ( 
.A(n_773),
.B(n_784),
.C(n_787),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_810),
.B(n_696),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_782),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_784),
.B(n_632),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_807),
.B(n_697),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_813),
.A2(n_684),
.B1(n_710),
.B2(n_702),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_853),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_756),
.B(n_697),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_776),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_812),
.B(n_347),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_823),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_739),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_867),
.B(n_701),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_852),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_745),
.B(n_701),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_752),
.B(n_854),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_812),
.B(n_359),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_742),
.A2(n_702),
.B1(n_233),
.B2(n_677),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_861),
.Y(n_994)
);

BUFx4f_ASAP7_75t_L g995 ( 
.A(n_782),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_871),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_815),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_854),
.B(n_673),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_813),
.Y(n_999)
);

OR2x4_ASAP7_75t_L g1000 ( 
.A(n_787),
.B(n_497),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_751),
.B(n_359),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_855),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_874),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_760),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_797),
.B(n_365),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_849),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_855),
.Y(n_1007)
);

AO22x1_ASAP7_75t_L g1008 ( 
.A1(n_797),
.A2(n_384),
.B1(n_283),
.B2(n_217),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_855),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_826),
.B(n_365),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_770),
.B(n_390),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_839),
.B(n_677),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_839),
.B(n_693),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_826),
.B(n_352),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_742),
.B(n_818),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_827),
.B(n_693),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_761),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_840),
.A2(n_693),
.B1(n_387),
.B2(n_727),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_763),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_774),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_780),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_786),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_789),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_793),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_803),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_794),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_886),
.Y(n_1027)
);

AND2x6_ASAP7_75t_SL g1028 ( 
.A(n_808),
.B(n_352),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_750),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_834),
.B(n_620),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_829),
.B(n_727),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_885),
.B(n_283),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_821),
.A2(n_345),
.B1(n_350),
.B2(n_351),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_860),
.A2(n_727),
.B1(n_343),
.B2(n_340),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_832),
.A2(n_277),
.B1(n_279),
.B2(n_281),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_876),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_869),
.B(n_720),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_795),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_837),
.B(n_282),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_837),
.A2(n_332),
.B(n_329),
.C(n_324),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_814),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_783),
.B(n_857),
.Y(n_1042)
);

AOI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_838),
.A2(n_303),
.B(n_295),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_846),
.B(n_720),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_879),
.A2(n_285),
.B1(n_294),
.B2(n_317),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_883),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_SL g1047 ( 
.A(n_769),
.B(n_379),
.C(n_345),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_864),
.B(n_350),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_868),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_976),
.A2(n_859),
.B(n_848),
.C(n_851),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_931),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_902),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_887),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_966),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_946),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1049),
.B(n_857),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_1005),
.A2(n_858),
.B1(n_880),
.B2(n_846),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_918),
.B(n_866),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_988),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_1011),
.A2(n_775),
.B(n_880),
.C(n_856),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_926),
.B(n_875),
.Y(n_1061)
);

AOI22x1_ASAP7_75t_L g1062 ( 
.A1(n_1046),
.A2(n_802),
.B1(n_775),
.B2(n_318),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_973),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_975),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_941),
.A2(n_805),
.B1(n_858),
.B2(n_882),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_991),
.A2(n_923),
.B1(n_914),
.B2(n_891),
.Y(n_1066)
);

AOI21xp33_ASAP7_75t_L g1067 ( 
.A1(n_985),
.A2(n_371),
.B(n_370),
.Y(n_1067)
);

NAND3xp33_ASAP7_75t_L g1068 ( 
.A(n_1032),
.B(n_373),
.C(n_379),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_890),
.A2(n_799),
.B(n_817),
.C(n_831),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_987),
.B(n_805),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_988),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_991),
.A2(n_678),
.B(n_647),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_943),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_911),
.B(n_805),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_999),
.B(n_799),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_930),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_998),
.A2(n_653),
.B(n_678),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_942),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_890),
.B(n_817),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_933),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_943),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_966),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_932),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_997),
.A2(n_319),
.B1(n_337),
.B2(n_322),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_891),
.A2(n_844),
.B1(n_824),
.B2(n_828),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_SL g1086 ( 
.A(n_900),
.B(n_915),
.C(n_949),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_894),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_943),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_888),
.B(n_830),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_953),
.Y(n_1090)
);

AO32x1_ASAP7_75t_L g1091 ( 
.A1(n_1014),
.A2(n_602),
.A3(n_642),
.B1(n_830),
.B2(n_836),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_889),
.A2(n_374),
.B1(n_355),
.B2(n_357),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_998),
.A2(n_678),
.B(n_653),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_929),
.B(n_352),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_889),
.A2(n_374),
.B1(n_355),
.B2(n_357),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_937),
.B(n_351),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_922),
.A2(n_678),
.B(n_653),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_924),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_925),
.B(n_647),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_934),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_978),
.B(n_720),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_922),
.A2(n_678),
.B(n_653),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1036),
.B(n_360),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_894),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1015),
.A2(n_375),
.B1(n_366),
.B2(n_370),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_928),
.A2(n_602),
.B(n_642),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_962),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_910),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_979),
.B(n_1048),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1003),
.A2(n_373),
.B1(n_366),
.B2(n_383),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_910),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1000),
.B(n_360),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1001),
.B(n_371),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1027),
.B(n_372),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_928),
.B(n_372),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1004),
.B(n_1020),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1015),
.A2(n_383),
.B1(n_375),
.B2(n_647),
.Y(n_1117)
);

INVxp67_ASAP7_75t_SL g1118 ( 
.A(n_973),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1000),
.B(n_0),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_994),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_956),
.B(n_0),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_912),
.A2(n_156),
.B(n_149),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_SL g1123 ( 
.A(n_1033),
.B(n_3),
.C(n_4),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_965),
.Y(n_1124)
);

NOR3xp33_ASAP7_75t_L g1125 ( 
.A(n_927),
.B(n_7),
.C(n_12),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_901),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1030),
.A2(n_147),
.B(n_146),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_963),
.B(n_15),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1029),
.B(n_16),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_SL g1130 ( 
.A1(n_1042),
.A2(n_142),
.B(n_136),
.C(n_129),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1023),
.B(n_1024),
.Y(n_1131)
);

OAI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_992),
.A2(n_18),
.B(n_19),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_895),
.A2(n_18),
.B(n_20),
.C(n_22),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_990),
.A2(n_127),
.B(n_122),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_939),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_978),
.B(n_100),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_962),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_939),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_962),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_971),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_921),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1006),
.B(n_1010),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_990),
.A2(n_121),
.B(n_118),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_955),
.A2(n_977),
.B(n_906),
.C(n_908),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_952),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_945),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_958),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_921),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1026),
.B(n_23),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_957),
.B(n_33),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_971),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_945),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1038),
.B(n_34),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_958),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_904),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_912),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_980),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_969),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_967),
.Y(n_1159)
);

INVx4_ASAP7_75t_L g1160 ( 
.A(n_887),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_980),
.B(n_113),
.Y(n_1161)
);

OAI22x1_ASAP7_75t_L g1162 ( 
.A1(n_909),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_887),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_955),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_969),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_940),
.B(n_43),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_977),
.B(n_43),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_893),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_896),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_906),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_898),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_947),
.A2(n_67),
.B(n_51),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_L g1173 ( 
.A(n_986),
.B(n_50),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_938),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_908),
.A2(n_50),
.B(n_52),
.C(n_53),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_947),
.A2(n_55),
.B(n_56),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_969),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1025),
.B(n_60),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1039),
.B(n_60),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1040),
.A2(n_63),
.B(n_64),
.C(n_66),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_SL g1181 ( 
.A(n_940),
.B(n_64),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_940),
.A2(n_950),
.B(n_917),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_950),
.A2(n_917),
.B(n_1016),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_899),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1073),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_1077),
.Y(n_1186)
);

AO21x2_ASAP7_75t_L g1187 ( 
.A1(n_1183),
.A2(n_1031),
.B(n_944),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1164),
.B(n_1041),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_SL g1189 ( 
.A(n_1113),
.B(n_960),
.C(n_1047),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1060),
.A2(n_950),
.B(n_897),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1144),
.A2(n_950),
.B(n_1016),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1109),
.B(n_899),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1051),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1085),
.A2(n_1012),
.A3(n_1013),
.B(n_892),
.Y(n_1194)
);

OR2x6_ASAP7_75t_L g1195 ( 
.A(n_1136),
.B(n_899),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1059),
.B(n_1022),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1071),
.B(n_1019),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1144),
.A2(n_983),
.B(n_1013),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1116),
.A2(n_919),
.B1(n_935),
.B2(n_936),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1135),
.B(n_1017),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1097),
.A2(n_1102),
.B(n_1072),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1179),
.A2(n_1043),
.B(n_1035),
.C(n_1034),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1080),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1050),
.A2(n_995),
.B(n_1021),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1050),
.A2(n_1089),
.B(n_1079),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1138),
.B(n_936),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1128),
.A2(n_1043),
.B(n_974),
.C(n_970),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1057),
.A2(n_995),
.B(n_982),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_SL g1209 ( 
.A(n_1125),
.B(n_1033),
.C(n_1018),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1142),
.B(n_1008),
.Y(n_1210)
);

AOI21xp33_ASAP7_75t_L g1211 ( 
.A1(n_1180),
.A2(n_989),
.B(n_996),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1083),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1080),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1069),
.A2(n_951),
.B(n_981),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1061),
.B(n_903),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1167),
.A2(n_954),
.A3(n_920),
.B(n_984),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1068),
.B(n_1045),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1131),
.A2(n_1007),
.B(n_982),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1146),
.B(n_907),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1152),
.A2(n_1007),
.B(n_982),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1074),
.A2(n_905),
.B(n_907),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1055),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1122),
.A2(n_993),
.B(n_964),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1114),
.B(n_1094),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1172),
.A2(n_968),
.B(n_959),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1115),
.B(n_972),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1053),
.B(n_905),
.Y(n_1227)
);

AOI221x1_ASAP7_75t_L g1228 ( 
.A1(n_1125),
.A2(n_1176),
.B1(n_1132),
.B2(n_1156),
.C(n_1162),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1096),
.B(n_938),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1070),
.A2(n_905),
.B(n_1044),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1053),
.A2(n_1044),
.B(n_1009),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_1073),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_L g1233 ( 
.A(n_1052),
.B(n_948),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1160),
.A2(n_1002),
.B(n_1037),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1055),
.Y(n_1235)
);

NAND3x1_ASAP7_75t_L g1236 ( 
.A(n_1121),
.B(n_916),
.C(n_1028),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1062),
.A2(n_948),
.B(n_961),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1167),
.B(n_1075),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1075),
.B(n_1129),
.Y(n_1239)
);

O2A1O1Ixp5_ASAP7_75t_L g1240 ( 
.A1(n_1056),
.A2(n_1099),
.B(n_1153),
.C(n_1149),
.Y(n_1240)
);

NOR2x1_ASAP7_75t_L g1241 ( 
.A(n_1160),
.B(n_1163),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1090),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1168),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1129),
.B(n_1169),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1103),
.B(n_1104),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1100),
.B(n_1067),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1073),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1100),
.B(n_1064),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1154),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1171),
.B(n_1058),
.Y(n_1250)
);

AO21x1_ASAP7_75t_L g1251 ( 
.A1(n_1133),
.A2(n_1180),
.B(n_1170),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1110),
.A2(n_1126),
.B1(n_1155),
.B2(n_1123),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1134),
.A2(n_1143),
.B(n_1127),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1073),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1163),
.A2(n_1091),
.B(n_1065),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1110),
.A2(n_1123),
.B1(n_1161),
.B2(n_1151),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1119),
.A2(n_1112),
.B(n_1175),
.Y(n_1257)
);

AOI221xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1145),
.A2(n_1133),
.B1(n_1175),
.B2(n_1170),
.C(n_1117),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_SL g1259 ( 
.A(n_1086),
.B(n_1084),
.C(n_1112),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1178),
.A2(n_1086),
.B(n_1130),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1064),
.B(n_1108),
.Y(n_1261)
);

OAI21xp33_ASAP7_75t_L g1262 ( 
.A1(n_1105),
.A2(n_1092),
.B(n_1095),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1140),
.B(n_1151),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1140),
.B(n_1157),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1091),
.A2(n_1063),
.B(n_1118),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1076),
.A2(n_1120),
.B(n_1078),
.Y(n_1266)
);

AOI221x1_ASAP7_75t_L g1267 ( 
.A1(n_1161),
.A2(n_1150),
.B1(n_1174),
.B2(n_1136),
.C(n_1165),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1157),
.B(n_1111),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_R g1269 ( 
.A(n_1159),
.B(n_1098),
.Y(n_1269)
);

AO21x1_ASAP7_75t_L g1270 ( 
.A1(n_1166),
.A2(n_1118),
.B(n_1063),
.Y(n_1270)
);

NAND2x1_ASAP7_75t_L g1271 ( 
.A(n_1088),
.B(n_1158),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1184),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1091),
.A2(n_1173),
.B(n_1181),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1081),
.B(n_1137),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1177),
.Y(n_1275)
);

AOI21xp33_ASAP7_75t_L g1276 ( 
.A1(n_1087),
.A2(n_1137),
.B(n_1081),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1141),
.A2(n_1148),
.B1(n_1124),
.B2(n_1147),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1081),
.A2(n_1107),
.B(n_1137),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1081),
.B(n_1107),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1107),
.B(n_1137),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1107),
.A2(n_1139),
.B(n_1177),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1139),
.B(n_1177),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1177),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1139),
.A2(n_1101),
.B(n_1054),
.C(n_1082),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1101),
.A2(n_914),
.B(n_991),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1115),
.B(n_918),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1183),
.A2(n_1106),
.B(n_998),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1066),
.B(n_1164),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1115),
.B(n_918),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1066),
.A2(n_914),
.B(n_991),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_1077),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1066),
.B(n_1164),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1066),
.A2(n_914),
.B(n_991),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1066),
.A2(n_914),
.B(n_991),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1113),
.A2(n_1005),
.B1(n_976),
.B2(n_926),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1066),
.A2(n_914),
.B(n_991),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1066),
.B(n_1164),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1183),
.A2(n_1060),
.A3(n_895),
.B(n_1066),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_1077),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1066),
.B(n_1164),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_1077),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1066),
.B(n_1164),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1083),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1115),
.B(n_918),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1051),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1060),
.A2(n_991),
.B(n_914),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1066),
.A2(n_914),
.B(n_991),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1051),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1115),
.B(n_918),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1066),
.B(n_1164),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_1077),
.Y(n_1311)
);

O2A1O1Ixp5_ASAP7_75t_L g1312 ( 
.A1(n_1113),
.A2(n_1005),
.B(n_976),
.C(n_747),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1083),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1115),
.B(n_918),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1179),
.A2(n_976),
.B(n_1005),
.C(n_1113),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1183),
.A2(n_1060),
.A3(n_895),
.B(n_1066),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1109),
.B(n_913),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_1077),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1083),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1066),
.A2(n_914),
.B(n_991),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1066),
.B(n_1164),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1066),
.A2(n_914),
.B(n_991),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1051),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1183),
.A2(n_1106),
.B(n_998),
.Y(n_1324)
);

INVxp67_ASAP7_75t_SL g1325 ( 
.A(n_1080),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_SL g1326 ( 
.A1(n_1156),
.A2(n_747),
.B(n_976),
.C(n_742),
.Y(n_1326)
);

OR2x6_ASAP7_75t_L g1327 ( 
.A(n_1136),
.B(n_1161),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1060),
.A2(n_991),
.B(n_914),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1183),
.A2(n_1106),
.B(n_998),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1212),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1301),
.A2(n_1318),
.B(n_1311),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1224),
.B(n_1229),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1193),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1239),
.B(n_1238),
.Y(n_1335)
);

AO21x2_ASAP7_75t_L g1336 ( 
.A1(n_1255),
.A2(n_1191),
.B(n_1306),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1264),
.B(n_1268),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1244),
.B(n_1245),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1249),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1295),
.A2(n_1259),
.B1(n_1210),
.B2(n_1217),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1315),
.A2(n_1312),
.B(n_1257),
.C(n_1238),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1327),
.B(n_1233),
.Y(n_1342)
);

OAI222xp33_ASAP7_75t_L g1343 ( 
.A1(n_1239),
.A2(n_1256),
.B1(n_1252),
.B2(n_1244),
.C1(n_1250),
.C2(n_1297),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1305),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1317),
.A2(n_1189),
.B1(n_1262),
.B2(n_1257),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1209),
.A2(n_1251),
.B1(n_1256),
.B2(n_1252),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1203),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1325),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1250),
.A2(n_1228),
.B1(n_1267),
.B2(n_1289),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_SL g1350 ( 
.A1(n_1202),
.A2(n_1207),
.B(n_1297),
.C(n_1321),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1306),
.A2(n_1328),
.B(n_1214),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1328),
.A2(n_1205),
.B(n_1265),
.Y(n_1352)
);

NAND2x1p5_ASAP7_75t_L g1353 ( 
.A(n_1241),
.B(n_1192),
.Y(n_1353)
);

A2O1A1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1290),
.A2(n_1293),
.B(n_1296),
.C(n_1294),
.Y(n_1354)
);

INVx5_ASAP7_75t_L g1355 ( 
.A(n_1185),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1214),
.A2(n_1198),
.B(n_1322),
.Y(n_1356)
);

AOI21xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1286),
.A2(n_1304),
.B(n_1309),
.Y(n_1357)
);

NAND2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1278),
.B(n_1281),
.Y(n_1358)
);

AOI222xp33_ASAP7_75t_L g1359 ( 
.A1(n_1246),
.A2(n_1226),
.B1(n_1313),
.B2(n_1303),
.C1(n_1243),
.C2(n_1319),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1232),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1307),
.A2(n_1320),
.B(n_1285),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1242),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1258),
.A2(n_1273),
.B(n_1211),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1208),
.A2(n_1204),
.B(n_1220),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1314),
.B(n_1226),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1213),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1260),
.A2(n_1302),
.B1(n_1310),
.B2(n_1300),
.Y(n_1367)
);

AOI221xp5_ASAP7_75t_L g1368 ( 
.A1(n_1258),
.A2(n_1326),
.B1(n_1260),
.B2(n_1292),
.C(n_1288),
.Y(n_1368)
);

AOI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1288),
.A2(n_1300),
.B(n_1302),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1292),
.A2(n_1310),
.B(n_1321),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1196),
.B(n_1197),
.Y(n_1371)
);

INVxp67_ASAP7_75t_SL g1372 ( 
.A(n_1219),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1215),
.A2(n_1211),
.B1(n_1200),
.B2(n_1188),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1195),
.B(n_1270),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1188),
.A2(n_1200),
.B1(n_1196),
.B2(n_1197),
.Y(n_1375)
);

AO21x1_ASAP7_75t_L g1376 ( 
.A1(n_1199),
.A2(n_1218),
.B(n_1219),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1206),
.A2(n_1195),
.B1(n_1261),
.B2(n_1222),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1266),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1206),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1263),
.A2(n_1235),
.B1(n_1199),
.B2(n_1223),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1287),
.A2(n_1187),
.B(n_1234),
.Y(n_1381)
);

AO32x2_ASAP7_75t_L g1382 ( 
.A1(n_1194),
.A2(n_1232),
.A3(n_1216),
.B1(n_1298),
.B2(n_1316),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_L g1383 ( 
.A(n_1240),
.B(n_1323),
.C(n_1308),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1237),
.A2(n_1225),
.B(n_1324),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1230),
.A2(n_1221),
.B(n_1231),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1223),
.A2(n_1253),
.B1(n_1272),
.B2(n_1287),
.Y(n_1386)
);

CKINVDCx14_ASAP7_75t_R g1387 ( 
.A(n_1277),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1253),
.A2(n_1329),
.B(n_1324),
.Y(n_1388)
);

AOI221xp5_ASAP7_75t_SL g1389 ( 
.A1(n_1276),
.A2(n_1275),
.B1(n_1283),
.B2(n_1280),
.C(n_1282),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1236),
.A2(n_1227),
.B1(n_1275),
.B2(n_1280),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1274),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1227),
.A2(n_1282),
.B(n_1274),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1187),
.A2(n_1279),
.B1(n_1185),
.B2(n_1254),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1216),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1185),
.B(n_1247),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1216),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1247),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1271),
.A2(n_1298),
.B(n_1316),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1247),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1284),
.A2(n_1194),
.B(n_1254),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1239),
.B(n_1238),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1239),
.B(n_1238),
.Y(n_1403)
);

AO31x2_ASAP7_75t_L g1404 ( 
.A1(n_1251),
.A2(n_1255),
.A3(n_1265),
.B(n_1191),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1255),
.A2(n_1191),
.B(n_1306),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1212),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1327),
.B(n_1233),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1239),
.B(n_1238),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1201),
.A2(n_1291),
.B(n_1186),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1306),
.A2(n_1328),
.B(n_1293),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1255),
.A2(n_1191),
.B(n_1306),
.Y(n_1413)
);

XNOR2xp5_ASAP7_75t_L g1414 ( 
.A(n_1236),
.B(n_671),
.Y(n_1414)
);

A2O1A1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1315),
.A2(n_1295),
.B(n_1312),
.C(n_976),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1193),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1249),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1248),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1209),
.A2(n_1125),
.B1(n_976),
.B2(n_1262),
.Y(n_1419)
);

INVx8_ASAP7_75t_L g1420 ( 
.A(n_1195),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1224),
.B(n_1229),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1295),
.A2(n_1239),
.B1(n_1238),
.B2(n_976),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1212),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1239),
.B(n_1238),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_SL g1426 ( 
.A1(n_1315),
.A2(n_1202),
.B(n_1207),
.C(n_1156),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1201),
.A2(n_1291),
.B(n_1186),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1295),
.A2(n_1315),
.B1(n_976),
.B2(n_1005),
.Y(n_1429)
);

AOI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1190),
.A2(n_1255),
.B(n_1191),
.Y(n_1430)
);

AO31x2_ASAP7_75t_L g1431 ( 
.A1(n_1251),
.A2(n_1255),
.A3(n_1265),
.B(n_1191),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1306),
.A2(n_1328),
.B(n_1293),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_SL g1433 ( 
.A1(n_1260),
.A2(n_1133),
.B(n_1204),
.Y(n_1433)
);

INVx6_ASAP7_75t_L g1434 ( 
.A(n_1193),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1201),
.A2(n_1291),
.B(n_1186),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1212),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1203),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1327),
.B(n_1233),
.Y(n_1441)
);

AOI21xp33_ASAP7_75t_L g1442 ( 
.A1(n_1295),
.A2(n_976),
.B(n_1005),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1212),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1445)
);

CKINVDCx16_ASAP7_75t_R g1446 ( 
.A(n_1269),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1447)
);

OAI21xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1295),
.A2(n_742),
.B(n_1122),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1315),
.A2(n_1312),
.B(n_1005),
.C(n_1257),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1212),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1295),
.A2(n_1315),
.B1(n_976),
.B2(n_1005),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1185),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1244),
.B(n_1245),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1193),
.Y(n_1455)
);

BUFx8_ASAP7_75t_SL g1456 ( 
.A(n_1249),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1224),
.B(n_1229),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_SL g1458 ( 
.A1(n_1260),
.A2(n_1133),
.B(n_1204),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1256),
.A2(n_791),
.B1(n_976),
.B2(n_405),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1212),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1295),
.A2(n_1315),
.B1(n_976),
.B2(n_1005),
.Y(n_1462)
);

AOI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1315),
.A2(n_1113),
.B1(n_976),
.B2(n_1295),
.C(n_648),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1209),
.A2(n_1125),
.B1(n_976),
.B2(n_1262),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1306),
.A2(n_1328),
.B(n_1293),
.Y(n_1466)
);

AOI222xp33_ASAP7_75t_L g1467 ( 
.A1(n_1209),
.A2(n_791),
.B1(n_941),
.B2(n_816),
.C1(n_1110),
.C2(n_558),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1212),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1186),
.A2(n_1299),
.B(n_1291),
.Y(n_1469)
);

CKINVDCx11_ASAP7_75t_R g1470 ( 
.A(n_1193),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1335),
.B(n_1402),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1429),
.A2(n_1451),
.B(n_1462),
.C(n_1442),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1403),
.B(n_1409),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1361),
.A2(n_1354),
.B(n_1412),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1425),
.B(n_1365),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1421),
.B(n_1457),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1338),
.B(n_1454),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1330),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1470),
.Y(n_1479)
);

AOI21x1_ASAP7_75t_SL g1480 ( 
.A1(n_1342),
.A2(n_1441),
.B(n_1408),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1460),
.A2(n_1387),
.B1(n_1346),
.B2(n_1446),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1460),
.A2(n_1346),
.B1(n_1465),
.B2(n_1419),
.Y(n_1482)
);

O2A1O1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1467),
.A2(n_1449),
.B(n_1415),
.C(n_1426),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1345),
.B(n_1391),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1418),
.B(n_1359),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1371),
.A2(n_1374),
.B1(n_1418),
.B2(n_1379),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1388),
.A2(n_1384),
.B(n_1354),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1422),
.B(n_1463),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1387),
.A2(n_1419),
.B1(n_1465),
.B2(n_1414),
.Y(n_1489)
);

AO21x1_ASAP7_75t_L g1490 ( 
.A1(n_1449),
.A2(n_1422),
.B(n_1341),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1348),
.B(n_1347),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1362),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1440),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1348),
.B(n_1415),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1357),
.B(n_1375),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1341),
.A2(n_1370),
.B(n_1368),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1426),
.A2(n_1350),
.B(n_1448),
.C(n_1343),
.Y(n_1497)
);

A2O1A1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1370),
.A2(n_1466),
.B(n_1432),
.C(n_1412),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1375),
.B(n_1373),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1373),
.B(n_1372),
.Y(n_1500)
);

AND2x2_ASAP7_75t_SL g1501 ( 
.A(n_1367),
.B(n_1380),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1372),
.B(n_1367),
.Y(n_1502)
);

OR2x6_ASAP7_75t_L g1503 ( 
.A(n_1374),
.B(n_1433),
.Y(n_1503)
);

BUFx2_ASAP7_75t_SL g1504 ( 
.A(n_1334),
.Y(n_1504)
);

NOR2xp67_ASAP7_75t_L g1505 ( 
.A(n_1383),
.B(n_1386),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1368),
.A2(n_1443),
.B1(n_1468),
.B2(n_1450),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1434),
.Y(n_1507)
);

O2A1O1Ixp5_ASAP7_75t_L g1508 ( 
.A1(n_1376),
.A2(n_1369),
.B(n_1349),
.C(n_1385),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1458),
.A2(n_1349),
.B(n_1377),
.C(n_1390),
.Y(n_1509)
);

NOR2xp67_ASAP7_75t_L g1510 ( 
.A(n_1386),
.B(n_1378),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1407),
.A2(n_1437),
.B1(n_1461),
.B2(n_1423),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1380),
.B(n_1366),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1397),
.B(n_1416),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1434),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1392),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1389),
.B(n_1377),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1344),
.B(n_1351),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1351),
.B(n_1374),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1404),
.B(n_1431),
.Y(n_1519)
);

A2O1A1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1364),
.A2(n_1400),
.B(n_1420),
.C(n_1398),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1356),
.A2(n_1455),
.B1(n_1420),
.B2(n_1393),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1396),
.Y(n_1522)
);

O2A1O1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1353),
.A2(n_1356),
.B(n_1405),
.C(n_1413),
.Y(n_1523)
);

AOI31xp33_ASAP7_75t_L g1524 ( 
.A1(n_1353),
.A2(n_1358),
.A3(n_1394),
.B(n_1395),
.Y(n_1524)
);

O2A1O1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1356),
.A2(n_1405),
.B(n_1413),
.C(n_1336),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1410),
.A2(n_1435),
.B(n_1427),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1470),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1410),
.A2(n_1435),
.B(n_1427),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1360),
.B(n_1453),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1355),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1331),
.A2(n_1332),
.B(n_1464),
.Y(n_1531)
);

AOI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1336),
.A2(n_1381),
.B1(n_1417),
.B2(n_1339),
.C(n_1399),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1404),
.B(n_1431),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1401),
.A2(n_1469),
.B(n_1438),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1406),
.A2(n_1459),
.B(n_1436),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1456),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1363),
.B(n_1404),
.Y(n_1537)
);

O2A1O1Ixp5_ASAP7_75t_L g1538 ( 
.A1(n_1430),
.A2(n_1382),
.B(n_1381),
.C(n_1352),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1339),
.A2(n_1417),
.B1(n_1358),
.B2(n_1382),
.C(n_1352),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1411),
.B(n_1424),
.Y(n_1540)
);

O2A1O1Ixp5_ASAP7_75t_L g1541 ( 
.A1(n_1428),
.A2(n_1439),
.B(n_1444),
.C(n_1445),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1447),
.A2(n_1295),
.B(n_1315),
.C(n_1463),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1452),
.B(n_1338),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1361),
.A2(n_1354),
.B(n_1412),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1460),
.A2(n_1295),
.B1(n_1346),
.B2(n_1340),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1338),
.B(n_1454),
.Y(n_1546)
);

A2O1A1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1463),
.A2(n_1295),
.B(n_1315),
.C(n_976),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1460),
.A2(n_1295),
.B1(n_1346),
.B2(n_1340),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1338),
.B(n_1454),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1361),
.A2(n_1354),
.B(n_1412),
.Y(n_1550)
);

OA22x2_ASAP7_75t_L g1551 ( 
.A1(n_1340),
.A2(n_1295),
.B1(n_1345),
.B2(n_1257),
.Y(n_1551)
);

CKINVDCx16_ASAP7_75t_R g1552 ( 
.A(n_1446),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1460),
.A2(n_1295),
.B1(n_1346),
.B2(n_1340),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1342),
.B(n_1408),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1342),
.B(n_1408),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1460),
.A2(n_1295),
.B1(n_1346),
.B2(n_1340),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1337),
.B(n_1333),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1340),
.A2(n_1295),
.B1(n_1460),
.B2(n_1315),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1429),
.A2(n_1315),
.B(n_1267),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1374),
.B(n_1341),
.Y(n_1560)
);

OA21x2_ASAP7_75t_L g1561 ( 
.A1(n_1388),
.A2(n_1384),
.B(n_1354),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1340),
.A2(n_1295),
.B1(n_1460),
.B2(n_1315),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1337),
.B(n_1333),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1338),
.B(n_1454),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1470),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1335),
.B(n_1402),
.Y(n_1566)
);

BUFx12f_ASAP7_75t_L g1567 ( 
.A(n_1470),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1361),
.A2(n_1354),
.B(n_1412),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1429),
.A2(n_1315),
.B(n_1462),
.C(n_1451),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1330),
.Y(n_1570)
);

INVx6_ASAP7_75t_L g1571 ( 
.A(n_1434),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1361),
.A2(n_1354),
.B(n_1412),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1335),
.B(n_1402),
.Y(n_1573)
);

A2O1A1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1463),
.A2(n_1295),
.B(n_1315),
.C(n_976),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1335),
.B(n_1402),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1337),
.B(n_1333),
.Y(n_1576)
);

AO21x2_ASAP7_75t_L g1577 ( 
.A1(n_1474),
.A2(n_1550),
.B(n_1544),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1500),
.B(n_1502),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1537),
.B(n_1519),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_1536),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1485),
.B(n_1499),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1533),
.B(n_1518),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1515),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1522),
.Y(n_1584)
);

OR2x6_ASAP7_75t_L g1585 ( 
.A(n_1568),
.B(n_1572),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1494),
.B(n_1488),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1526),
.A2(n_1528),
.B(n_1525),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1543),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1487),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1503),
.B(n_1520),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1498),
.B(n_1517),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1539),
.B(n_1561),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1510),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1478),
.Y(n_1594)
);

AO22x1_ASAP7_75t_L g1595 ( 
.A1(n_1545),
.A2(n_1556),
.B1(n_1553),
.B2(n_1548),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1484),
.B(n_1475),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1531),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1560),
.B(n_1510),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1492),
.Y(n_1599)
);

BUFx4f_ASAP7_75t_SL g1600 ( 
.A(n_1567),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1534),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1534),
.Y(n_1602)
);

AOI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1505),
.A2(n_1540),
.B(n_1490),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1535),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1538),
.B(n_1501),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1471),
.B(n_1473),
.Y(n_1606)
);

CKINVDCx11_ASAP7_75t_R g1607 ( 
.A(n_1479),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1503),
.B(n_1521),
.Y(n_1608)
);

AO21x2_ASAP7_75t_L g1609 ( 
.A1(n_1523),
.A2(n_1496),
.B(n_1542),
.Y(n_1609)
);

OA21x2_ASAP7_75t_L g1610 ( 
.A1(n_1508),
.A2(n_1541),
.B(n_1532),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1570),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1472),
.A2(n_1559),
.B(n_1524),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1511),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1511),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1506),
.B(n_1477),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1506),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1524),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1566),
.B(n_1573),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1569),
.A2(n_1483),
.B(n_1574),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1486),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1491),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1546),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1516),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1497),
.B(n_1509),
.Y(n_1624)
);

AO21x2_ASAP7_75t_L g1625 ( 
.A1(n_1547),
.A2(n_1558),
.B(n_1562),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1549),
.B(n_1564),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1495),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1551),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1486),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1545),
.A2(n_1556),
.B1(n_1553),
.B2(n_1548),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1530),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1529),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1512),
.B(n_1482),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1575),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1513),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1493),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1554),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1630),
.A2(n_1625),
.B1(n_1619),
.B2(n_1481),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1590),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1588),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1578),
.B(n_1576),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1583),
.Y(n_1642)
);

OAI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1630),
.A2(n_1489),
.B1(n_1514),
.B2(n_1565),
.C(n_1479),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1602),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1582),
.B(n_1514),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1582),
.B(n_1552),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1583),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1597),
.Y(n_1648)
);

AOI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1595),
.A2(n_1557),
.B1(n_1563),
.B2(n_1476),
.C(n_1565),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1597),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1579),
.B(n_1577),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1578),
.B(n_1554),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1585),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1584),
.Y(n_1654)
);

OAI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1619),
.A2(n_1624),
.B1(n_1628),
.B2(n_1633),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1616),
.B(n_1605),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1584),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1625),
.A2(n_1624),
.B1(n_1628),
.B2(n_1595),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1593),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1625),
.B(n_1507),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1605),
.B(n_1555),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1585),
.B(n_1601),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1585),
.B(n_1527),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1601),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1582),
.B(n_1504),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1585),
.B(n_1527),
.Y(n_1666)
);

AOI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1603),
.A2(n_1480),
.B(n_1571),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1638),
.A2(n_1625),
.B1(n_1624),
.B2(n_1628),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1654),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1659),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1654),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1638),
.A2(n_1624),
.B1(n_1628),
.B2(n_1633),
.Y(n_1672)
);

NOR4xp25_ASAP7_75t_SL g1673 ( 
.A(n_1643),
.B(n_1620),
.C(n_1617),
.D(n_1631),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1659),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_1667),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1665),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1655),
.B(n_1593),
.Y(n_1677)
);

OA21x2_ASAP7_75t_L g1678 ( 
.A1(n_1648),
.A2(n_1587),
.B(n_1601),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1661),
.B(n_1608),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1649),
.B(n_1586),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1654),
.Y(n_1681)
);

AOI33xp33_ASAP7_75t_L g1682 ( 
.A1(n_1658),
.A2(n_1620),
.A3(n_1623),
.B1(n_1592),
.B2(n_1627),
.B3(n_1634),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1657),
.Y(n_1683)
);

AOI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1643),
.A2(n_1581),
.B1(n_1586),
.B2(n_1629),
.C(n_1623),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1639),
.B(n_1590),
.Y(n_1685)
);

AOI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1667),
.A2(n_1603),
.B(n_1629),
.Y(n_1686)
);

AOI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1643),
.A2(n_1581),
.B1(n_1623),
.B2(n_1627),
.C(n_1634),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1645),
.B(n_1621),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1639),
.B(n_1590),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1645),
.B(n_1621),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1657),
.Y(n_1691)
);

OAI221xp5_ASAP7_75t_SL g1692 ( 
.A1(n_1658),
.A2(n_1624),
.B1(n_1633),
.B2(n_1649),
.C(n_1591),
.Y(n_1692)
);

OAI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1649),
.A2(n_1624),
.B1(n_1627),
.B2(n_1591),
.C(n_1596),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1657),
.Y(n_1694)
);

OAI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1646),
.A2(n_1617),
.B1(n_1596),
.B2(n_1591),
.Y(n_1695)
);

OAI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1646),
.A2(n_1598),
.B1(n_1606),
.B2(n_1618),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1646),
.A2(n_1606),
.B1(n_1618),
.B2(n_1622),
.C(n_1626),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1642),
.Y(n_1698)
);

AO21x2_ASAP7_75t_L g1699 ( 
.A1(n_1662),
.A2(n_1587),
.B(n_1604),
.Y(n_1699)
);

OAI211xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1660),
.A2(n_1622),
.B(n_1632),
.C(n_1607),
.Y(n_1700)
);

AOI33xp33_ASAP7_75t_L g1701 ( 
.A1(n_1651),
.A2(n_1592),
.A3(n_1615),
.B1(n_1632),
.B2(n_1614),
.B3(n_1613),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1642),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1659),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1641),
.A2(n_1652),
.B1(n_1598),
.B2(n_1665),
.Y(n_1704)
);

CKINVDCx16_ASAP7_75t_R g1705 ( 
.A(n_1639),
.Y(n_1705)
);

OAI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1660),
.A2(n_1626),
.B1(n_1636),
.B2(n_1592),
.C(n_1637),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1645),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1647),
.Y(n_1708)
);

OAI33xp33_ASAP7_75t_L g1709 ( 
.A1(n_1656),
.A2(n_1614),
.A3(n_1635),
.B1(n_1594),
.B2(n_1599),
.B3(n_1611),
.Y(n_1709)
);

NAND4xp25_ASAP7_75t_L g1710 ( 
.A(n_1656),
.B(n_1615),
.C(n_1635),
.D(n_1621),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1669),
.Y(n_1711)
);

INVxp67_ASAP7_75t_SL g1712 ( 
.A(n_1670),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_SL g1713 ( 
.A(n_1673),
.B(n_1666),
.C(n_1663),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1678),
.Y(n_1714)
);

INVx4_ASAP7_75t_SL g1715 ( 
.A(n_1675),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1674),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1686),
.A2(n_1589),
.B(n_1644),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1671),
.Y(n_1718)
);

OR2x2_ASAP7_75t_SL g1719 ( 
.A(n_1705),
.B(n_1653),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1685),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1678),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1681),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1710),
.B(n_1656),
.Y(n_1723)
);

AOI21xp33_ASAP7_75t_L g1724 ( 
.A1(n_1677),
.A2(n_1612),
.B(n_1609),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1683),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1679),
.B(n_1651),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1685),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1701),
.B(n_1663),
.Y(n_1728)
);

AOI21x1_ASAP7_75t_L g1729 ( 
.A1(n_1677),
.A2(n_1664),
.B(n_1650),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1680),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1691),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1685),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1694),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1698),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1703),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1702),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1697),
.B(n_1641),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1708),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1688),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1684),
.B(n_1610),
.C(n_1653),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1679),
.B(n_1651),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1690),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1711),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1726),
.B(n_1741),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1721),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1721),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1719),
.B(n_1707),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1730),
.B(n_1701),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1730),
.A2(n_1612),
.B1(n_1609),
.B2(n_1653),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1718),
.Y(n_1751)
);

AO21x2_ASAP7_75t_L g1752 ( 
.A1(n_1740),
.A2(n_1699),
.B(n_1680),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1737),
.B(n_1682),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1718),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1722),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1723),
.B(n_1704),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1737),
.B(n_1600),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1721),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1721),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1716),
.Y(n_1760)
);

NOR2xp67_ASAP7_75t_L g1761 ( 
.A(n_1713),
.B(n_1706),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1722),
.Y(n_1762)
);

NAND3xp33_ASAP7_75t_L g1763 ( 
.A(n_1740),
.B(n_1668),
.C(n_1692),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1725),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1727),
.B(n_1676),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1715),
.B(n_1689),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1727),
.B(n_1676),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1731),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1719),
.B(n_1640),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1714),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1727),
.B(n_1689),
.Y(n_1771)
);

INVxp67_ASAP7_75t_SL g1772 ( 
.A(n_1716),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1733),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1720),
.B(n_1689),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1714),
.Y(n_1775)
);

OAI211xp5_ASAP7_75t_L g1776 ( 
.A1(n_1724),
.A2(n_1668),
.B(n_1687),
.C(n_1693),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1734),
.B(n_1682),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1733),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1734),
.B(n_1736),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1720),
.B(n_1675),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1780),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1756),
.B(n_1719),
.Y(n_1782)
);

OAI21xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1753),
.A2(n_1728),
.B(n_1732),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1760),
.Y(n_1784)
);

NAND2x1p5_ASAP7_75t_L g1785 ( 
.A(n_1769),
.B(n_1735),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1760),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1743),
.Y(n_1787)
);

NAND2x1p5_ASAP7_75t_L g1788 ( 
.A(n_1769),
.B(n_1735),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1757),
.B(n_1753),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1756),
.B(n_1723),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1748),
.B(n_1712),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1766),
.B(n_1715),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1766),
.B(n_1732),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1748),
.B(n_1712),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1772),
.B(n_1736),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1743),
.Y(n_1796)
);

OR2x2_ASAP7_75t_SL g1797 ( 
.A(n_1763),
.B(n_1713),
.Y(n_1797)
);

OAI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1763),
.A2(n_1724),
.B1(n_1672),
.B2(n_1728),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1777),
.B(n_1723),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1761),
.A2(n_1729),
.B(n_1666),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1749),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1777),
.B(n_1739),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1780),
.Y(n_1803)
);

BUFx2_ASAP7_75t_L g1804 ( 
.A(n_1766),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1749),
.Y(n_1805)
);

OAI31xp33_ASAP7_75t_L g1806 ( 
.A1(n_1776),
.A2(n_1700),
.A3(n_1695),
.B(n_1696),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1772),
.B(n_1738),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1747),
.B(n_1739),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1747),
.B(n_1742),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1766),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1751),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1766),
.Y(n_1812)
);

CKINVDCx16_ASAP7_75t_R g1813 ( 
.A(n_1747),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1776),
.B(n_1607),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1751),
.Y(n_1815)
);

NOR2x1_ASAP7_75t_L g1816 ( 
.A(n_1752),
.B(n_1580),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1745),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1754),
.B(n_1738),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1765),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1816),
.B(n_1752),
.Y(n_1820)
);

AOI222xp33_ASAP7_75t_L g1821 ( 
.A1(n_1814),
.A2(n_1761),
.B1(n_1750),
.B2(n_1600),
.C1(n_1709),
.C2(n_1779),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1784),
.B(n_1754),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1810),
.B(n_1752),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1785),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1791),
.B(n_1779),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1813),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1806),
.B(n_1769),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1786),
.B(n_1755),
.Y(n_1828)
);

INVx1_ASAP7_75t_SL g1829 ( 
.A(n_1804),
.Y(n_1829)
);

AND2x6_ASAP7_75t_L g1830 ( 
.A(n_1792),
.B(n_1527),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1810),
.B(n_1812),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1792),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1812),
.B(n_1752),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1785),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1793),
.B(n_1744),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1788),
.B(n_1744),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1787),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1788),
.B(n_1744),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1796),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1801),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1797),
.B(n_1755),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1781),
.Y(n_1842)
);

OAI21x1_ASAP7_75t_L g1843 ( 
.A1(n_1800),
.A2(n_1729),
.B(n_1717),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1803),
.B(n_1774),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1814),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1805),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1817),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1832),
.B(n_1842),
.Y(n_1848)
);

AOI21xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1827),
.A2(n_1798),
.B(n_1789),
.Y(n_1849)
);

OAI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1826),
.A2(n_1798),
.B1(n_1782),
.B2(n_1799),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1842),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1826),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1845),
.A2(n_1789),
.B1(n_1783),
.B2(n_1791),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1829),
.B(n_1819),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1821),
.B(n_1808),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1832),
.B(n_1771),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1845),
.A2(n_1794),
.B1(n_1802),
.B2(n_1612),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1829),
.B(n_1845),
.Y(n_1858)
);

OAI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1841),
.A2(n_1794),
.B1(n_1790),
.B2(n_1809),
.C(n_1795),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1831),
.B(n_1771),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1836),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1842),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1841),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1836),
.Y(n_1864)
);

AOI211xp5_ASAP7_75t_L g1865 ( 
.A1(n_1841),
.A2(n_1795),
.B(n_1807),
.C(n_1811),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1847),
.Y(n_1866)
);

OAI322xp33_ASAP7_75t_L g1867 ( 
.A1(n_1825),
.A2(n_1807),
.A3(n_1815),
.B1(n_1818),
.B2(n_1817),
.C1(n_1762),
.C2(n_1778),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1820),
.A2(n_1729),
.B(n_1818),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1821),
.A2(n_1653),
.B1(n_1609),
.B2(n_1771),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1820),
.A2(n_1765),
.B1(n_1767),
.B2(n_1732),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1852),
.B(n_1835),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1848),
.B(n_1861),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1848),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1853),
.B(n_1835),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1848),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1858),
.B(n_1835),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1849),
.B(n_1861),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1851),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1854),
.B(n_1825),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1863),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1864),
.B(n_1835),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1860),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1864),
.B(n_1835),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1850),
.A2(n_1820),
.B1(n_1836),
.B2(n_1838),
.Y(n_1884)
);

AOI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1884),
.A2(n_1859),
.B1(n_1855),
.B2(n_1863),
.C(n_1865),
.Y(n_1885)
);

NAND4xp25_ASAP7_75t_SL g1886 ( 
.A(n_1874),
.B(n_1869),
.C(n_1857),
.D(n_1870),
.Y(n_1886)
);

NAND4xp25_ASAP7_75t_L g1887 ( 
.A(n_1876),
.B(n_1824),
.C(n_1834),
.D(n_1851),
.Y(n_1887)
);

AOI211x1_ASAP7_75t_SL g1888 ( 
.A1(n_1871),
.A2(n_1834),
.B(n_1824),
.C(n_1822),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1879),
.B(n_1824),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1873),
.B(n_1856),
.Y(n_1890)
);

A2O1A1Ixp33_ASAP7_75t_L g1891 ( 
.A1(n_1877),
.A2(n_1868),
.B(n_1834),
.C(n_1843),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1880),
.A2(n_1867),
.B(n_1828),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1880),
.A2(n_1828),
.B(n_1822),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1875),
.B(n_1856),
.Y(n_1894)
);

NAND3xp33_ASAP7_75t_L g1895 ( 
.A(n_1881),
.B(n_1862),
.C(n_1866),
.Y(n_1895)
);

AOI221xp5_ASAP7_75t_L g1896 ( 
.A1(n_1882),
.A2(n_1862),
.B1(n_1846),
.B2(n_1837),
.C(n_1839),
.Y(n_1896)
);

AOI21xp33_ASAP7_75t_L g1897 ( 
.A1(n_1885),
.A2(n_1889),
.B(n_1894),
.Y(n_1897)
);

OAI211xp5_ASAP7_75t_L g1898 ( 
.A1(n_1892),
.A2(n_1883),
.B(n_1878),
.C(n_1866),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1890),
.B(n_1872),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1893),
.B(n_1872),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1895),
.Y(n_1901)
);

AO22x2_ASAP7_75t_L g1902 ( 
.A1(n_1888),
.A2(n_1839),
.B1(n_1846),
.B2(n_1837),
.Y(n_1902)
);

AOI211xp5_ASAP7_75t_L g1903 ( 
.A1(n_1886),
.A2(n_1838),
.B(n_1840),
.C(n_1860),
.Y(n_1903)
);

AOI21xp33_ASAP7_75t_L g1904 ( 
.A1(n_1891),
.A2(n_1831),
.B(n_1840),
.Y(n_1904)
);

OAI21xp33_ASAP7_75t_SL g1905 ( 
.A1(n_1887),
.A2(n_1838),
.B(n_1843),
.Y(n_1905)
);

NOR3xp33_ASAP7_75t_L g1906 ( 
.A(n_1897),
.B(n_1896),
.C(n_1831),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1899),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1900),
.B(n_1901),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1903),
.B(n_1830),
.Y(n_1909)
);

AND2x2_ASAP7_75t_SL g1910 ( 
.A(n_1898),
.B(n_1565),
.Y(n_1910)
);

NOR3xp33_ASAP7_75t_L g1911 ( 
.A(n_1904),
.B(n_1847),
.C(n_1844),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1902),
.B(n_1830),
.Y(n_1912)
);

NOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1905),
.B(n_1847),
.Y(n_1913)
);

OAI211xp5_ASAP7_75t_SL g1914 ( 
.A1(n_1907),
.A2(n_1830),
.B(n_1759),
.C(n_1745),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_SL g1915 ( 
.A1(n_1910),
.A2(n_1830),
.B1(n_1833),
.B2(n_1823),
.Y(n_1915)
);

AND3x2_ASAP7_75t_L g1916 ( 
.A(n_1908),
.B(n_1833),
.C(n_1823),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1906),
.A2(n_1830),
.B1(n_1844),
.B2(n_1823),
.Y(n_1917)
);

AOI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1911),
.A2(n_1833),
.B1(n_1844),
.B2(n_1775),
.C(n_1770),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_R g1919 ( 
.A(n_1909),
.B(n_1580),
.Y(n_1919)
);

OAI22xp5_ASAP7_75t_SL g1920 ( 
.A1(n_1917),
.A2(n_1912),
.B1(n_1913),
.B2(n_1571),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1919),
.B(n_1830),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_L g1922 ( 
.A(n_1914),
.B(n_1780),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1915),
.B(n_1765),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1922),
.B(n_1916),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1920),
.Y(n_1925)
);

NOR3xp33_ASAP7_75t_L g1926 ( 
.A(n_1924),
.B(n_1921),
.C(n_1923),
.Y(n_1926)
);

OAI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1925),
.A2(n_1918),
.B1(n_1775),
.B2(n_1770),
.C(n_1746),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1926),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1927),
.B(n_1830),
.Y(n_1929)
);

NAND2xp33_ASAP7_75t_SL g1930 ( 
.A(n_1928),
.B(n_1929),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1929),
.A2(n_1830),
.B1(n_1770),
.B2(n_1775),
.Y(n_1931)
);

AOI22x1_ASAP7_75t_L g1932 ( 
.A1(n_1930),
.A2(n_1758),
.B1(n_1759),
.B2(n_1745),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1931),
.A2(n_1746),
.B1(n_1758),
.B2(n_1759),
.Y(n_1933)
);

XNOR2xp5_ASAP7_75t_L g1934 ( 
.A(n_1932),
.B(n_1830),
.Y(n_1934)
);

OAI21x1_ASAP7_75t_L g1935 ( 
.A1(n_1934),
.A2(n_1933),
.B(n_1843),
.Y(n_1935)
);

NOR2x1_ASAP7_75t_L g1936 ( 
.A(n_1935),
.B(n_1746),
.Y(n_1936)
);

OAI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1936),
.A2(n_1758),
.B(n_1767),
.Y(n_1937)
);

OAI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1937),
.A2(n_1778),
.B1(n_1762),
.B2(n_1764),
.Y(n_1938)
);

AOI211xp5_ASAP7_75t_L g1939 ( 
.A1(n_1938),
.A2(n_1764),
.B(n_1773),
.C(n_1768),
.Y(n_1939)
);


endmodule