module fake_jpeg_5296_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx5_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx4f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx24_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_5),
.B(n_2),
.Y(n_12)
);

FAx1_ASAP7_75t_SL g13 ( 
.A(n_7),
.B(n_0),
.CI(n_2),
.CON(n_13),
.SN(n_13)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_14),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_0),
.C(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_12),
.A2(n_0),
.B(n_3),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_16),
.A2(n_17),
.B1(n_18),
.B2(n_10),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_6),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_17)
);

AOI22x1_ASAP7_75t_L g18 ( 
.A1(n_9),
.A2(n_11),
.B1(n_6),
.B2(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_16),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_10),
.C(n_9),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_17),
.B1(n_9),
.B2(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_13),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_23),
.B1(n_21),
.B2(n_24),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_30),
.B(n_31),
.Y(n_34)
);

NOR2xp67_ASAP7_75t_R g30 ( 
.A(n_25),
.B(n_14),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_20),
.B1(n_27),
.B2(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_20),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_34),
.Y(n_36)
);


endmodule