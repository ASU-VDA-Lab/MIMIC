module fake_aes_6326_n_1323 (n_120, n_136, n_260, n_155, n_107, n_103, n_157, n_52, n_162, n_114, n_156, n_154, n_50, n_7, n_239, n_222, n_253, n_286, n_3, n_34, n_142, n_273, n_231, n_25, n_9, n_163, n_96, n_204, n_72, n_77, n_90, n_169, n_178, n_214, n_227, n_180, n_250, n_99, n_43, n_73, n_190, n_62, n_167, n_97, n_229, n_133, n_199, n_268, n_33, n_192, n_279, n_4, n_59, n_76, n_6, n_74, n_8, n_61, n_44, n_189, n_216, n_153, n_187, n_226, n_66, n_88, n_46, n_121, n_174, n_240, n_188, n_108, n_161, n_37, n_122, n_165, n_224, n_18, n_247, n_65, n_87, n_207, n_5, n_197, n_81, n_285, n_211, n_85, n_112, n_215, n_264, n_102, n_172, n_283, n_47, n_109, n_198, n_290, n_1, n_201, n_16, n_78, n_95, n_217, n_277, n_40, n_68, n_281, n_105, n_210, n_251, n_36, n_228, n_259, n_11, n_244, n_278, n_115, n_270, n_276, n_225, n_179, n_289, n_208, n_237, n_252, n_15, n_168, n_271, n_139, n_152, n_151, n_71, n_117, n_238, n_176, n_70, n_256, n_288, n_94, n_2, n_194, n_17, n_221, n_58, n_282, n_195, n_113, n_242, n_209, n_241, n_284, n_20, n_84, n_130, n_266, n_12, n_56, n_80, n_223, n_67, n_116, n_292, n_22, n_118, n_19, n_233, n_257, n_275, n_202, n_26, n_203, n_261, n_274, n_243, n_39, n_101, n_98, n_150, n_220, n_235, n_38, n_230, n_245, n_104, n_272, n_291, n_100, n_159, n_24, n_141, n_280, n_35, n_91, n_146, n_160, n_32, n_148, n_149, n_246, n_263, n_93, n_191, n_143, n_134, n_48, n_63, n_255, n_54, n_193, n_232, n_125, n_41, n_147, n_55, n_145, n_185, n_29, n_166, n_218, n_267, n_173, n_181, n_123, n_171, n_219, n_60, n_135, n_138, n_140, n_111, n_10, n_212, n_30, n_13, n_254, n_92, n_75, n_82, n_53, n_183, n_64, n_132, n_69, n_196, n_213, n_175, n_248, n_127, n_128, n_170, n_293, n_83, n_200, n_158, n_205, n_23, n_0, n_126, n_258, n_110, n_249, n_262, n_234, n_184, n_182, n_269, n_119, n_265, n_57, n_51, n_287, n_144, n_106, n_186, n_45, n_42, n_21, n_137, n_236, n_131, n_86, n_27, n_124, n_89, n_177, n_28, n_79, n_129, n_164, n_49, n_206, n_14, n_31, n_1323, n_1321);
input n_120;
input n_136;
input n_260;
input n_155;
input n_107;
input n_103;
input n_157;
input n_52;
input n_162;
input n_114;
input n_156;
input n_154;
input n_50;
input n_7;
input n_239;
input n_222;
input n_253;
input n_286;
input n_3;
input n_34;
input n_142;
input n_273;
input n_231;
input n_25;
input n_9;
input n_163;
input n_96;
input n_204;
input n_72;
input n_77;
input n_90;
input n_169;
input n_178;
input n_214;
input n_227;
input n_180;
input n_250;
input n_99;
input n_43;
input n_73;
input n_190;
input n_62;
input n_167;
input n_97;
input n_229;
input n_133;
input n_199;
input n_268;
input n_33;
input n_192;
input n_279;
input n_4;
input n_59;
input n_76;
input n_6;
input n_74;
input n_8;
input n_61;
input n_44;
input n_189;
input n_216;
input n_153;
input n_187;
input n_226;
input n_66;
input n_88;
input n_46;
input n_121;
input n_174;
input n_240;
input n_188;
input n_108;
input n_161;
input n_37;
input n_122;
input n_165;
input n_224;
input n_18;
input n_247;
input n_65;
input n_87;
input n_207;
input n_5;
input n_197;
input n_81;
input n_285;
input n_211;
input n_85;
input n_112;
input n_215;
input n_264;
input n_102;
input n_172;
input n_283;
input n_47;
input n_109;
input n_198;
input n_290;
input n_1;
input n_201;
input n_16;
input n_78;
input n_95;
input n_217;
input n_277;
input n_40;
input n_68;
input n_281;
input n_105;
input n_210;
input n_251;
input n_36;
input n_228;
input n_259;
input n_11;
input n_244;
input n_278;
input n_115;
input n_270;
input n_276;
input n_225;
input n_179;
input n_289;
input n_208;
input n_237;
input n_252;
input n_15;
input n_168;
input n_271;
input n_139;
input n_152;
input n_151;
input n_71;
input n_117;
input n_238;
input n_176;
input n_70;
input n_256;
input n_288;
input n_94;
input n_2;
input n_194;
input n_17;
input n_221;
input n_58;
input n_282;
input n_195;
input n_113;
input n_242;
input n_209;
input n_241;
input n_284;
input n_20;
input n_84;
input n_130;
input n_266;
input n_12;
input n_56;
input n_80;
input n_223;
input n_67;
input n_116;
input n_292;
input n_22;
input n_118;
input n_19;
input n_233;
input n_257;
input n_275;
input n_202;
input n_26;
input n_203;
input n_261;
input n_274;
input n_243;
input n_39;
input n_101;
input n_98;
input n_150;
input n_220;
input n_235;
input n_38;
input n_230;
input n_245;
input n_104;
input n_272;
input n_291;
input n_100;
input n_159;
input n_24;
input n_141;
input n_280;
input n_35;
input n_91;
input n_146;
input n_160;
input n_32;
input n_148;
input n_149;
input n_246;
input n_263;
input n_93;
input n_191;
input n_143;
input n_134;
input n_48;
input n_63;
input n_255;
input n_54;
input n_193;
input n_232;
input n_125;
input n_41;
input n_147;
input n_55;
input n_145;
input n_185;
input n_29;
input n_166;
input n_218;
input n_267;
input n_173;
input n_181;
input n_123;
input n_171;
input n_219;
input n_60;
input n_135;
input n_138;
input n_140;
input n_111;
input n_10;
input n_212;
input n_30;
input n_13;
input n_254;
input n_92;
input n_75;
input n_82;
input n_53;
input n_183;
input n_64;
input n_132;
input n_69;
input n_196;
input n_213;
input n_175;
input n_248;
input n_127;
input n_128;
input n_170;
input n_293;
input n_83;
input n_200;
input n_158;
input n_205;
input n_23;
input n_0;
input n_126;
input n_258;
input n_110;
input n_249;
input n_262;
input n_234;
input n_184;
input n_182;
input n_269;
input n_119;
input n_265;
input n_57;
input n_51;
input n_287;
input n_144;
input n_106;
input n_186;
input n_45;
input n_42;
input n_21;
input n_137;
input n_236;
input n_131;
input n_86;
input n_27;
input n_124;
input n_89;
input n_177;
input n_28;
input n_79;
input n_129;
input n_164;
input n_49;
input n_206;
input n_14;
input n_31;
output n_1323;
output n_1321;
wire n_890;
wire n_107;
wire n_759;
wire n_987;
wire n_658;
wire n_1202;
wire n_309;
wire n_356;
wire n_327;
wire n_1267;
wire n_1041;
wire n_1084;
wire n_169;
wire n_384;
wire n_959;
wire n_1152;
wire n_279;
wire n_1129;
wire n_1149;
wire n_357;
wire n_1207;
wire n_886;
wire n_595;
wire n_875;
wire n_952;
wire n_47;
wire n_766;
wire n_744;
wire n_399;
wire n_942;
wire n_295;
wire n_139;
wire n_151;
wire n_900;
wire n_869;
wire n_935;
wire n_359;
wire n_300;
wire n_487;
wire n_405;
wire n_482;
wire n_1050;
wire n_707;
wire n_220;
wire n_159;
wire n_301;
wire n_340;
wire n_963;
wire n_1278;
wire n_246;
wire n_676;
wire n_143;
wire n_446;
wire n_402;
wire n_54;
wire n_876;
wire n_1198;
wire n_145;
wire n_166;
wire n_1059;
wire n_621;
wire n_981;
wire n_213;
wire n_196;
wire n_1167;
wire n_1089;
wire n_1286;
wire n_1045;
wire n_424;
wire n_110;
wire n_1019;
wire n_1024;
wire n_433;
wire n_660;
wire n_392;
wire n_155;
wire n_1171;
wire n_331;
wire n_814;
wire n_678;
wire n_991;
wire n_1091;
wire n_133;
wire n_1244;
wire n_548;
wire n_443;
wire n_304;
wire n_682;
wire n_441;
wire n_868;
wire n_920;
wire n_517;
wire n_386;
wire n_1209;
wire n_653;
wire n_351;
wire n_1;
wire n_1218;
wire n_829;
wire n_984;
wire n_366;
wire n_837;
wire n_549;
wire n_720;
wire n_1092;
wire n_17;
wire n_711;
wire n_221;
wire n_773;
wire n_266;
wire n_1311;
wire n_793;
wire n_679;
wire n_684;
wire n_879;
wire n_544;
wire n_275;
wire n_691;
wire n_1122;
wire n_274;
wire n_1110;
wire n_38;
wire n_965;
wire n_100;
wire n_1277;
wire n_844;
wire n_695;
wire n_344;
wire n_878;
wire n_367;
wire n_795;
wire n_687;
wire n_212;
wire n_1203;
wire n_254;
wire n_728;
wire n_704;
wire n_435;
wire n_841;
wire n_69;
wire n_1021;
wire n_1186;
wire n_1300;
wire n_1012;
wire n_124;
wire n_1175;
wire n_1127;
wire n_904;
wire n_1016;
wire n_103;
wire n_253;
wire n_677;
wire n_692;
wire n_951;
wire n_163;
wire n_77;
wire n_214;
wire n_167;
wire n_1134;
wire n_76;
wire n_1320;
wire n_470;
wire n_61;
wire n_355;
wire n_153;
wire n_216;
wire n_1066;
wire n_286;
wire n_408;
wire n_1003;
wire n_247;
wire n_1090;
wire n_165;
wire n_413;
wire n_1126;
wire n_290;
wire n_1031;
wire n_792;
wire n_277;
wire n_885;
wire n_631;
wire n_854;
wire n_523;
wire n_985;
wire n_901;
wire n_419;
wire n_1183;
wire n_519;
wire n_271;
wire n_1132;
wire n_785;
wire n_1137;
wire n_94;
wire n_1085;
wire n_997;
wire n_858;
wire n_1191;
wire n_58;
wire n_242;
wire n_284;
wire n_321;
wire n_811;
wire n_734;
wire n_233;
wire n_698;
wire n_257;
wire n_26;
wire n_1173;
wire n_477;
wire n_318;
wire n_98;
wire n_714;
wire n_32;
wire n_531;
wire n_406;
wire n_372;
wire n_820;
wire n_923;
wire n_702;
wire n_1301;
wire n_647;
wire n_445;
wire n_1303;
wire n_732;
wire n_926;
wire n_845;
wire n_10;
wire n_1036;
wire n_761;
wire n_1075;
wire n_510;
wire n_360;
wire n_1040;
wire n_1067;
wire n_296;
wire n_975;
wire n_89;
wire n_130;
wire n_639;
wire n_1008;
wire n_34;
wire n_395;
wire n_250;
wire n_1120;
wire n_565;
wire n_323;
wire n_1101;
wire n_1275;
wire n_240;
wire n_768;
wire n_568;
wire n_1287;
wire n_46;
wire n_174;
wire n_108;
wire n_335;
wire n_37;
wire n_515;
wire n_802;
wire n_672;
wire n_87;
wire n_466;
wire n_1027;
wire n_572;
wire n_81;
wire n_1292;
wire n_36;
wire n_917;
wire n_680;
wire n_767;
wire n_237;
wire n_1034;
wire n_633;
wire n_803;
wire n_398;
wire n_796;
wire n_1263;
wire n_662;
wire n_391;
wire n_241;
wire n_874;
wire n_449;
wire n_1070;
wire n_56;
wire n_455;
wire n_67;
wire n_401;
wire n_1159;
wire n_877;
wire n_725;
wire n_930;
wire n_1318;
wire n_1063;
wire n_291;
wire n_1233;
wire n_664;
wire n_35;
wire n_1196;
wire n_659;
wire n_968;
wire n_1093;
wire n_336;
wire n_1241;
wire n_556;
wire n_648;
wire n_60;
wire n_936;
wire n_1289;
wire n_924;
wire n_305;
wire n_1158;
wire n_358;
wire n_627;
wire n_750;
wire n_589;
wire n_128;
wire n_697;
wire n_642;
wire n_234;
wire n_848;
wire n_1005;
wire n_1153;
wire n_514;
wire n_625;
wire n_403;
wire n_995;
wire n_738;
wire n_511;
wire n_49;
wire n_646;
wire n_156;
wire n_154;
wire n_1099;
wire n_994;
wire n_1257;
wire n_204;
wire n_439;
wire n_180;
wire n_73;
wire n_1172;
wire n_74;
wire n_308;
wire n_518;
wire n_681;
wire n_189;
wire n_447;
wire n_903;
wire n_66;
wire n_379;
wire n_626;
wire n_475;
wire n_281;
wire n_1296;
wire n_516;
wire n_1282;
wire n_342;
wire n_557;
wire n_438;
wire n_461;
wire n_830;
wire n_562;
wire n_967;
wire n_526;
wire n_261;
wire n_104;
wire n_709;
wire n_1200;
wire n_821;
wire n_468;
wire n_91;
wire n_148;
wire n_378;
wire n_752;
wire n_823;
wire n_191;
wire n_63;
wire n_387;
wire n_961;
wire n_492;
wire n_1100;
wire n_1128;
wire n_219;
wire n_343;
wire n_555;
wire n_1259;
wire n_880;
wire n_312;
wire n_742;
wire n_23;
wire n_1048;
wire n_269;
wire n_751;
wire n_186;
wire n_164;
wire n_114;
wire n_1229;
wire n_50;
wire n_1322;
wire n_574;
wire n_478;
wire n_1225;
wire n_1141;
wire n_998;
wire n_824;
wire n_601;
wire n_736;
wire n_215;
wire n_172;
wire n_979;
wire n_332;
wire n_670;
wire n_1112;
wire n_755;
wire n_1193;
wire n_765;
wire n_179;
wire n_289;
wire n_721;
wire n_485;
wire n_354;
wire n_980;
wire n_70;
wire n_458;
wire n_322;
wire n_1123;
wire n_317;
wire n_800;
wire n_973;
wire n_522;
wire n_1055;
wire n_326;
wire n_532;
wire n_1206;
wire n_635;
wire n_1107;
wire n_1023;
wire n_299;
wire n_1072;
wire n_509;
wire n_1043;
wire n_263;
wire n_1230;
wire n_193;
wire n_267;
wire n_638;
wire n_873;
wire n_450;
wire n_585;
wire n_140;
wire n_779;
wire n_13;
wire n_64;
wire n_970;
wire n_921;
wire n_927;
wire n_339;
wire n_696;
wire n_748;
wire n_774;
wire n_1080;
wire n_1280;
wire n_743;
wire n_944;
wire n_96;
wire n_669;
wire n_770;
wire n_364;
wire n_33;
wire n_464;
wire n_1279;
wire n_1119;
wire n_590;
wire n_121;
wire n_161;
wire n_224;
wire n_537;
wire n_1117;
wire n_843;
wire n_85;
wire n_264;
wire n_733;
wire n_846;
wire n_791;
wire n_1157;
wire n_932;
wire n_244;
wire n_1061;
wire n_297;
wire n_350;
wire n_616;
wire n_208;
wire n_528;
wire n_168;
wire n_1271;
wire n_1011;
wire n_1087;
wire n_758;
wire n_775;
wire n_113;
wire n_498;
wire n_538;
wire n_1214;
wire n_302;
wire n_292;
wire n_547;
wire n_741;
wire n_705;
wire n_828;
wire n_988;
wire n_996;
wire n_1283;
wire n_1164;
wire n_146;
wire n_641;
wire n_93;
wire n_1294;
wire n_41;
wire n_826;
wire n_1009;
wire n_1079;
wire n_898;
wire n_417;
wire n_1215;
wire n_1192;
wire n_1248;
wire n_818;
wire n_1297;
wire n_75;
wire n_82;
wire n_183;
wire n_550;
wire n_582;
wire n_784;
wire n_170;
wire n_915;
wire n_363;
wire n_1078;
wire n_724;
wire n_21;
wire n_1148;
wire n_939;
wire n_640;
wire n_1228;
wire n_976;
wire n_938;
wire n_657;
wire n_964;
wire n_385;
wire n_454;
wire n_227;
wire n_551;
wire n_268;
wire n_190;
wire n_62;
wire n_4;
wire n_956;
wire n_781;
wire n_1071;
wire n_376;
wire n_694;
wire n_88;
wire n_807;
wire n_613;
wire n_207;
wire n_1258;
wire n_1190;
wire n_298;
wire n_630;
wire n_1290;
wire n_983;
wire n_1052;
wire n_78;
wire n_68;
wire n_919;
wire n_598;
wire n_251;
wire n_810;
wire n_916;
wire n_465;
wire n_881;
wire n_520;
wire n_668;
wire n_338;
wire n_907;
wire n_20;
wire n_782;
wire n_832;
wire n_790;
wire n_504;
wire n_456;
wire n_319;
wire n_1227;
wire n_933;
wire n_719;
wire n_788;
wire n_655;
wire n_1208;
wire n_1103;
wire n_472;
wire n_1010;
wire n_1142;
wire n_457;
wire n_255;
wire n_1170;
wire n_513;
wire n_29;
wire n_893;
wire n_382;
wire n_894;
wire n_536;
wire n_474;
wire n_745;
wire n_706;
wire n_1165;
wire n_1210;
wire n_958;
wire n_0;
wire n_619;
wire n_258;
wire n_974;
wire n_1155;
wire n_607;
wire n_184;
wire n_1251;
wire n_144;
wire n_1130;
wire n_420;
wire n_86;
wire n_28;
wire n_206;
wire n_349;
wire n_673;
wire n_1124;
wire n_25;
wire n_592;
wire n_1238;
wire n_545;
wire n_99;
wire n_43;
wire n_199;
wire n_1184;
wire n_831;
wire n_1295;
wire n_729;
wire n_394;
wire n_44;
wire n_352;
wire n_689;
wire n_1268;
wire n_1306;
wire n_316;
wire n_586;
wire n_1252;
wire n_1131;
wire n_645;
wire n_497;
wire n_11;
wire n_1314;
wire n_1088;
wire n_1242;
wire n_1197;
wire n_805;
wire n_1315;
wire n_373;
wire n_753;
wire n_288;
wire n_71;
wire n_176;
wire n_931;
wire n_195;
wire n_723;
wire n_833;
wire n_1281;
wire n_409;
wire n_838;
wire n_534;
wire n_483;
wire n_423;
wire n_353;
wire n_303;
wire n_1187;
wire n_566;
wire n_149;
wire n_567;
wire n_780;
wire n_1224;
wire n_864;
wire n_125;
wire n_596;
wire n_1046;
wire n_1111;
wire n_1243;
wire n_494;
wire n_1115;
wire n_481;
wire n_135;
wire n_797;
wire n_1147;
wire n_127;
wire n_182;
wire n_529;
wire n_656;
wire n_1246;
wire n_1226;
wire n_137;
wire n_1274;
wire n_651;
wire n_882;
wire n_999;
wire n_636;
wire n_614;
wire n_737;
wire n_428;
wire n_178;
wire n_1276;
wire n_708;
wire n_229;
wire n_442;
wire n_1176;
wire n_699;
wire n_857;
wire n_1273;
wire n_1199;
wire n_8;
wire n_1185;
wire n_578;
wire n_928;
wire n_187;
wire n_188;
wire n_18;
wire n_628;
wire n_425;
wire n_905;
wire n_109;
wire n_198;
wire n_1310;
wire n_426;
wire n_716;
wire n_892;
wire n_115;
wire n_476;
wire n_989;
wire n_599;
wire n_1232;
wire n_715;
wire n_849;
wire n_1077;
wire n_404;
wire n_1288;
wire n_362;
wire n_688;
wire n_152;
wire n_1102;
wire n_1177;
wire n_506;
wire n_328;
wire n_1305;
wire n_388;
wire n_1260;
wire n_763;
wire n_632;
wire n_906;
wire n_615;
wire n_1145;
wire n_701;
wire n_888;
wire n_661;
wire n_909;
wire n_493;
wire n_972;
wire n_690;
wire n_272;
wire n_561;
wire n_1057;
wire n_581;
wire n_280;
wire n_1068;
wire n_377;
wire n_1044;
wire n_1013;
wire n_1143;
wire n_185;
wire n_955;
wire n_1007;
wire n_950;
wire n_171;
wire n_899;
wire n_111;
wire n_978;
wire n_30;
wire n_634;
wire n_559;
wire n_407;
wire n_527;
wire n_200;
wire n_986;
wire n_262;
wire n_503;
wire n_969;
wire n_1138;
wire n_856;
wire n_1081;
wire n_347;
wire n_79;
wire n_1265;
wire n_1284;
wire n_521;
wire n_157;
wire n_808;
wire n_1113;
wire n_1038;
wire n_434;
wire n_624;
wire n_1240;
wire n_273;
wire n_325;
wire n_571;
wire n_524;
wire n_1118;
wire n_530;
wire n_348;
wire n_762;
wire n_685;
wire n_90;
wire n_72;
wire n_594;
wire n_1114;
wire n_1030;
wire n_1253;
wire n_861;
wire n_809;
wire n_908;
wire n_1239;
wire n_1022;
wire n_463;
wire n_1125;
wire n_484;
wire n_431;
wire n_860;
wire n_710;
wire n_560;
wire n_525;
wire n_1174;
wire n_393;
wire n_211;
wire n_283;
wire n_217;
wire n_1264;
wire n_259;
wire n_1178;
wire n_666;
wire n_276;
wire n_225;
wire n_815;
wire n_922;
wire n_839;
wire n_1109;
wire n_739;
wire n_1221;
wire n_501;
wire n_593;
wire n_597;
wire n_1097;
wire n_1234;
wire n_1151;
wire n_203;
wire n_460;
wire n_1235;
wire n_637;
wire n_957;
wire n_872;
wire n_539;
wire n_713;
wire n_467;
wire n_760;
wire n_665;
wire n_390;
wire n_1001;
wire n_1161;
wire n_1321;
wire n_778;
wire n_925;
wire n_158;
wire n_249;
wire n_749;
wire n_1069;
wire n_1098;
wire n_106;
wire n_605;
wire n_835;
wire n_437;
wire n_940;
wire n_1150;
wire n_700;
wire n_1033;
wire n_1236;
wire n_822;
wire n_381;
wire n_142;
wire n_754;
wire n_453;
wire n_59;
wire n_1121;
wire n_914;
wire n_945;
wire n_852;
wire n_122;
wire n_374;
wire n_1042;
wire n_197;
wire n_541;
wire n_1285;
wire n_112;
wire n_735;
wire n_552;
wire n_962;
wire n_416;
wire n_1299;
wire n_1205;
wire n_414;
wire n_469;
wire n_1313;
wire n_429;
wire n_1270;
wire n_804;
wire n_117;
wire n_238;
wire n_577;
wire n_294;
wire n_2;
wire n_1256;
wire n_412;
wire n_618;
wire n_22;
wire n_683;
wire n_479;
wire n_1266;
wire n_584;
wire n_311;
wire n_813;
wire n_819;
wire n_1096;
wire n_39;
wire n_953;
wire n_489;
wire n_245;
wire n_764;
wire n_486;
wire n_794;
wire n_1261;
wire n_1017;
wire n_1195;
wire n_1291;
wire n_543;
wire n_218;
wire n_173;
wire n_488;
wire n_1105;
wire n_799;
wire n_937;
wire n_462;
wire n_495;
wire n_430;
wire n_418;
wire n_175;
wire n_897;
wire n_512;
wire n_1188;
wire n_265;
wire n_57;
wire n_51;
wire n_1231;
wire n_131;
wire n_27;
wire n_1180;
wire n_448;
wire n_415;
wire n_31;
wire n_1309;
wire n_239;
wire n_7;
wire n_895;
wire n_1029;
wire n_1014;
wire n_929;
wire n_769;
wire n_370;
wire n_1015;
wire n_604;
wire n_440;
wire n_786;
wire n_1249;
wire n_226;
wire n_535;
wire n_1116;
wire n_285;
wire n_564;
wire n_1047;
wire n_471;
wire n_1049;
wire n_949;
wire n_1035;
wire n_1104;
wire n_371;
wire n_579;
wire n_608;
wire n_368;
wire n_1020;
wire n_859;
wire n_223;
wire n_19;
wire n_971;
wire n_569;
wire n_410;
wire n_502;
wire n_1262;
wire n_1312;
wire n_1136;
wire n_1298;
wire n_629;
wire n_1189;
wire n_558;
wire n_181;
wire n_123;
wire n_553;
wire n_817;
wire n_776;
wire n_315;
wire n_397;
wire n_53;
wire n_1201;
wire n_1058;
wire n_836;
wire n_293;
wire n_1028;
wire n_990;
wire n_663;
wire n_887;
wire n_507;
wire n_334;
wire n_1095;
wire n_1062;
wire n_993;
wire n_806;
wire n_120;
wire n_1053;
wire n_650;
wire n_162;
wire n_977;
wire n_772;
wire n_816;
wire n_789;
wire n_1255;
wire n_3;
wire n_330;
wire n_884;
wire n_231;
wire n_1307;
wire n_9;
wire n_1211;
wire n_1083;
wire n_652;
wire n_97;
wire n_982;
wire n_324;
wire n_422;
wire n_192;
wire n_329;
wire n_6;
wire n_1293;
wire n_1160;
wire n_883;
wire n_801;
wire n_912;
wire n_314;
wire n_307;
wire n_934;
wire n_16;
wire n_95;
wire n_40;
wire n_210;
wire n_228;
wire n_863;
wire n_671;
wire n_1144;
wire n_278;
wire n_270;
wire n_1135;
wire n_617;
wire n_396;
wire n_1139;
wire n_851;
wire n_588;
wire n_375;
wire n_1162;
wire n_855;
wire n_911;
wire n_491;
wire n_1216;
wire n_80;
wire n_1237;
wire n_546;
wire n_756;
wire n_992;
wire n_576;
wire n_622;
wire n_910;
wire n_150;
wire n_235;
wire n_533;
wire n_686;
wire n_1269;
wire n_141;
wire n_160;
wire n_1182;
wire n_499;
wire n_757;
wire n_1060;
wire n_232;
wire n_812;
wire n_783;
wire n_147;
wire n_1065;
wire n_644;
wire n_746;
wire n_1064;
wire n_583;
wire n_248;
wire n_866;
wire n_83;
wire n_1106;
wire n_603;
wire n_1032;
wire n_119;
wire n_667;
wire n_1076;
wire n_1018;
wire n_129;
wire n_611;
wire n_421;
wire n_52;
wire n_1179;
wire n_850;
wire n_1308;
wire n_1074;
wire n_787;
wire n_1272;
wire n_1108;
wire n_609;
wire n_946;
wire n_1082;
wire n_65;
wire n_5;
wire n_496;
wire n_1181;
wire n_1316;
wire n_320;
wire n_102;
wire n_201;
wire n_612;
wire n_771;
wire n_827;
wire n_1037;
wire n_747;
wire n_252;
wire n_966;
wire n_693;
wire n_896;
wire n_1212;
wire n_1056;
wire n_194;
wire n_825;
wire n_282;
wire n_1223;
wire n_703;
wire n_1254;
wire n_116;
wire n_1213;
wire n_1247;
wire n_118;
wire n_587;
wire n_554;
wire n_722;
wire n_1245;
wire n_243;
wire n_346;
wire n_1154;
wire n_345;
wire n_230;
wire n_452;
wire n_337;
wire n_726;
wire n_847;
wire n_842;
wire n_918;
wire n_623;
wire n_451;
wire n_500;
wire n_948;
wire n_1026;
wire n_575;
wire n_600;
wire n_731;
wire n_1006;
wire n_132;
wire n_643;
wire n_205;
wire n_126;
wire n_473;
wire n_389;
wire n_834;
wire n_427;
wire n_1194;
wire n_42;
wire n_1086;
wire n_871;
wire n_620;
wire n_480;
wire n_1073;
wire n_1039;
wire n_310;
wire n_341;
wire n_14;
wire n_236;
wire n_727;
wire n_260;
wire n_136;
wire n_891;
wire n_1317;
wire n_1002;
wire n_1004;
wire n_580;
wire n_610;
wire n_222;
wire n_1302;
wire n_853;
wire n_798;
wire n_943;
wire n_606;
wire n_712;
wire n_777;
wire n_954;
wire n_902;
wire n_459;
wire n_717;
wire n_865;
wire n_380;
wire n_867;
wire n_649;
wire n_602;
wire n_444;
wire n_105;
wire n_1220;
wire n_870;
wire n_889;
wire n_432;
wire n_913;
wire n_730;
wire n_369;
wire n_1146;
wire n_361;
wire n_1163;
wire n_654;
wire n_15;
wire n_960;
wire n_256;
wire n_365;
wire n_1222;
wire n_591;
wire n_1025;
wire n_209;
wire n_84;
wire n_12;
wire n_1133;
wire n_1250;
wire n_1169;
wire n_383;
wire n_202;
wire n_542;
wire n_862;
wire n_101;
wire n_1168;
wire n_941;
wire n_1304;
wire n_508;
wire n_24;
wire n_1204;
wire n_490;
wire n_540;
wire n_947;
wire n_840;
wire n_400;
wire n_1094;
wire n_134;
wire n_48;
wire n_563;
wire n_55;
wire n_718;
wire n_1140;
wire n_1156;
wire n_138;
wire n_573;
wire n_505;
wire n_740;
wire n_313;
wire n_92;
wire n_333;
wire n_306;
wire n_675;
wire n_1219;
wire n_1000;
wire n_674;
wire n_570;
wire n_411;
wire n_287;
wire n_45;
wire n_1217;
wire n_177;
wire n_1054;
wire n_1166;
wire n_436;
wire n_1051;
INVx1_ASAP7_75t_SL g294 ( .A(n_6), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_16), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_127), .Y(n_296) );
NOR2xp67_ASAP7_75t_L g297 ( .A(n_74), .B(n_289), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_209), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_70), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_194), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_165), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_290), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_281), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_52), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_243), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_101), .Y(n_306) );
INVxp33_ASAP7_75t_L g307 ( .A(n_110), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_288), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_230), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_87), .Y(n_310) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_129), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_54), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_158), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_16), .Y(n_314) );
CKINVDCx16_ASAP7_75t_R g315 ( .A(n_20), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_20), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_25), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_41), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_244), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_4), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_65), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_49), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_241), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_155), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_166), .Y(n_325) );
CKINVDCx16_ASAP7_75t_R g326 ( .A(n_276), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_75), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_98), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_19), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_106), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_278), .Y(n_331) );
CKINVDCx14_ASAP7_75t_R g332 ( .A(n_121), .Y(n_332) );
INVxp33_ASAP7_75t_L g333 ( .A(n_130), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_179), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_95), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_273), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_126), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_53), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_233), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_71), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_78), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_214), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_254), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_213), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_261), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_275), .B(n_123), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_89), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_133), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_218), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_242), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_34), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_116), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_184), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_154), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_169), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_228), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_204), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_232), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_150), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_60), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_33), .Y(n_361) );
INVxp67_ASAP7_75t_SL g362 ( .A(n_292), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_28), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_138), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_287), .Y(n_365) );
CKINVDCx16_ASAP7_75t_R g366 ( .A(n_239), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_69), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_22), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_76), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_167), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_11), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_37), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_272), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_277), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_279), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_240), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_177), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_252), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_198), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_156), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_74), .Y(n_381) );
BUFx2_ASAP7_75t_SL g382 ( .A(n_70), .Y(n_382) );
INVxp33_ASAP7_75t_L g383 ( .A(n_6), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_128), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_250), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_112), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_248), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_190), .Y(n_388) );
INVxp33_ASAP7_75t_SL g389 ( .A(n_293), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_24), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_19), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_91), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_168), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_122), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_197), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_119), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_81), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_53), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_172), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_79), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_229), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_24), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_152), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_117), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_201), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_134), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_183), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_175), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_124), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g410 ( .A(n_105), .Y(n_410) );
INVxp33_ASAP7_75t_L g411 ( .A(n_4), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_271), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_83), .Y(n_413) );
INVxp33_ASAP7_75t_SL g414 ( .A(n_61), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_15), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_22), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_56), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_46), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_196), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_8), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_108), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_88), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_238), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_13), .Y(n_424) );
INVxp33_ASAP7_75t_SL g425 ( .A(n_3), .Y(n_425) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_262), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_54), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_265), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_264), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_266), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_25), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_39), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_64), .Y(n_433) );
CKINVDCx16_ASAP7_75t_R g434 ( .A(n_77), .Y(n_434) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_160), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_139), .Y(n_436) );
INVxp33_ASAP7_75t_L g437 ( .A(n_171), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_246), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_284), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_207), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_141), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_315), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_415), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_303), .Y(n_444) );
BUFx8_ASAP7_75t_L g445 ( .A(n_303), .Y(n_445) );
INVxp33_ASAP7_75t_SL g446 ( .A(n_299), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_415), .B(n_0), .Y(n_447) );
AND3x2_ASAP7_75t_L g448 ( .A(n_305), .B(n_1), .C(n_2), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_415), .B(n_3), .Y(n_449) );
INVxp33_ASAP7_75t_SL g450 ( .A(n_351), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_303), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_338), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_303), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_363), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_381), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_383), .B(n_411), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_384), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_363), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_384), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_381), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_338), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_368), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_368), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_296), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_326), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_307), .B(n_5), .Y(n_466) );
INVx3_ASAP7_75t_L g467 ( .A(n_309), .Y(n_467) );
OAI22xp5_ASAP7_75t_SL g468 ( .A1(n_418), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_383), .B(n_7), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_298), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_384), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_300), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_384), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_334), .Y(n_474) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_334), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_301), .Y(n_476) );
AND2x6_ASAP7_75t_L g477 ( .A(n_447), .B(n_341), .Y(n_477) );
INVx4_ASAP7_75t_L g478 ( .A(n_447), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_456), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_474), .Y(n_480) );
AND2x6_ASAP7_75t_L g481 ( .A(n_447), .B(n_341), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_456), .B(n_366), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_458), .B(n_379), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_447), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_450), .Y(n_485) );
AND2x6_ASAP7_75t_L g486 ( .A(n_449), .B(n_302), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_445), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_458), .B(n_307), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_445), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_449), .Y(n_490) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_466), .B(n_372), .C(n_312), .Y(n_491) );
AND2x6_ASAP7_75t_L g492 ( .A(n_449), .B(n_308), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_449), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_443), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_474), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_464), .B(n_411), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_443), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_465), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_452), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g500 ( .A(n_464), .B(n_310), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_470), .B(n_333), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_470), .B(n_333), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_472), .B(n_437), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_462), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_474), .Y(n_505) );
AND3x4_ASAP7_75t_L g506 ( .A(n_446), .B(n_297), .C(n_414), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_461), .Y(n_507) );
INVx4_ASAP7_75t_L g508 ( .A(n_454), .Y(n_508) );
AND2x2_ASAP7_75t_SL g509 ( .A(n_466), .B(n_410), .Y(n_509) );
AND2x6_ASAP7_75t_L g510 ( .A(n_454), .B(n_319), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_472), .B(n_437), .Y(n_511) );
INVxp33_ASAP7_75t_L g512 ( .A(n_469), .Y(n_512) );
INVx3_ASAP7_75t_R g513 ( .A(n_444), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_476), .B(n_396), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_454), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_454), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_476), .B(n_358), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_462), .B(n_351), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_474), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_463), .B(n_426), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_463), .B(n_434), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_478), .B(n_323), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_484), .A2(n_467), .B1(n_425), .B2(n_414), .Y(n_523) );
INVx3_ASAP7_75t_L g524 ( .A(n_478), .Y(n_524) );
OR2x6_ASAP7_75t_L g525 ( .A(n_485), .B(n_468), .Y(n_525) );
NOR2x1p5_ASAP7_75t_L g526 ( .A(n_498), .B(n_361), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_514), .B(n_448), .Y(n_527) );
OAI21xp33_ASAP7_75t_L g528 ( .A1(n_512), .A2(n_389), .B(n_304), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_497), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_501), .B(n_306), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_502), .B(n_313), .Y(n_531) );
INVx4_ASAP7_75t_L g532 ( .A(n_487), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_497), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_484), .A2(n_346), .B(n_336), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_487), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_494), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_503), .B(n_313), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_511), .B(n_339), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_496), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_515), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_489), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_498), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_520), .B(n_389), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_479), .B(n_361), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_499), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_488), .B(n_442), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_518), .A2(n_442), .B(n_425), .C(n_455), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_516), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_496), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_504), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_518), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_516), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_480), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_478), .B(n_324), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_514), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_521), .B(n_455), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_514), .B(n_460), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_500), .B(n_325), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_493), .A2(n_467), .B1(n_460), .B2(n_295), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_483), .B(n_339), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_491), .B(n_467), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_483), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_483), .B(n_486), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_493), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_500), .B(n_328), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_486), .B(n_448), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_500), .B(n_335), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_517), .B(n_343), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_480), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_509), .A2(n_344), .B1(n_349), .B2(n_345), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_507), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_482), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_477), .Y(n_573) );
INVx3_ASAP7_75t_L g574 ( .A(n_490), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_505), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_490), .Y(n_576) );
INVx5_ASAP7_75t_L g577 ( .A(n_477), .Y(n_577) );
BUFx3_ASAP7_75t_L g578 ( .A(n_489), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_505), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_519), .Y(n_580) );
OR2x6_ASAP7_75t_L g581 ( .A(n_490), .B(n_468), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_508), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_499), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_519), .Y(n_584) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_495), .Y(n_585) );
O2A1O1Ixp33_ASAP7_75t_L g586 ( .A1(n_506), .A2(n_314), .B(n_317), .C(n_316), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_508), .Y(n_587) );
INVxp67_ASAP7_75t_SL g588 ( .A(n_508), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_477), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_486), .A2(n_467), .B1(n_320), .B2(n_321), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_477), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_477), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_477), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_481), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_486), .B(n_492), .Y(n_595) );
BUFx2_ASAP7_75t_L g596 ( .A(n_481), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g597 ( .A1(n_509), .A2(n_322), .B(n_327), .C(n_318), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_481), .B(n_343), .Y(n_598) );
BUFx2_ASAP7_75t_L g599 ( .A(n_481), .Y(n_599) );
BUFx3_ASAP7_75t_L g600 ( .A(n_486), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_506), .A2(n_345), .B1(n_349), .B2(n_344), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_495), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_481), .B(n_354), .Y(n_603) );
OR2x6_ASAP7_75t_L g604 ( .A(n_486), .B(n_382), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_555), .B(n_492), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_574), .Y(n_606) );
INVx4_ASAP7_75t_L g607 ( .A(n_563), .Y(n_607) );
BUFx12f_ASAP7_75t_L g608 ( .A(n_545), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_574), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_536), .Y(n_610) );
AO22x1_ASAP7_75t_L g611 ( .A1(n_542), .A2(n_492), .B1(n_390), .B2(n_417), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_571), .Y(n_612) );
BUFx2_ASAP7_75t_L g613 ( .A(n_563), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_529), .A2(n_360), .B(n_371), .C(n_340), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_597), .A2(n_391), .B(n_402), .C(n_398), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_542), .Y(n_616) );
A2O1A1Ixp33_ASAP7_75t_L g617 ( .A1(n_533), .A2(n_424), .B(n_431), .C(n_416), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_535), .Y(n_618) );
INVx3_ASAP7_75t_L g619 ( .A(n_532), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_535), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_550), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_522), .A2(n_495), .B(n_362), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_551), .A2(n_492), .B1(n_510), .B2(n_378), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_597), .A2(n_294), .B(n_432), .C(n_418), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_564), .B(n_492), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_527), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_522), .A2(n_495), .B(n_377), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_532), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_544), .B(n_432), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_576), .Y(n_630) );
BUFx8_ASAP7_75t_SL g631 ( .A(n_545), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_524), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_563), .B(n_492), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_581), .A2(n_510), .B1(n_378), .B2(n_413), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_583), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_535), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_524), .Y(n_637) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_535), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_554), .A2(n_435), .B(n_311), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_557), .B(n_510), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_539), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_549), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_570), .B(n_367), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_562), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_557), .A2(n_342), .B(n_347), .C(n_337), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_527), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_552), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_540), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_523), .A2(n_420), .B1(n_417), .B2(n_390), .C(n_367), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_601), .Y(n_650) );
A2O1A1Ixp33_ASAP7_75t_L g651 ( .A1(n_561), .A2(n_350), .B(n_352), .C(n_348), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_546), .B(n_420), .Y(n_652) );
NOR2x1_ASAP7_75t_R g653 ( .A(n_527), .B(n_354), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_590), .A2(n_413), .B1(n_412), .B2(n_433), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_566), .B(n_510), .Y(n_655) );
INVx2_ASAP7_75t_SL g656 ( .A(n_526), .Y(n_656) );
INVx4_ASAP7_75t_L g657 ( .A(n_595), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_540), .Y(n_658) );
AOI21x1_ASAP7_75t_L g659 ( .A1(n_558), .A2(n_357), .B(n_353), .Y(n_659) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_578), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_604), .Y(n_661) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_578), .Y(n_662) );
OR2x6_ASAP7_75t_L g663 ( .A(n_595), .B(n_433), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_548), .Y(n_664) );
INVx4_ASAP7_75t_L g665 ( .A(n_595), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_556), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_572), .B(n_412), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_566), .A2(n_510), .B1(n_445), .B2(n_332), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_523), .A2(n_427), .B1(n_329), .B2(n_439), .C(n_438), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_561), .A2(n_365), .B(n_369), .C(n_359), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_560), .B(n_510), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_532), .B(n_355), .Y(n_672) );
AO21x2_ASAP7_75t_L g673 ( .A1(n_534), .A2(n_565), .B(n_558), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_543), .A2(n_373), .B(n_374), .C(n_370), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_582), .Y(n_675) );
OA22x2_ASAP7_75t_L g676 ( .A1(n_525), .A2(n_356), .B1(n_380), .B2(n_355), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_L g677 ( .A1(n_543), .A2(n_386), .B(n_387), .C(n_385), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_556), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_587), .Y(n_679) );
INVx4_ASAP7_75t_L g680 ( .A(n_604), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_565), .A2(n_393), .B(n_388), .Y(n_681) );
AND2x4_ASAP7_75t_L g682 ( .A(n_566), .B(n_394), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_528), .B(n_356), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_590), .A2(n_397), .B1(n_399), .B2(n_395), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_530), .B(n_380), .Y(n_685) );
NAND2x1_ASAP7_75t_L g686 ( .A(n_604), .B(n_309), .Y(n_686) );
INVx3_ASAP7_75t_L g687 ( .A(n_600), .Y(n_687) );
BUFx12f_ASAP7_75t_L g688 ( .A(n_525), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_600), .B(n_392), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_559), .A2(n_401), .B1(n_403), .B2(n_400), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_567), .A2(n_407), .B(n_404), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_553), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_577), .B(n_409), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_553), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g695 ( .A1(n_525), .A2(n_405), .B1(n_441), .B2(n_392), .Y(n_695) );
INVx5_ASAP7_75t_L g696 ( .A(n_577), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_594), .Y(n_697) );
INVx5_ASAP7_75t_L g698 ( .A(n_577), .Y(n_698) );
BUFx2_ASAP7_75t_L g699 ( .A(n_541), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_581), .Y(n_700) );
BUFx2_ASAP7_75t_L g701 ( .A(n_581), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_531), .B(n_441), .Y(n_702) );
INVxp67_ASAP7_75t_L g703 ( .A(n_537), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_567), .A2(n_421), .B(n_419), .Y(n_704) );
INVx2_ASAP7_75t_SL g705 ( .A(n_538), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_559), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_588), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_589), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_568), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_598), .B(n_445), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_603), .A2(n_592), .B(n_591), .Y(n_711) );
AND2x4_ASAP7_75t_SL g712 ( .A(n_594), .B(n_422), .Y(n_712) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_577), .Y(n_713) );
AOI222xp33_ASAP7_75t_L g714 ( .A1(n_547), .A2(n_429), .B1(n_428), .B2(n_423), .C1(n_430), .C2(n_375), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_593), .A2(n_364), .B(n_336), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_586), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_569), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_596), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_599), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_573), .B(n_376), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_585), .B(n_330), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_569), .B(n_406), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_610), .Y(n_723) );
NAND2x1_ASAP7_75t_L g724 ( .A(n_680), .B(n_575), .Y(n_724) );
OAI21x1_ASAP7_75t_SL g725 ( .A1(n_680), .A2(n_436), .B(n_602), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_666), .B(n_575), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g727 ( .A1(n_711), .A2(n_580), .B(n_579), .Y(n_727) );
AO21x2_ASAP7_75t_L g728 ( .A1(n_715), .A2(n_451), .B(n_444), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_615), .A2(n_451), .B(n_453), .C(n_444), .Y(n_729) );
OAI21x1_ASAP7_75t_L g730 ( .A1(n_659), .A2(n_580), .B(n_579), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_703), .B(n_584), .Y(n_731) );
OAI21x1_ASAP7_75t_L g732 ( .A1(n_686), .A2(n_584), .B(n_453), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_631), .Y(n_733) );
OAI21x1_ASAP7_75t_L g734 ( .A1(n_722), .A2(n_453), .B(n_451), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g735 ( .A1(n_678), .A2(n_459), .B(n_473), .C(n_471), .Y(n_735) );
INVx2_ASAP7_75t_SL g736 ( .A(n_612), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_621), .Y(n_737) );
AO32x2_ASAP7_75t_L g738 ( .A1(n_690), .A2(n_474), .A3(n_475), .B1(n_457), .B2(n_473), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_641), .Y(n_739) );
OAI21xp5_ASAP7_75t_L g740 ( .A1(n_625), .A2(n_459), .B(n_457), .Y(n_740) );
O2A1O1Ixp33_ASAP7_75t_L g741 ( .A1(n_614), .A2(n_457), .B(n_459), .C(n_471), .Y(n_741) );
OAI21x1_ASAP7_75t_SL g742 ( .A1(n_623), .A2(n_473), .B(n_471), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_624), .A2(n_475), .B1(n_474), .B2(n_440), .C(n_408), .Y(n_743) );
O2A1O1Ixp33_ASAP7_75t_L g744 ( .A1(n_617), .A2(n_677), .B(n_674), .C(n_716), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_706), .A2(n_475), .B1(n_331), .B2(n_585), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_646), .B(n_9), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_629), .B(n_9), .Y(n_747) );
OAI21x1_ASAP7_75t_L g748 ( .A1(n_722), .A2(n_585), .B(n_513), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_622), .A2(n_513), .B(n_475), .Y(n_749) );
AOI22x1_ASAP7_75t_L g750 ( .A1(n_627), .A2(n_475), .B1(n_142), .B2(n_143), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_623), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_751) );
OAI21x1_ASAP7_75t_L g752 ( .A1(n_619), .A2(n_82), .B(n_80), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_634), .A2(n_10), .B1(n_12), .B2(n_13), .Y(n_753) );
OAI21xp5_ASAP7_75t_L g754 ( .A1(n_625), .A2(n_14), .B(n_15), .Y(n_754) );
NAND2x1p5_ASAP7_75t_L g755 ( .A(n_607), .B(n_14), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_608), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_642), .Y(n_757) );
BUFx6f_ASAP7_75t_L g758 ( .A(n_618), .Y(n_758) );
CKINVDCx9p33_ASAP7_75t_R g759 ( .A(n_661), .Y(n_759) );
AOI222xp33_ASAP7_75t_L g760 ( .A1(n_700), .A2(n_17), .B1(n_18), .B2(n_21), .C1(n_23), .C2(n_26), .Y(n_760) );
OA21x2_ASAP7_75t_L g761 ( .A1(n_651), .A2(n_670), .B(n_681), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_647), .B(n_17), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_644), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_709), .A2(n_18), .B1(n_21), .B2(n_23), .Y(n_764) );
OAI21x1_ASAP7_75t_L g765 ( .A1(n_619), .A2(n_85), .B(n_84), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_652), .B(n_26), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_616), .Y(n_767) );
AO31x2_ASAP7_75t_L g768 ( .A1(n_645), .A2(n_27), .A3(n_28), .B(n_29), .Y(n_768) );
AOI221xp5_ASAP7_75t_L g769 ( .A1(n_669), .A2(n_27), .B1(n_29), .B2(n_30), .C(n_31), .Y(n_769) );
OAI21x1_ASAP7_75t_L g770 ( .A1(n_628), .A2(n_90), .B(n_86), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_648), .Y(n_771) );
OAI21x1_ASAP7_75t_L g772 ( .A1(n_628), .A2(n_664), .B(n_658), .Y(n_772) );
AOI21x1_ASAP7_75t_L g773 ( .A1(n_710), .A2(n_93), .B(n_92), .Y(n_773) );
OAI21x1_ASAP7_75t_SL g774 ( .A1(n_634), .A2(n_30), .B(n_31), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_675), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_630), .Y(n_776) );
CKINVDCx8_ASAP7_75t_R g777 ( .A(n_635), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_663), .B(n_32), .Y(n_778) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_654), .Y(n_779) );
AOI21xp33_ASAP7_75t_L g780 ( .A1(n_676), .A2(n_690), .B(n_684), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_679), .Y(n_781) );
CKINVDCx6p67_ASAP7_75t_R g782 ( .A(n_663), .Y(n_782) );
O2A1O1Ixp33_ASAP7_75t_SL g783 ( .A1(n_721), .A2(n_161), .B(n_286), .C(n_285), .Y(n_783) );
OAI21x1_ASAP7_75t_L g784 ( .A1(n_692), .A2(n_96), .B(n_94), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_626), .Y(n_785) );
AOI222xp33_ASAP7_75t_L g786 ( .A1(n_701), .A2(n_32), .B1(n_33), .B2(n_34), .C1(n_35), .C2(n_36), .Y(n_786) );
OAI21x1_ASAP7_75t_L g787 ( .A1(n_694), .A2(n_99), .B(n_97), .Y(n_787) );
INVx2_ASAP7_75t_SL g788 ( .A(n_663), .Y(n_788) );
OAI21x1_ASAP7_75t_L g789 ( .A1(n_717), .A2(n_102), .B(n_100), .Y(n_789) );
AO21x2_ASAP7_75t_L g790 ( .A1(n_691), .A2(n_104), .B(n_103), .Y(n_790) );
INVx1_ASAP7_75t_SL g791 ( .A(n_699), .Y(n_791) );
OA21x2_ASAP7_75t_L g792 ( .A1(n_704), .A2(n_109), .B(n_107), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_682), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_682), .Y(n_794) );
OAI21x1_ASAP7_75t_L g795 ( .A1(n_697), .A2(n_609), .B(n_606), .Y(n_795) );
INVx1_ASAP7_75t_SL g796 ( .A(n_654), .Y(n_796) );
AO21x2_ASAP7_75t_L g797 ( .A1(n_673), .A2(n_113), .B(n_111), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_705), .Y(n_798) );
OAI21x1_ASAP7_75t_L g799 ( .A1(n_697), .A2(n_115), .B(n_114), .Y(n_799) );
OAI21x1_ASAP7_75t_L g800 ( .A1(n_639), .A2(n_120), .B(n_118), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_684), .A2(n_35), .B1(n_36), .B2(n_37), .Y(n_801) );
NAND2x1p5_ASAP7_75t_L g802 ( .A(n_607), .B(n_38), .Y(n_802) );
BUFx3_ASAP7_75t_L g803 ( .A(n_688), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_707), .Y(n_804) );
OAI21x1_ASAP7_75t_SL g805 ( .A1(n_633), .A2(n_38), .B(n_39), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_632), .Y(n_806) );
AOI21x1_ASAP7_75t_L g807 ( .A1(n_693), .A2(n_180), .B(n_283), .Y(n_807) );
NAND2x1p5_ASAP7_75t_L g808 ( .A(n_655), .B(n_40), .Y(n_808) );
AND2x4_ASAP7_75t_L g809 ( .A(n_655), .B(n_40), .Y(n_809) );
OAI21x1_ASAP7_75t_L g810 ( .A1(n_672), .A2(n_181), .B(n_282), .Y(n_810) );
OAI21x1_ASAP7_75t_L g811 ( .A1(n_637), .A2(n_178), .B(n_280), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_613), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_685), .Y(n_813) );
OAI21xp5_ASAP7_75t_L g814 ( .A1(n_640), .A2(n_41), .B(n_42), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_643), .B(n_42), .Y(n_815) );
INVx4_ASAP7_75t_L g816 ( .A(n_696), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_695), .B(n_43), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_673), .Y(n_818) );
OAI21x1_ASAP7_75t_L g819 ( .A1(n_687), .A2(n_182), .B(n_274), .Y(n_819) );
OAI21x1_ASAP7_75t_L g820 ( .A1(n_687), .A2(n_176), .B(n_270), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_714), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_821) );
OAI21xp33_ASAP7_75t_L g822 ( .A1(n_702), .A2(n_44), .B(n_45), .Y(n_822) );
OAI21xp5_ASAP7_75t_L g823 ( .A1(n_671), .A2(n_46), .B(n_47), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_693), .Y(n_824) );
O2A1O1Ixp33_ASAP7_75t_SL g825 ( .A1(n_689), .A2(n_186), .B(n_269), .C(n_268), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_605), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_826) );
INVx2_ASAP7_75t_SL g827 ( .A(n_656), .Y(n_827) );
NAND2xp33_ASAP7_75t_R g828 ( .A(n_605), .B(n_48), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_660), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_714), .B(n_50), .Y(n_830) );
OAI21x1_ASAP7_75t_L g831 ( .A1(n_668), .A2(n_187), .B(n_267), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_633), .A2(n_185), .B(n_263), .Y(n_832) );
O2A1O1Ixp33_ASAP7_75t_L g833 ( .A1(n_649), .A2(n_50), .B(n_51), .C(n_52), .Y(n_833) );
AO21x2_ASAP7_75t_L g834 ( .A1(n_719), .A2(n_188), .B(n_260), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_708), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_611), .B(n_51), .Y(n_836) );
INVx3_ASAP7_75t_L g837 ( .A(n_657), .Y(n_837) );
AND2x4_ASAP7_75t_L g838 ( .A(n_657), .B(n_55), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_660), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_660), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_667), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_841) );
OR2x6_ASAP7_75t_L g842 ( .A(n_665), .B(n_57), .Y(n_842) );
AO22x2_ASAP7_75t_L g843 ( .A1(n_653), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_665), .B(n_58), .Y(n_844) );
BUFx2_ASAP7_75t_L g845 ( .A(n_653), .Y(n_845) );
OAI21x1_ASAP7_75t_L g846 ( .A1(n_720), .A2(n_192), .B(n_259), .Y(n_846) );
OAI21x1_ASAP7_75t_L g847 ( .A1(n_618), .A2(n_191), .B(n_258), .Y(n_847) );
AND2x4_ASAP7_75t_L g848 ( .A(n_696), .B(n_59), .Y(n_848) );
AO21x2_ASAP7_75t_L g849 ( .A1(n_683), .A2(n_189), .B(n_257), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_650), .Y(n_850) );
BUFx3_ASAP7_75t_L g851 ( .A(n_662), .Y(n_851) );
OA21x2_ASAP7_75t_L g852 ( .A1(n_718), .A2(n_174), .B(n_256), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_771), .Y(n_853) );
NAND3xp33_ASAP7_75t_L g854 ( .A(n_769), .B(n_618), .C(n_620), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_779), .B(n_712), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g856 ( .A1(n_813), .A2(n_662), .B1(n_638), .B2(n_636), .C(n_620), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_779), .A2(n_662), .B1(n_638), .B2(n_636), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_727), .A2(n_638), .B(n_636), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_723), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_737), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_842), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_842), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_796), .A2(n_620), .B1(n_713), .B2(n_696), .Y(n_863) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_744), .A2(n_713), .B1(n_698), .B2(n_63), .C(n_64), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_744), .B(n_713), .Y(n_865) );
AOI221xp5_ASAP7_75t_L g866 ( .A1(n_766), .A2(n_753), .B1(n_780), .B2(n_815), .C(n_751), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_804), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_828), .A2(n_698), .B1(n_62), .B2(n_63), .Y(n_868) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_778), .A2(n_698), .B1(n_62), .B2(n_65), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_842), .Y(n_870) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_782), .A2(n_61), .B1(n_66), .B2(n_67), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_776), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_808), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_873) );
OA21x2_ASAP7_75t_L g874 ( .A1(n_818), .A2(n_199), .B(n_255), .Y(n_874) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_791), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_780), .A2(n_68), .B1(n_69), .B2(n_71), .Y(n_876) );
OAI221xp5_ASAP7_75t_L g877 ( .A1(n_766), .A2(n_72), .B1(n_73), .B2(n_75), .C(n_125), .Y(n_877) );
BUFx6f_ASAP7_75t_L g878 ( .A(n_758), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_762), .Y(n_879) );
OAI211xp5_ASAP7_75t_SL g880 ( .A1(n_760), .A2(n_72), .B(n_73), .C(n_131), .Y(n_880) );
AO21x1_ASAP7_75t_L g881 ( .A1(n_751), .A2(n_132), .B(n_135), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_830), .A2(n_136), .B1(n_137), .B2(n_140), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_843), .A2(n_144), .B1(n_145), .B2(n_146), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_727), .A2(n_147), .B(n_148), .Y(n_884) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_758), .Y(n_885) );
OAI22xp33_ASAP7_75t_SL g886 ( .A1(n_753), .A2(n_149), .B1(n_151), .B2(n_153), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_762), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_736), .B(n_747), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g889 ( .A1(n_843), .A2(n_157), .B1(n_159), .B2(n_162), .Y(n_889) );
BUFx4f_ASAP7_75t_L g890 ( .A(n_808), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_843), .A2(n_163), .B1(n_164), .B2(n_170), .Y(n_891) );
INVx4_ASAP7_75t_L g892 ( .A(n_816), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_815), .A2(n_173), .B1(n_193), .B2(n_195), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_726), .A2(n_200), .B(n_202), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_755), .A2(n_203), .B1(n_205), .B2(n_206), .Y(n_895) );
AOI222xp33_ASAP7_75t_L g896 ( .A1(n_845), .A2(n_208), .B1(n_210), .B2(n_211), .C1(n_212), .C2(n_215), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_755), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_802), .Y(n_898) );
A2O1A1Ixp33_ASAP7_75t_L g899 ( .A1(n_833), .A2(n_216), .B(n_217), .C(n_219), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_731), .B(n_291), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_731), .B(n_220), .Y(n_901) );
CKINVDCx6p67_ASAP7_75t_R g902 ( .A(n_767), .Y(n_902) );
AO21x2_ASAP7_75t_L g903 ( .A1(n_735), .A2(n_221), .B(n_222), .Y(n_903) );
OAI211xp5_ASAP7_75t_SL g904 ( .A1(n_786), .A2(n_223), .B(n_224), .C(n_225), .Y(n_904) );
AOI21xp5_ASAP7_75t_L g905 ( .A1(n_726), .A2(n_226), .B(n_227), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_802), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_821), .B(n_231), .Y(n_907) );
AOI21xp5_ASAP7_75t_L g908 ( .A1(n_730), .A2(n_234), .B(n_235), .Y(n_908) );
INVx4_ASAP7_75t_L g909 ( .A(n_816), .Y(n_909) );
AOI222xp33_ASAP7_75t_L g910 ( .A1(n_788), .A2(n_236), .B1(n_237), .B2(n_245), .C1(n_247), .C2(n_249), .Y(n_910) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_817), .A2(n_251), .B1(n_253), .B2(n_774), .Y(n_911) );
OR2x6_ASAP7_75t_L g912 ( .A(n_809), .B(n_838), .Y(n_912) );
INVx3_ASAP7_75t_L g913 ( .A(n_851), .Y(n_913) );
OAI22x1_ASAP7_75t_L g914 ( .A1(n_841), .A2(n_850), .B1(n_809), .B2(n_848), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_821), .A2(n_826), .B1(n_801), .B2(n_823), .Y(n_915) );
AOI221xp5_ASAP7_75t_L g916 ( .A1(n_833), .A2(n_769), .B1(n_743), .B2(n_739), .C(n_757), .Y(n_916) );
AND2x4_ASAP7_75t_L g917 ( .A(n_837), .B(n_793), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_763), .Y(n_918) );
OAI22xp33_ASAP7_75t_L g919 ( .A1(n_828), .A2(n_777), .B1(n_767), .B2(n_836), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_801), .Y(n_920) );
OAI22xp33_ASAP7_75t_L g921 ( .A1(n_836), .A2(n_826), .B1(n_823), .B2(n_798), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_835), .B(n_812), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_775), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_746), .A2(n_838), .B1(n_794), .B2(n_743), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_764), .B(n_781), .Y(n_925) );
BUFx4f_ASAP7_75t_SL g926 ( .A(n_803), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_844), .Y(n_927) );
INVx4_ASAP7_75t_L g928 ( .A(n_756), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_746), .A2(n_844), .B1(n_824), .B2(n_761), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_764), .B(n_848), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_761), .A2(n_742), .B1(n_822), .B2(n_754), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_785), .B(n_806), .Y(n_932) );
OA21x2_ASAP7_75t_L g933 ( .A1(n_772), .A2(n_734), .B(n_832), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_768), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_814), .A2(n_754), .B1(n_852), .B2(n_729), .Y(n_935) );
AOI21xp33_ASAP7_75t_L g936 ( .A1(n_741), .A2(n_814), .B(n_805), .Y(n_936) );
AO21x2_ASAP7_75t_L g937 ( .A1(n_735), .A2(n_797), .B(n_773), .Y(n_937) );
HB1xp67_ASAP7_75t_L g938 ( .A(n_829), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g939 ( .A1(n_740), .A2(n_749), .B(n_795), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g940 ( .A1(n_827), .A2(n_729), .B1(n_741), .B2(n_740), .C(n_745), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_837), .A2(n_725), .B1(n_852), .B2(n_840), .Y(n_941) );
AOI211xp5_ASAP7_75t_L g942 ( .A1(n_825), .A2(n_783), .B(n_831), .C(n_759), .Y(n_942) );
OAI22xp5_ASAP7_75t_SL g943 ( .A1(n_733), .A2(n_759), .B1(n_724), .B2(n_792), .Y(n_943) );
AOI221xp5_ASAP7_75t_L g944 ( .A1(n_825), .A2(n_745), .B1(n_783), .B2(n_728), .C(n_839), .Y(n_944) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_834), .A2(n_849), .B1(n_770), .B2(n_765), .Y(n_945) );
AOI21xp5_ASAP7_75t_L g946 ( .A1(n_792), .A2(n_748), .B(n_797), .Y(n_946) );
INVxp33_ASAP7_75t_L g947 ( .A(n_758), .Y(n_947) );
BUFx3_ASAP7_75t_L g948 ( .A(n_758), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_750), .A2(n_807), .B1(n_768), .B2(n_738), .Y(n_949) );
AND2x4_ASAP7_75t_L g950 ( .A(n_810), .B(n_846), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_768), .B(n_738), .Y(n_951) );
AOI21xp5_ASAP7_75t_L g952 ( .A1(n_834), .A2(n_790), .B(n_732), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_768), .B(n_849), .Y(n_953) );
OR2x6_ASAP7_75t_L g954 ( .A(n_752), .B(n_820), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_738), .B(n_790), .Y(n_955) );
OAI21x1_ASAP7_75t_L g956 ( .A1(n_784), .A2(n_787), .B(n_789), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_800), .B(n_819), .Y(n_957) );
AOI21xp5_ASAP7_75t_L g958 ( .A1(n_811), .A2(n_799), .B(n_847), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_779), .A2(n_525), .B1(n_581), .B2(n_796), .Y(n_959) );
AOI222xp33_ASAP7_75t_L g960 ( .A1(n_830), .A2(n_468), .B1(n_779), .B2(n_796), .C1(n_688), .C2(n_442), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_830), .B(n_512), .Y(n_961) );
AOI221xp5_ASAP7_75t_L g962 ( .A1(n_744), .A2(n_547), .B1(n_586), .B2(n_624), .C(n_716), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_830), .B(n_512), .Y(n_963) );
OAI211xp5_ASAP7_75t_L g964 ( .A1(n_821), .A2(n_786), .B(n_760), .C(n_714), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_779), .B(n_716), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_723), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_779), .A2(n_796), .B1(n_842), .B2(n_623), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_744), .A2(n_547), .B1(n_586), .B2(n_624), .C(n_716), .Y(n_968) );
NOR2x1_ASAP7_75t_SL g969 ( .A(n_842), .B(n_680), .Y(n_969) );
OAI221xp5_ASAP7_75t_L g970 ( .A1(n_813), .A2(n_703), .B1(n_586), .B2(n_601), .C(n_583), .Y(n_970) );
OA21x2_ASAP7_75t_L g971 ( .A1(n_953), .A2(n_952), .B(n_946), .Y(n_971) );
INVxp67_ASAP7_75t_SL g972 ( .A(n_890), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g973 ( .A1(n_959), .A2(n_964), .B1(n_970), .B2(n_968), .C(n_962), .Y(n_973) );
BUFx2_ASAP7_75t_L g974 ( .A(n_912), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_934), .Y(n_975) );
OR2x2_ASAP7_75t_L g976 ( .A(n_912), .B(n_920), .Y(n_976) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_961), .B(n_963), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_912), .B(n_853), .Y(n_978) );
OR2x2_ASAP7_75t_L g979 ( .A(n_965), .B(n_967), .Y(n_979) );
BUFx3_ASAP7_75t_L g980 ( .A(n_926), .Y(n_980) );
AOI21xp5_ASAP7_75t_SL g981 ( .A1(n_895), .A2(n_915), .B(n_969), .Y(n_981) );
OAI21xp5_ASAP7_75t_L g982 ( .A1(n_854), .A2(n_916), .B(n_866), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_865), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_878), .Y(n_984) );
OR2x2_ASAP7_75t_L g985 ( .A(n_967), .B(n_927), .Y(n_985) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_875), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_915), .B(n_879), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_878), .Y(n_988) );
INVx2_ASAP7_75t_L g989 ( .A(n_885), .Y(n_989) );
OR2x2_ASAP7_75t_L g990 ( .A(n_887), .B(n_855), .Y(n_990) );
BUFx3_ASAP7_75t_L g991 ( .A(n_892), .Y(n_991) );
BUFx3_ASAP7_75t_L g992 ( .A(n_892), .Y(n_992) );
CKINVDCx8_ASAP7_75t_R g993 ( .A(n_902), .Y(n_993) );
OR2x2_ASAP7_75t_L g994 ( .A(n_867), .B(n_859), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_880), .A2(n_960), .B1(n_919), .B2(n_914), .Y(n_995) );
AND2x4_ASAP7_75t_L g996 ( .A(n_897), .B(n_898), .Y(n_996) );
OAI31xp33_ASAP7_75t_L g997 ( .A1(n_871), .A2(n_904), .A3(n_873), .B(n_921), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_960), .B(n_860), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_923), .B(n_872), .Y(n_999) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_890), .Y(n_1000) );
INVxp67_ASAP7_75t_L g1001 ( .A(n_888), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_966), .B(n_925), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_930), .B(n_951), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_865), .Y(n_1004) );
INVxp67_ASAP7_75t_L g1005 ( .A(n_922), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_918), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_933), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_906), .B(n_932), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_954), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_929), .B(n_873), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_907), .B(n_924), .Y(n_1011) );
INVxp67_ASAP7_75t_L g1012 ( .A(n_861), .Y(n_1012) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_909), .B(n_870), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_874), .Y(n_1014) );
OAI221xp5_ASAP7_75t_SL g1015 ( .A1(n_868), .A2(n_877), .B1(n_876), .B2(n_864), .C(n_869), .Y(n_1015) );
OR2x2_ASAP7_75t_L g1016 ( .A(n_862), .B(n_909), .Y(n_1016) );
OA21x2_ASAP7_75t_L g1017 ( .A1(n_939), .A2(n_949), .B(n_957), .Y(n_1017) );
BUFx2_ASAP7_75t_L g1018 ( .A(n_948), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_917), .B(n_938), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_896), .B(n_917), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_896), .B(n_913), .Y(n_1021) );
INVxp67_ASAP7_75t_R g1022 ( .A(n_943), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_954), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_913), .B(n_910), .Y(n_1024) );
OA21x2_ASAP7_75t_L g1025 ( .A1(n_949), .A2(n_956), .B(n_958), .Y(n_1025) );
BUFx3_ASAP7_75t_L g1026 ( .A(n_856), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_895), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_955), .Y(n_1028) );
INVxp67_ASAP7_75t_L g1029 ( .A(n_910), .Y(n_1029) );
AO22x1_ASAP7_75t_L g1030 ( .A1(n_935), .A2(n_947), .B1(n_950), .B2(n_928), .Y(n_1030) );
AND2x4_ASAP7_75t_L g1031 ( .A(n_950), .B(n_903), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_854), .B(n_935), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_903), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_931), .B(n_857), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_883), .B(n_891), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_889), .B(n_911), .Y(n_1036) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_863), .B(n_884), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_881), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_940), .A2(n_936), .B1(n_882), .B2(n_886), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_937), .Y(n_1040) );
INVx5_ASAP7_75t_L g1041 ( .A(n_928), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_899), .B(n_936), .Y(n_1042) );
BUFx8_ASAP7_75t_SL g1043 ( .A(n_900), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_937), .Y(n_1044) );
AND2x4_ASAP7_75t_L g1045 ( .A(n_858), .B(n_908), .Y(n_1045) );
INVx2_ASAP7_75t_L g1046 ( .A(n_901), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_893), .B(n_941), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_942), .B(n_945), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_942), .B(n_944), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_894), .B(n_905), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_912), .B(n_853), .Y(n_1051) );
INVx1_ASAP7_75t_SL g1052 ( .A(n_902), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_912), .B(n_853), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_912), .B(n_920), .Y(n_1054) );
OR2x6_ASAP7_75t_L g1055 ( .A(n_912), .B(n_842), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_912), .B(n_853), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_934), .Y(n_1057) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_912), .B(n_920), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_934), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_912), .B(n_853), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_934), .Y(n_1061) );
INVxp67_ASAP7_75t_SL g1062 ( .A(n_1027), .Y(n_1062) );
BUFx2_ASAP7_75t_L g1063 ( .A(n_1055), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_998), .B(n_1002), .Y(n_1064) );
AND2x4_ASAP7_75t_SL g1065 ( .A(n_1055), .B(n_1020), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_1020), .A2(n_1029), .B1(n_1021), .B2(n_995), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_1021), .A2(n_973), .B1(n_1024), .B2(n_1011), .Y(n_1067) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_1055), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1003), .B(n_1002), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_975), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_975), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_1003), .B(n_985), .Y(n_1072) );
A2O1A1Ixp33_ASAP7_75t_SL g1073 ( .A1(n_977), .A2(n_1038), .B(n_1012), .C(n_982), .Y(n_1073) );
OAI211xp5_ASAP7_75t_L g1074 ( .A1(n_981), .A2(n_993), .B(n_997), .C(n_1000), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1057), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1028), .B(n_987), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1057), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1059), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1028), .B(n_987), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1059), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_983), .B(n_1004), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_983), .B(n_1004), .Y(n_1082) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_1055), .Y(n_1083) );
NAND3xp33_ASAP7_75t_L g1084 ( .A(n_1038), .B(n_1039), .C(n_981), .Y(n_1084) );
INVx4_ASAP7_75t_L g1085 ( .A(n_991), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_999), .B(n_1061), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1061), .Y(n_1087) );
NOR2x1_ASAP7_75t_SL g1088 ( .A(n_991), .B(n_992), .Y(n_1088) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_1024), .A2(n_1015), .B1(n_1041), .B2(n_1000), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_999), .B(n_1008), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1008), .B(n_1010), .Y(n_1091) );
OR2x2_ASAP7_75t_L g1092 ( .A(n_985), .B(n_979), .Y(n_1092) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_1005), .A2(n_1001), .B1(n_1010), .B2(n_986), .C(n_1011), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_990), .B(n_1006), .Y(n_1094) );
NOR2xp33_ASAP7_75t_L g1095 ( .A(n_1052), .B(n_972), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_979), .B(n_1058), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_976), .B(n_1058), .Y(n_1097) );
OAI221xp5_ASAP7_75t_L g1098 ( .A1(n_990), .A2(n_976), .B1(n_1054), .B2(n_993), .C(n_1016), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1009), .Y(n_1099) );
INVxp67_ASAP7_75t_SL g1100 ( .A(n_992), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1006), .B(n_1023), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_1054), .B(n_994), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1009), .B(n_1023), .Y(n_1103) );
NOR2xp33_ASAP7_75t_L g1104 ( .A(n_980), .B(n_1041), .Y(n_1104) );
INVx2_ASAP7_75t_SL g1105 ( .A(n_1041), .Y(n_1105) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_1036), .A2(n_1035), .B1(n_1049), .B2(n_996), .C(n_974), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1049), .B(n_994), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_978), .B(n_1060), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_978), .B(n_1060), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1032), .B(n_1056), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1032), .B(n_1056), .Y(n_1111) );
INVx3_ASAP7_75t_L g1112 ( .A(n_1031), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1051), .B(n_1053), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1048), .B(n_1022), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_1036), .A2(n_1035), .B1(n_974), .B2(n_1043), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1022), .B(n_1042), .Y(n_1116) );
INVxp67_ASAP7_75t_L g1117 ( .A(n_1019), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1007), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1042), .B(n_996), .Y(n_1119) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_1018), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_996), .B(n_1044), .Y(n_1121) );
INVx2_ASAP7_75t_SL g1122 ( .A(n_1041), .Y(n_1122) );
OR2x2_ASAP7_75t_L g1123 ( .A(n_1016), .B(n_1018), .Y(n_1123) );
NOR2xp33_ASAP7_75t_L g1124 ( .A(n_980), .B(n_1041), .Y(n_1124) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_1034), .B(n_1013), .Y(n_1125) );
AND2x4_ASAP7_75t_L g1126 ( .A(n_1112), .B(n_1031), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1086), .Y(n_1127) );
BUFx2_ASAP7_75t_L g1128 ( .A(n_1085), .Y(n_1128) );
NAND3xp33_ASAP7_75t_SL g1129 ( .A(n_1074), .B(n_1041), .C(n_1047), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1069), .B(n_1013), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1069), .B(n_1013), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1110), .B(n_1031), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1110), .B(n_1040), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1086), .Y(n_1134) );
NOR2xp33_ASAP7_75t_L g1135 ( .A(n_1114), .B(n_1026), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1090), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1090), .Y(n_1137) );
NOR2xp33_ASAP7_75t_L g1138 ( .A(n_1114), .B(n_1026), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1107), .B(n_1046), .Y(n_1139) );
NOR2xp33_ASAP7_75t_L g1140 ( .A(n_1116), .B(n_1064), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1070), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1111), .B(n_1040), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1070), .Y(n_1143) );
AND2x4_ASAP7_75t_L g1144 ( .A(n_1112), .B(n_1045), .Y(n_1144) );
INVxp67_ASAP7_75t_SL g1145 ( .A(n_1088), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1111), .B(n_1033), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1076), .B(n_1033), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1076), .B(n_971), .Y(n_1148) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_1072), .B(n_1034), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1150 ( .A(n_1112), .B(n_1045), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1079), .B(n_971), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1079), .B(n_971), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1107), .B(n_1046), .Y(n_1153) );
INVx1_ASAP7_75t_SL g1154 ( .A(n_1085), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1091), .B(n_971), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1091), .B(n_1017), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1072), .B(n_1030), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1094), .B(n_1030), .Y(n_1158) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1118), .Y(n_1159) );
NOR2x1_ASAP7_75t_L g1160 ( .A(n_1085), .B(n_984), .Y(n_1160) );
INVx2_ASAP7_75t_SL g1161 ( .A(n_1085), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1071), .Y(n_1162) );
OR2x2_ASAP7_75t_L g1163 ( .A(n_1092), .B(n_1017), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1101), .B(n_1017), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_1102), .B(n_1123), .Y(n_1165) );
INVx1_ASAP7_75t_SL g1166 ( .A(n_1123), .Y(n_1166) );
OR2x2_ASAP7_75t_L g1167 ( .A(n_1108), .B(n_988), .Y(n_1167) );
NAND4xp25_ASAP7_75t_L g1168 ( .A(n_1106), .B(n_1050), .C(n_1037), .D(n_1045), .Y(n_1168) );
NAND4xp25_ASAP7_75t_L g1169 ( .A(n_1066), .B(n_1050), .C(n_1037), .D(n_1045), .Y(n_1169) );
NOR2xp67_ASAP7_75t_L g1170 ( .A(n_1105), .B(n_1014), .Y(n_1170) );
INVx3_ASAP7_75t_L g1171 ( .A(n_1105), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1109), .B(n_989), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1071), .Y(n_1173) );
OR2x2_ASAP7_75t_SL g1174 ( .A(n_1084), .B(n_1017), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1075), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1092), .B(n_1025), .Y(n_1176) );
INVx2_ASAP7_75t_SL g1177 ( .A(n_1122), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1075), .Y(n_1178) );
NOR2xp33_ASAP7_75t_L g1179 ( .A(n_1116), .B(n_1037), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1077), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1101), .B(n_1025), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1141), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1143), .Y(n_1183) );
INVx2_ASAP7_75t_SL g1184 ( .A(n_1128), .Y(n_1184) );
NOR2xp33_ASAP7_75t_L g1185 ( .A(n_1140), .B(n_1135), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1155), .B(n_1119), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_1149), .B(n_1096), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1136), .B(n_1093), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1155), .B(n_1119), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1162), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1173), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1175), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1137), .B(n_1067), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1127), .B(n_1134), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1178), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1180), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1156), .B(n_1103), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1165), .B(n_1096), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1140), .B(n_1117), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1139), .B(n_1082), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1166), .Y(n_1201) );
INVx2_ASAP7_75t_SL g1202 ( .A(n_1161), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1153), .B(n_1082), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_1147), .B(n_1081), .Y(n_1204) );
OR2x2_ASAP7_75t_L g1205 ( .A(n_1163), .B(n_1097), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1147), .B(n_1081), .Y(n_1206) );
OR2x2_ASAP7_75t_L g1207 ( .A(n_1130), .B(n_1125), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1156), .B(n_1103), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1148), .B(n_1078), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1148), .B(n_1121), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1151), .B(n_1078), .Y(n_1211) );
OAI31xp33_ASAP7_75t_L g1212 ( .A1(n_1154), .A2(n_1065), .A3(n_1089), .B(n_1073), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1151), .B(n_1121), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1152), .B(n_1099), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1215 ( .A(n_1163), .B(n_1097), .Y(n_1215) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1159), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1131), .Y(n_1217) );
BUFx2_ASAP7_75t_L g1218 ( .A(n_1145), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1152), .B(n_1080), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1167), .Y(n_1220) );
AOI22xp5_ASAP7_75t_L g1221 ( .A1(n_1135), .A2(n_1065), .B1(n_1115), .B2(n_1098), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1146), .B(n_1077), .Y(n_1222) );
AOI221xp5_ASAP7_75t_L g1223 ( .A1(n_1169), .A2(n_1084), .B1(n_1099), .B2(n_1062), .C(n_1087), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1172), .Y(n_1224) );
AND2x2_ASAP7_75t_SL g1225 ( .A(n_1157), .B(n_1083), .Y(n_1225) );
INVx2_ASAP7_75t_L g1226 ( .A(n_1159), .Y(n_1226) );
OR2x6_ASAP7_75t_L g1227 ( .A(n_1161), .B(n_1063), .Y(n_1227) );
OAI21xp33_ASAP7_75t_L g1228 ( .A1(n_1185), .A2(n_1168), .B(n_1179), .Y(n_1228) );
INVxp67_ASAP7_75t_L g1229 ( .A(n_1202), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_1221), .A2(n_1100), .B1(n_1138), .B2(n_1179), .Y(n_1230) );
AOI222xp33_ASAP7_75t_L g1231 ( .A1(n_1188), .A2(n_1138), .B1(n_1158), .B2(n_1164), .C1(n_1181), .C2(n_1146), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1198), .Y(n_1232) );
OAI22xp33_ASAP7_75t_L g1233 ( .A1(n_1218), .A2(n_1157), .B1(n_1083), .B2(n_1063), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1198), .Y(n_1234) );
NOR2xp33_ASAP7_75t_L g1235 ( .A(n_1185), .B(n_1129), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1205), .Y(n_1236) );
NOR3xp33_ASAP7_75t_L g1237 ( .A(n_1223), .B(n_1095), .C(n_1124), .Y(n_1237) );
OAI31xp33_ASAP7_75t_L g1238 ( .A1(n_1212), .A2(n_1104), .A3(n_1068), .B(n_1177), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1205), .Y(n_1239) );
AOI211xp5_ASAP7_75t_L g1240 ( .A1(n_1202), .A2(n_1176), .B(n_1068), .C(n_1125), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1187), .B(n_1133), .Y(n_1241) );
INVxp67_ASAP7_75t_L g1242 ( .A(n_1184), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1215), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1186), .B(n_1164), .Y(n_1244) );
INVx4_ASAP7_75t_L g1245 ( .A(n_1227), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1214), .B(n_1181), .Y(n_1246) );
AOI221xp5_ASAP7_75t_L g1247 ( .A1(n_1193), .A2(n_1132), .B1(n_1087), .B2(n_1080), .C(n_1133), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1186), .B(n_1132), .Y(n_1248) );
OR2x2_ASAP7_75t_L g1249 ( .A(n_1187), .B(n_1142), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1214), .B(n_1217), .Y(n_1250) );
AND2x4_ASAP7_75t_L g1251 ( .A(n_1184), .B(n_1144), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1215), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1182), .Y(n_1253) );
NOR2xp33_ASAP7_75t_L g1254 ( .A(n_1201), .B(n_1177), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1189), .B(n_1142), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1220), .B(n_1176), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1189), .B(n_1144), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1197), .B(n_1126), .Y(n_1258) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1253), .Y(n_1259) );
AND3x1_ASAP7_75t_L g1260 ( .A(n_1238), .B(n_1199), .C(n_1122), .Y(n_1260) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1241), .Y(n_1261) );
INVx2_ASAP7_75t_L g1262 ( .A(n_1249), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1244), .B(n_1197), .Y(n_1263) );
NOR2xp67_ASAP7_75t_L g1264 ( .A(n_1245), .B(n_1171), .Y(n_1264) );
NAND2xp5_ASAP7_75t_SL g1265 ( .A(n_1245), .B(n_1225), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1256), .Y(n_1266) );
XNOR2xp5_ASAP7_75t_L g1267 ( .A(n_1230), .B(n_1224), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1236), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1239), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1244), .B(n_1208), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1231), .B(n_1208), .Y(n_1271) );
AOI211xp5_ASAP7_75t_L g1272 ( .A1(n_1235), .A2(n_1170), .B(n_1171), .C(n_1120), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1243), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1252), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1232), .Y(n_1275) );
NAND2xp5_ASAP7_75t_SL g1276 ( .A(n_1245), .B(n_1225), .Y(n_1276) );
OAI321xp33_ASAP7_75t_L g1277 ( .A1(n_1235), .A2(n_1227), .A3(n_1211), .B1(n_1209), .B2(n_1219), .C(n_1222), .Y(n_1277) );
INVx1_ASAP7_75t_SL g1278 ( .A(n_1255), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1263), .B(n_1257), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_1271), .A2(n_1228), .B1(n_1237), .B2(n_1267), .Y(n_1280) );
OAI31xp33_ASAP7_75t_SL g1281 ( .A1(n_1267), .A2(n_1233), .A3(n_1247), .B(n_1254), .Y(n_1281) );
NAND2xp5_ASAP7_75t_SL g1282 ( .A(n_1260), .B(n_1233), .Y(n_1282) );
O2A1O1Ixp33_ASAP7_75t_L g1283 ( .A1(n_1277), .A2(n_1242), .B(n_1229), .C(n_1254), .Y(n_1283) );
NAND2xp33_ASAP7_75t_L g1284 ( .A(n_1265), .B(n_1171), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1259), .Y(n_1285) );
AOI22x1_ASAP7_75t_L g1286 ( .A1(n_1278), .A2(n_1251), .B1(n_1088), .B2(n_1257), .Y(n_1286) );
OAI21xp5_ASAP7_75t_L g1287 ( .A1(n_1272), .A2(n_1240), .B(n_1258), .Y(n_1287) );
NAND4xp25_ASAP7_75t_SL g1288 ( .A(n_1272), .B(n_1234), .C(n_1255), .D(n_1248), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1259), .Y(n_1289) );
XNOR2x1_ASAP7_75t_L g1290 ( .A(n_1263), .B(n_1251), .Y(n_1290) );
OAI21xp5_ASAP7_75t_L g1291 ( .A1(n_1276), .A2(n_1251), .B(n_1227), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1268), .Y(n_1292) );
NAND3xp33_ASAP7_75t_SL g1293 ( .A(n_1282), .B(n_1270), .C(n_1262), .Y(n_1293) );
AOI221xp5_ASAP7_75t_L g1294 ( .A1(n_1280), .A2(n_1266), .B1(n_1275), .B2(n_1273), .C(n_1274), .Y(n_1294) );
OAI221xp5_ASAP7_75t_SL g1295 ( .A1(n_1281), .A2(n_1266), .B1(n_1227), .B2(n_1262), .C(n_1261), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1292), .Y(n_1296) );
NAND4xp75_ASAP7_75t_L g1297 ( .A(n_1291), .B(n_1264), .C(n_1275), .D(n_1274), .Y(n_1297) );
OAI21xp5_ASAP7_75t_L g1298 ( .A1(n_1288), .A2(n_1264), .B(n_1270), .Y(n_1298) );
AOI221xp5_ASAP7_75t_L g1299 ( .A1(n_1283), .A2(n_1273), .B1(n_1269), .B2(n_1268), .C(n_1261), .Y(n_1299) );
AOI211xp5_ASAP7_75t_L g1300 ( .A1(n_1284), .A2(n_1269), .B(n_1250), .C(n_1150), .Y(n_1300) );
AOI221xp5_ASAP7_75t_L g1301 ( .A1(n_1287), .A2(n_1194), .B1(n_1246), .B2(n_1196), .C(n_1195), .Y(n_1301) );
HB1xp67_ASAP7_75t_L g1302 ( .A(n_1296), .Y(n_1302) );
NOR2xp33_ASAP7_75t_L g1303 ( .A(n_1295), .B(n_1290), .Y(n_1303) );
NAND2xp5_ASAP7_75t_SL g1304 ( .A(n_1298), .B(n_1286), .Y(n_1304) );
OAI321xp33_ASAP7_75t_L g1305 ( .A1(n_1293), .A2(n_1292), .A3(n_1279), .B1(n_1284), .B2(n_1285), .C(n_1289), .Y(n_1305) );
AND2x4_ASAP7_75t_L g1306 ( .A(n_1297), .B(n_1279), .Y(n_1306) );
AOI21xp5_ASAP7_75t_L g1307 ( .A1(n_1299), .A2(n_1286), .B(n_1290), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1302), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1303), .B(n_1294), .Y(n_1309) );
OAI22xp33_ASAP7_75t_L g1310 ( .A1(n_1305), .A2(n_1301), .B1(n_1300), .B2(n_1207), .Y(n_1310) );
AND2x4_ASAP7_75t_SL g1311 ( .A(n_1306), .B(n_1113), .Y(n_1311) );
OR4x2_ASAP7_75t_L g1312 ( .A(n_1304), .B(n_1174), .C(n_1204), .D(n_1206), .Y(n_1312) );
HB1xp67_ASAP7_75t_L g1313 ( .A(n_1308), .Y(n_1313) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1311), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1309), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1310), .Y(n_1316) );
OAI221xp5_ASAP7_75t_L g1317 ( .A1(n_1316), .A2(n_1307), .B1(n_1312), .B2(n_1160), .C(n_1192), .Y(n_1317) );
OAI22xp5_ASAP7_75t_L g1318 ( .A1(n_1315), .A2(n_1190), .B1(n_1191), .B2(n_1183), .Y(n_1318) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_1317), .A2(n_1314), .B1(n_1313), .B2(n_1203), .Y(n_1319) );
AO22x2_ASAP7_75t_L g1320 ( .A1(n_1318), .A2(n_1200), .B1(n_1226), .B2(n_1216), .Y(n_1320) );
UNKNOWN g1321 ( );
AOI22xp5_ASAP7_75t_SL g1322 ( .A1(n_1321), .A2(n_1320), .B1(n_1150), .B2(n_1144), .Y(n_1322) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_1322), .A2(n_1150), .B1(n_1126), .B2(n_1213), .C(n_1210), .Y(n_1323) );
endmodule