module fake_jpeg_28990_n_61 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_61);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_61;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVxp67_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_2),
.B(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NAND2x1_ASAP7_75t_SL g23 ( 
.A(n_8),
.B(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_7),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_25),
.B(n_23),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

AND2x6_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_9),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_10),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_40),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_51),
.C(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_40),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_11),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_56),
.B(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);


endmodule