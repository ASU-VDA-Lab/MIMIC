module fake_jpeg_10632_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx4f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_20),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_7),
.Y(n_20)
);

HAxp5_ASAP7_75t_SL g21 ( 
.A(n_11),
.B(n_7),
.CON(n_21),
.SN(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_35),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_19),
.B1(n_13),
.B2(n_16),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_18),
.B1(n_26),
.B2(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

AO22x2_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_31),
.B1(n_33),
.B2(n_26),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_44),
.B1(n_12),
.B2(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_25),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

OAI32xp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_9),
.A3(n_10),
.B1(n_29),
.B2(n_24),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_12),
.B(n_24),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_47),
.B(n_51),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_51),
.B1(n_41),
.B2(n_44),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_24),
.B(n_9),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_24),
.C(n_27),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_41),
.C(n_38),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_10),
.B1(n_9),
.B2(n_27),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_10),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_56),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_0),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_59),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_65),
.B(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_59),
.Y(n_65)
);

NOR3xp33_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_53),
.C(n_57),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_65),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_64),
.B(n_62),
.C(n_61),
.Y(n_73)
);

INVxp33_ASAP7_75t_SL g71 ( 
.A(n_68),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_67),
.C(n_5),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_72),
.B(n_5),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_7),
.B1(n_4),
.B2(n_6),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_76),
.B(n_6),
.Y(n_79)
);


endmodule