module fake_jpeg_12771_n_92 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_92);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_92;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_27),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_48),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_36),
.B(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_56),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_38),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_7),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_26),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_72),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_13),
.C(n_23),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_65),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_1),
.B(n_2),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_1),
.B(n_3),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_4),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_70),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_16),
.B(n_22),
.C(n_20),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_12),
.C(n_19),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_4),
.B(n_6),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_73),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_64),
.B1(n_67),
.B2(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_80),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_84),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_79),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_78),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_85),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_85),
.C(n_86),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_76),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_76),
.B(n_77),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_90),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_78),
.Y(n_92)
);


endmodule