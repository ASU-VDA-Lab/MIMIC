module fake_jpeg_19851_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_0),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_1),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_48),
.B1(n_49),
.B2(n_46),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_66),
.B1(n_2),
.B2(n_3),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_46),
.B1(n_52),
.B2(n_51),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_41),
.B1(n_4),
.B2(n_5),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_53),
.B1(n_50),
.B2(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_69),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_40),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_2),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_79),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_77),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_85),
.B1(n_72),
.B2(n_4),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_23),
.B(n_37),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_12),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_3),
.B1(n_6),
.B2(n_11),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_85),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_90),
.B(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_97),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_79),
.C(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_6),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_101),
.B1(n_86),
.B2(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_105),
.B(n_106),
.Y(n_107)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_89),
.B1(n_94),
.B2(n_100),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_102),
.B(n_18),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_93),
.C(n_20),
.Y(n_110)
);

AOI211xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_16),
.B(n_27),
.C(n_29),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_30),
.B(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_32),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_33),
.Y(n_114)
);


endmodule