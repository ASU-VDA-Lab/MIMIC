module real_aes_16117_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1600;
wire n_805;
wire n_619;
wire n_1250;
wire n_1284;
wire n_1583;
wire n_360;
wire n_1095;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_1584;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_0), .A2(n_53), .B1(n_453), .B2(n_782), .Y(n_781) );
INVxp67_ASAP7_75t_SL g810 ( .A(n_0), .Y(n_810) );
INVx1_ASAP7_75t_L g322 ( .A(n_1), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_1), .B(n_332), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_2), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_3), .A2(n_230), .B1(n_1143), .B2(n_1278), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1294 ( .A1(n_3), .A2(n_175), .B1(n_1105), .B2(n_1221), .Y(n_1294) );
INVx1_ASAP7_75t_L g611 ( .A(n_4), .Y(n_611) );
INVx1_ASAP7_75t_L g962 ( .A(n_5), .Y(n_962) );
OAI22xp5_ASAP7_75t_SL g976 ( .A1(n_6), .A2(n_199), .B1(n_466), .B2(n_533), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_6), .A2(n_199), .B1(n_980), .B2(n_981), .Y(n_979) );
OAI22xp33_ASAP7_75t_SL g872 ( .A1(n_7), .A2(n_302), .B1(n_791), .B2(n_873), .Y(n_872) );
OAI22xp33_ASAP7_75t_L g887 ( .A1(n_7), .A2(n_163), .B1(n_477), .B2(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g1072 ( .A(n_8), .Y(n_1072) );
INVx1_ASAP7_75t_L g949 ( .A(n_9), .Y(n_949) );
INVx1_ASAP7_75t_L g1270 ( .A(n_10), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g1299 ( .A1(n_10), .A2(n_230), .B1(n_1089), .B2(n_1221), .Y(n_1299) );
AOI22xp5_ASAP7_75t_L g1336 ( .A1(n_11), .A2(n_52), .B1(n_1311), .B2(n_1317), .Y(n_1336) );
CKINVDCx5p33_ASAP7_75t_R g680 ( .A(n_12), .Y(n_680) );
INVx1_ASAP7_75t_L g757 ( .A(n_13), .Y(n_757) );
OAI22xp33_ASAP7_75t_L g977 ( .A1(n_14), .A2(n_134), .B1(n_324), .B2(n_538), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g987 ( .A1(n_14), .A2(n_134), .B1(n_517), .B2(n_602), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_15), .A2(n_45), .B1(n_475), .B2(n_517), .Y(n_516) );
OAI22xp33_ASAP7_75t_L g537 ( .A1(n_15), .A2(n_45), .B1(n_324), .B2(n_538), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_16), .A2(n_278), .B1(n_533), .B2(n_588), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_16), .A2(n_278), .B1(n_501), .B2(n_503), .Y(n_655) );
INVx2_ASAP7_75t_L g392 ( .A(n_17), .Y(n_392) );
INVx1_ASAP7_75t_L g1117 ( .A(n_18), .Y(n_1117) );
INVx1_ASAP7_75t_L g1113 ( .A(n_19), .Y(n_1113) );
XNOR2xp5_ASAP7_75t_L g745 ( .A(n_20), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g364 ( .A(n_21), .Y(n_364) );
INVx1_ASAP7_75t_L g1180 ( .A(n_22), .Y(n_1180) );
INVx1_ASAP7_75t_L g1020 ( .A(n_23), .Y(n_1020) );
INVx1_ASAP7_75t_L g1067 ( .A(n_24), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_25), .A2(n_162), .B1(n_1216), .B2(n_1218), .Y(n_1215) );
AOI22xp33_ASAP7_75t_SL g1238 ( .A1(n_25), .A2(n_119), .B1(n_1152), .B2(n_1239), .Y(n_1238) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_26), .A2(n_83), .B1(n_689), .B2(n_1094), .C(n_1097), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_26), .A2(n_42), .B1(n_1150), .B2(n_1152), .Y(n_1149) );
INVx1_ASAP7_75t_L g348 ( .A(n_27), .Y(n_348) );
OAI211xp5_ASAP7_75t_L g441 ( .A1(n_28), .A2(n_442), .B(n_446), .C(n_458), .Y(n_441) );
INVx1_ASAP7_75t_L g499 ( .A(n_28), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g1350 ( .A1(n_29), .A2(n_196), .B1(n_1307), .B2(n_1314), .Y(n_1350) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_30), .A2(n_281), .B1(n_931), .B2(n_1050), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_30), .A2(n_281), .B1(n_502), .B2(n_505), .Y(n_1060) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_31), .Y(n_318) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_31), .B(n_316), .Y(n_1308) );
AOI22xp5_ASAP7_75t_L g1335 ( .A1(n_32), .A2(n_173), .B1(n_1307), .B2(n_1314), .Y(n_1335) );
OAI22xp33_ASAP7_75t_SL g587 ( .A1(n_33), .A2(n_152), .B1(n_533), .B2(n_588), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_33), .A2(n_152), .B1(n_501), .B2(n_592), .Y(n_591) );
OAI222xp33_ASAP7_75t_L g1208 ( .A1(n_34), .A2(n_179), .B1(n_300), .B2(n_813), .C1(n_814), .C2(n_1209), .Y(n_1208) );
OAI222xp33_ASAP7_75t_L g1244 ( .A1(n_34), .A2(n_179), .B1(n_300), .B2(n_453), .C1(n_619), .C2(n_782), .Y(n_1244) );
AOI22xp5_ASAP7_75t_L g1341 ( .A1(n_35), .A2(n_242), .B1(n_1307), .B2(n_1314), .Y(n_1341) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_36), .Y(n_906) );
INVx1_ASAP7_75t_L g1531 ( .A(n_37), .Y(n_1531) );
INVx1_ASAP7_75t_L g974 ( .A(n_38), .Y(n_974) );
INVx1_ASAP7_75t_L g716 ( .A(n_39), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g1330 ( .A1(n_40), .A2(n_107), .B1(n_1307), .B2(n_1314), .Y(n_1330) );
INVxp67_ASAP7_75t_SL g780 ( .A(n_41), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_41), .A2(n_53), .B1(n_813), .B2(n_814), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_42), .A2(n_69), .B1(n_689), .B2(n_1094), .C(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1537 ( .A(n_43), .Y(n_1537) );
INVx1_ASAP7_75t_L g1009 ( .A(n_44), .Y(n_1009) );
AOI22xp5_ASAP7_75t_L g1328 ( .A1(n_46), .A2(n_153), .B1(n_1317), .B2(n_1329), .Y(n_1328) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_47), .A2(n_238), .B1(n_435), .B2(n_873), .Y(n_1051) );
OAI22xp33_ASAP7_75t_SL g1053 ( .A1(n_47), .A2(n_238), .B1(n_477), .B2(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g543 ( .A(n_48), .Y(n_543) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_49), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g1268 ( .A(n_50), .Y(n_1268) );
INVx1_ASAP7_75t_L g1106 ( .A(n_51), .Y(n_1106) );
AOI22xp33_ASAP7_75t_SL g1141 ( .A1(n_51), .A2(n_232), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
INVx1_ASAP7_75t_L g959 ( .A(n_54), .Y(n_959) );
INVx1_ASAP7_75t_L g1188 ( .A(n_55), .Y(n_1188) );
OAI211xp5_ASAP7_75t_SL g518 ( .A1(n_56), .A2(n_483), .B(n_486), .C(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g531 ( .A(n_56), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_57), .A2(n_211), .B1(n_1311), .B2(n_1317), .Y(n_1408) );
OAI211xp5_ASAP7_75t_L g993 ( .A1(n_58), .A2(n_597), .B(n_657), .C(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g1002 ( .A(n_58), .Y(n_1002) );
OAI211xp5_ASAP7_75t_L g863 ( .A1(n_59), .A2(n_864), .B(n_865), .C(n_869), .Y(n_863) );
INVx1_ASAP7_75t_L g886 ( .A(n_59), .Y(n_886) );
OAI22xp33_ASAP7_75t_L g522 ( .A1(n_60), .A2(n_158), .B1(n_501), .B2(n_503), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_60), .A2(n_158), .B1(n_533), .B2(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g957 ( .A(n_61), .Y(n_957) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_62), .Y(n_835) );
INVx1_ASAP7_75t_L g784 ( .A(n_63), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g1525 ( .A1(n_64), .A2(n_71), .B1(n_1526), .B2(n_1527), .Y(n_1525) );
OAI22xp33_ASAP7_75t_L g1565 ( .A1(n_64), .A2(n_71), .B1(n_981), .B2(n_1566), .Y(n_1565) );
OAI222xp33_ASAP7_75t_L g1257 ( .A1(n_65), .A2(n_165), .B1(n_384), .B2(n_734), .C1(n_1258), .C2(n_1259), .Y(n_1257) );
OAI222xp33_ASAP7_75t_L g1284 ( .A1(n_65), .A2(n_165), .B1(n_200), .B2(n_1285), .C1(n_1286), .C2(n_1287), .Y(n_1284) );
INVx1_ASAP7_75t_L g1071 ( .A(n_66), .Y(n_1071) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_67), .A2(n_266), .B1(n_324), .B2(n_538), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g738 ( .A1(n_67), .A2(n_266), .B1(n_517), .B2(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g457 ( .A(n_68), .Y(n_457) );
OAI211xp5_ASAP7_75t_L g482 ( .A1(n_68), .A2(n_483), .B(n_486), .C(n_490), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_69), .A2(n_83), .B1(n_1145), .B2(n_1147), .Y(n_1144) );
INVx1_ASAP7_75t_L g1019 ( .A(n_70), .Y(n_1019) );
INVx1_ASAP7_75t_L g789 ( .A(n_72), .Y(n_789) );
INVx1_ASAP7_75t_L g1015 ( .A(n_73), .Y(n_1015) );
INVx1_ASAP7_75t_L g1544 ( .A(n_74), .Y(n_1544) );
INVx1_ASAP7_75t_L g557 ( .A(n_75), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g1592 ( .A(n_76), .Y(n_1592) );
OAI211xp5_ASAP7_75t_L g1044 ( .A1(n_77), .A2(n_865), .B(n_1045), .C(n_1046), .Y(n_1044) );
INVx1_ASAP7_75t_L g1057 ( .A(n_77), .Y(n_1057) );
INVx1_ASAP7_75t_L g775 ( .A(n_78), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_79), .A2(n_155), .B1(n_1314), .B2(n_1317), .Y(n_1313) );
INVx1_ASAP7_75t_L g631 ( .A(n_80), .Y(n_631) );
XNOR2xp5_ASAP7_75t_L g893 ( .A(n_81), .B(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_82), .A2(n_264), .B1(n_1307), .B2(n_1311), .Y(n_1306) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_84), .A2(n_174), .B1(n_477), .B2(n_502), .Y(n_1110) );
INVx1_ASAP7_75t_L g1123 ( .A(n_84), .Y(n_1123) );
AOI22xp5_ASAP7_75t_L g1353 ( .A1(n_85), .A2(n_140), .B1(n_1317), .B2(n_1326), .Y(n_1353) );
INVx1_ASAP7_75t_L g371 ( .A(n_86), .Y(n_371) );
INVx1_ASAP7_75t_L g1606 ( .A(n_87), .Y(n_1606) );
OAI211xp5_ASAP7_75t_L g1611 ( .A1(n_87), .A2(n_430), .B(n_597), .C(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g556 ( .A(n_88), .Y(n_556) );
INVx1_ASAP7_75t_L g996 ( .A(n_89), .Y(n_996) );
OAI211xp5_ASAP7_75t_L g999 ( .A1(n_89), .A2(n_647), .B(n_1000), .C(n_1001), .Y(n_999) );
INVx1_ASAP7_75t_L g1075 ( .A(n_90), .Y(n_1075) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_91), .A2(n_146), .B1(n_324), .B2(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_91), .A2(n_146), .B1(n_475), .B2(n_478), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_92), .Y(n_833) );
INVx1_ASAP7_75t_L g1118 ( .A(n_93), .Y(n_1118) );
XOR2xp5_ASAP7_75t_L g828 ( .A(n_94), .B(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_95), .A2(n_293), .B1(n_1307), .B2(n_1314), .Y(n_1409) );
INVx1_ASAP7_75t_L g759 ( .A(n_96), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_96), .A2(n_255), .B1(n_800), .B2(n_807), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g910 ( .A(n_97), .Y(n_910) );
INVx1_ASAP7_75t_L g1014 ( .A(n_98), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1523 ( .A1(n_99), .A2(n_125), .B1(n_1253), .B2(n_1524), .Y(n_1523) );
OAI22xp5_ASAP7_75t_L g1558 ( .A1(n_99), .A2(n_125), .B1(n_1559), .B2(n_1560), .Y(n_1558) );
INVx1_ASAP7_75t_L g1048 ( .A(n_100), .Y(n_1048) );
INVx1_ASAP7_75t_L g722 ( .A(n_101), .Y(n_722) );
OAI211xp5_ASAP7_75t_L g1603 ( .A1(n_102), .A2(n_572), .B(n_865), .C(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1613 ( .A(n_102), .Y(n_1613) );
INVx1_ASAP7_75t_L g316 ( .A(n_103), .Y(n_316) );
INVx1_ASAP7_75t_L g952 ( .A(n_104), .Y(n_952) );
INVx1_ASAP7_75t_L g771 ( .A(n_105), .Y(n_771) );
OAI22xp33_ASAP7_75t_L g1608 ( .A1(n_106), .A2(n_262), .B1(n_465), .B2(n_538), .Y(n_1608) );
OAI22xp33_ASAP7_75t_L g1614 ( .A1(n_106), .A2(n_142), .B1(n_502), .B2(n_505), .Y(n_1614) );
XOR2xp5_ASAP7_75t_L g1249 ( .A(n_107), .B(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g585 ( .A(n_108), .Y(n_585) );
INVx1_ASAP7_75t_L g710 ( .A(n_109), .Y(n_710) );
INVx1_ASAP7_75t_L g755 ( .A(n_110), .Y(n_755) );
INVx1_ASAP7_75t_L g616 ( .A(n_111), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g1340 ( .A1(n_112), .A2(n_189), .B1(n_1311), .B2(n_1317), .Y(n_1340) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_113), .A2(n_228), .B1(n_1206), .B2(n_1207), .Y(n_1205) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_113), .A2(n_228), .B1(n_464), .B2(n_791), .Y(n_1243) );
INVx1_ASAP7_75t_L g995 ( .A(n_114), .Y(n_995) );
INVx1_ASAP7_75t_L g1183 ( .A(n_115), .Y(n_1183) );
INVx1_ASAP7_75t_L g561 ( .A(n_116), .Y(n_561) );
INVx1_ASAP7_75t_L g1187 ( .A(n_117), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_118), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_119), .A2(n_253), .B1(n_1094), .B2(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1012 ( .A(n_120), .Y(n_1012) );
INVx1_ASAP7_75t_L g1185 ( .A(n_121), .Y(n_1185) );
AOI31xp33_ASAP7_75t_L g1085 ( .A1(n_122), .A2(n_1086), .A3(n_1109), .B(n_1121), .Y(n_1085) );
NAND2xp33_ASAP7_75t_SL g1137 ( .A(n_122), .B(n_1138), .Y(n_1137) );
INVxp67_ASAP7_75t_SL g1155 ( .A(n_122), .Y(n_1155) );
INVx1_ASAP7_75t_L g1539 ( .A(n_123), .Y(n_1539) );
INVx1_ASAP7_75t_L g351 ( .A(n_124), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_126), .Y(n_679) );
CKINVDCx5p33_ASAP7_75t_R g908 ( .A(n_127), .Y(n_908) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_128), .A2(n_168), .B1(n_538), .B2(n_931), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g938 ( .A1(n_128), .A2(n_161), .B1(n_502), .B2(n_505), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_129), .Y(n_898) );
OAI22xp33_ASAP7_75t_L g997 ( .A1(n_130), .A2(n_145), .B1(n_602), .B2(n_604), .Y(n_997) );
OAI22xp33_ASAP7_75t_L g1004 ( .A1(n_130), .A2(n_145), .B1(n_538), .B2(n_873), .Y(n_1004) );
OAI211xp5_ASAP7_75t_L g583 ( .A1(n_131), .A2(n_525), .B(n_528), .C(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g600 ( .A(n_131), .Y(n_600) );
INVx1_ASAP7_75t_L g586 ( .A(n_132), .Y(n_586) );
OAI211xp5_ASAP7_75t_L g594 ( .A1(n_132), .A2(n_595), .B(n_597), .C(n_598), .Y(n_594) );
INVx1_ASAP7_75t_L g549 ( .A(n_133), .Y(n_549) );
INVx1_ASAP7_75t_L g520 ( .A(n_135), .Y(n_520) );
INVx1_ASAP7_75t_L g373 ( .A(n_136), .Y(n_373) );
INVx1_ASAP7_75t_L g613 ( .A(n_137), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_138), .Y(n_837) );
OAI211xp5_ASAP7_75t_L g729 ( .A1(n_139), .A2(n_527), .B(n_528), .C(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g743 ( .A(n_139), .Y(n_743) );
INVx1_ASAP7_75t_L g731 ( .A(n_141), .Y(n_731) );
OAI22xp33_ASAP7_75t_L g1607 ( .A1(n_142), .A2(n_240), .B1(n_536), .B2(n_873), .Y(n_1607) );
INVx1_ASAP7_75t_L g928 ( .A(n_143), .Y(n_928) );
OAI211xp5_ASAP7_75t_L g934 ( .A1(n_143), .A2(n_430), .B(n_597), .C(n_935), .Y(n_934) );
CKINVDCx5p33_ASAP7_75t_R g1583 ( .A(n_144), .Y(n_1583) );
OAI211xp5_ASAP7_75t_SL g972 ( .A1(n_147), .A2(n_442), .B(n_528), .C(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g986 ( .A(n_147), .Y(n_986) );
INVx1_ASAP7_75t_L g1181 ( .A(n_148), .Y(n_1181) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_149), .A2(n_252), .B1(n_533), .B2(n_588), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_149), .A2(n_252), .B1(n_501), .B2(n_592), .Y(n_744) );
OAI211xp5_ASAP7_75t_L g923 ( .A1(n_150), .A2(n_572), .B(n_865), .C(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g937 ( .A(n_150), .Y(n_937) );
INVx1_ASAP7_75t_L g1011 ( .A(n_151), .Y(n_1011) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_154), .Y(n_842) );
INVx1_ASAP7_75t_L g630 ( .A(n_156), .Y(n_630) );
INVx1_ASAP7_75t_L g721 ( .A(n_157), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g929 ( .A1(n_159), .A2(n_161), .B1(n_536), .B2(n_873), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g933 ( .A1(n_159), .A2(n_168), .B1(n_477), .B2(n_888), .Y(n_933) );
INVx1_ASAP7_75t_L g521 ( .A(n_160), .Y(n_521) );
OAI211xp5_ASAP7_75t_L g524 ( .A1(n_160), .A2(n_525), .B(n_528), .C(n_529), .Y(n_524) );
AOI22xp33_ASAP7_75t_SL g1230 ( .A1(n_162), .A2(n_253), .B1(n_1231), .B2(n_1235), .Y(n_1230) );
OAI22xp33_ASAP7_75t_SL g874 ( .A1(n_163), .A2(n_269), .B1(n_465), .B2(n_538), .Y(n_874) );
INVx1_ASAP7_75t_L g705 ( .A(n_164), .Y(n_705) );
INVx1_ASAP7_75t_L g1177 ( .A(n_166), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_167), .B(n_1310), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_167), .B(n_263), .Y(n_1312) );
INVx2_ASAP7_75t_L g1316 ( .A(n_167), .Y(n_1316) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_169), .Y(n_904) );
INVx1_ASAP7_75t_L g545 ( .A(n_170), .Y(n_545) );
INVx1_ASAP7_75t_L g1521 ( .A(n_171), .Y(n_1521) );
AOI22xp5_ASAP7_75t_L g1324 ( .A1(n_172), .A2(n_222), .B1(n_1307), .B2(n_1317), .Y(n_1324) );
XNOR2xp5_ASAP7_75t_L g943 ( .A(n_173), .B(n_944), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g1127 ( .A1(n_174), .A2(n_245), .B1(n_931), .B2(n_1050), .Y(n_1127) );
INVx1_ASAP7_75t_L g1271 ( .A(n_175), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_176), .A2(n_291), .B1(n_1213), .B2(n_1220), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_176), .A2(n_221), .B1(n_1231), .B2(n_1235), .Y(n_1237) );
XNOR2x2_ASAP7_75t_L g338 ( .A(n_177), .B(n_339), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g1325 ( .A1(n_177), .A2(n_183), .B1(n_1314), .B2(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g1164 ( .A(n_178), .Y(n_1164) );
CKINVDCx5p33_ASAP7_75t_R g1590 ( .A(n_180), .Y(n_1590) );
OAI211xp5_ASAP7_75t_L g1519 ( .A1(n_181), .A2(n_458), .B(n_1184), .C(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1564 ( .A(n_181), .Y(n_1564) );
INVx1_ASAP7_75t_L g1047 ( .A(n_182), .Y(n_1047) );
XOR2x2_ASAP7_75t_L g1041 ( .A(n_184), .B(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g956 ( .A(n_185), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_186), .Y(n_649) );
OAI211xp5_ASAP7_75t_L g1252 ( .A1(n_187), .A2(n_1253), .B(n_1254), .C(n_1263), .Y(n_1252) );
INVx1_ASAP7_75t_L g1290 ( .A(n_187), .Y(n_1290) );
INVx1_ASAP7_75t_L g711 ( .A(n_188), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_190), .A2(n_207), .B1(n_501), .B2(n_981), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_190), .A2(n_207), .B1(n_464), .B2(n_466), .Y(n_1003) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_191), .A2(n_254), .B1(n_324), .B2(n_538), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g601 ( .A1(n_191), .A2(n_254), .B1(n_602), .B2(n_604), .Y(n_601) );
INVx2_ASAP7_75t_L g391 ( .A(n_192), .Y(n_391) );
INVx1_ASAP7_75t_L g428 ( .A(n_192), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g1584 ( .A(n_193), .Y(n_1584) );
AOI22xp5_ASAP7_75t_L g1354 ( .A1(n_194), .A2(n_299), .B1(n_1307), .B2(n_1314), .Y(n_1354) );
OAI22xp33_ASAP7_75t_L g1160 ( .A1(n_195), .A2(n_244), .B1(n_931), .B2(n_1050), .Y(n_1160) );
OAI22xp5_ASAP7_75t_SL g1167 ( .A1(n_195), .A2(n_219), .B1(n_477), .B2(n_502), .Y(n_1167) );
XOR2xp5_ASAP7_75t_L g1198 ( .A(n_197), .B(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1262 ( .A(n_198), .Y(n_1262) );
OAI22xp5_ASAP7_75t_L g1288 ( .A1(n_198), .A2(n_225), .B1(n_502), .B2(n_505), .Y(n_1288) );
INVx1_ASAP7_75t_L g1255 ( .A(n_200), .Y(n_1255) );
BUFx3_ASAP7_75t_L g398 ( .A(n_201), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g1594 ( .A(n_202), .Y(n_1594) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_203), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_204), .Y(n_913) );
XOR2xp5_ASAP7_75t_L g700 ( .A(n_205), .B(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_206), .A2(n_221), .B1(n_1114), .B2(n_1213), .Y(n_1212) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_206), .A2(n_291), .B1(n_1228), .B2(n_1229), .Y(n_1227) );
OA22x2_ASAP7_75t_L g989 ( .A1(n_208), .A2(n_990), .B1(n_1032), .B2(n_1033), .Y(n_989) );
INVxp67_ASAP7_75t_L g1033 ( .A(n_208), .Y(n_1033) );
INVx1_ASAP7_75t_L g764 ( .A(n_209), .Y(n_764) );
INVx1_ASAP7_75t_L g651 ( .A(n_210), .Y(n_651) );
OAI211xp5_ASAP7_75t_L g656 ( .A1(n_210), .A2(n_597), .B(n_657), .C(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g1267 ( .A(n_212), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_212), .B(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g706 ( .A(n_213), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_214), .Y(n_902) );
INVx1_ASAP7_75t_L g1535 ( .A(n_215), .Y(n_1535) );
CKINVDCx5p33_ASAP7_75t_R g1587 ( .A(n_216), .Y(n_1587) );
INVx1_ASAP7_75t_L g618 ( .A(n_217), .Y(n_618) );
INVx1_ASAP7_75t_L g1163 ( .A(n_218), .Y(n_1163) );
OAI22xp33_ASAP7_75t_L g1165 ( .A1(n_219), .A2(n_247), .B1(n_435), .B2(n_873), .Y(n_1165) );
CKINVDCx5p33_ASAP7_75t_R g674 ( .A(n_220), .Y(n_674) );
INVx1_ASAP7_75t_L g769 ( .A(n_223), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_223), .A2(n_265), .B1(n_798), .B2(n_800), .Y(n_797) );
INVx1_ASAP7_75t_L g1069 ( .A(n_224), .Y(n_1069) );
INVx1_ASAP7_75t_L g1264 ( .A(n_225), .Y(n_1264) );
BUFx3_ASAP7_75t_L g332 ( .A(n_226), .Y(n_332) );
INVx1_ASAP7_75t_L g438 ( .A(n_226), .Y(n_438) );
INVx1_ASAP7_75t_L g451 ( .A(n_227), .Y(n_451) );
XOR2x2_ASAP7_75t_L g513 ( .A(n_229), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g1064 ( .A(n_231), .Y(n_1064) );
AOI22xp5_ASAP7_75t_L g1087 ( .A1(n_232), .A2(n_250), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
INVx1_ASAP7_75t_L g386 ( .A(n_233), .Y(n_386) );
INVx1_ASAP7_75t_L g1203 ( .A(n_234), .Y(n_1203) );
OAI211xp5_ASAP7_75t_L g1161 ( .A1(n_235), .A2(n_619), .B(n_865), .C(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1172 ( .A(n_235), .Y(n_1172) );
INVx1_ASAP7_75t_L g1522 ( .A(n_236), .Y(n_1522) );
OAI211xp5_ASAP7_75t_L g1561 ( .A1(n_236), .A2(n_401), .B(n_486), .C(n_1562), .Y(n_1561) );
CKINVDCx5p33_ASAP7_75t_R g840 ( .A(n_237), .Y(n_840) );
INVx1_ASAP7_75t_L g1540 ( .A(n_239), .Y(n_1540) );
OAI22xp33_ASAP7_75t_L g1610 ( .A1(n_240), .A2(n_262), .B1(n_477), .B2(n_888), .Y(n_1610) );
CKINVDCx5p33_ASAP7_75t_R g843 ( .A(n_241), .Y(n_843) );
XOR2x2_ASAP7_75t_L g579 ( .A(n_242), .B(n_580), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_243), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g1173 ( .A1(n_244), .A2(n_247), .B1(n_505), .B2(n_888), .Y(n_1173) );
OAI22xp5_ASAP7_75t_L g1119 ( .A1(n_245), .A2(n_282), .B1(n_505), .B2(n_888), .Y(n_1119) );
INVx1_ASAP7_75t_L g400 ( .A(n_246), .Y(n_400) );
INVx1_ASAP7_75t_L g406 ( .A(n_246), .Y(n_406) );
INVx1_ASAP7_75t_L g385 ( .A(n_248), .Y(n_385) );
INVx1_ASAP7_75t_L g359 ( .A(n_249), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_250), .A2(n_284), .B1(n_1145), .B2(n_1147), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_251), .A2(n_297), .B1(n_464), .B2(n_466), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g500 ( .A1(n_251), .A2(n_297), .B1(n_501), .B2(n_503), .Y(n_500) );
INVx1_ASAP7_75t_L g767 ( .A(n_255), .Y(n_767) );
INVx1_ASAP7_75t_L g870 ( .A(n_256), .Y(n_870) );
OAI211xp5_ASAP7_75t_SL g878 ( .A1(n_256), .A2(n_486), .B(n_813), .C(n_879), .Y(n_878) );
XNOR2xp5_ASAP7_75t_L g1577 ( .A(n_257), .B(n_1578), .Y(n_1577) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_258), .A2(n_260), .B1(n_324), .B2(n_538), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g662 ( .A1(n_258), .A2(n_260), .B1(n_517), .B2(n_602), .Y(n_662) );
INVx1_ASAP7_75t_L g551 ( .A(n_259), .Y(n_551) );
AOI22xp5_ASAP7_75t_SL g1349 ( .A1(n_261), .A2(n_305), .B1(n_1317), .B2(n_1326), .Y(n_1349) );
AOI22xp5_ASAP7_75t_L g1515 ( .A1(n_261), .A2(n_1516), .B1(n_1517), .B2(n_1567), .Y(n_1515) );
INVxp67_ASAP7_75t_SL g1567 ( .A(n_261), .Y(n_1567) );
AOI22xp33_ASAP7_75t_L g1573 ( .A1(n_261), .A2(n_1574), .B1(n_1576), .B2(n_1615), .Y(n_1573) );
INVx1_ASAP7_75t_L g1310 ( .A(n_263), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_263), .B(n_1316), .Y(n_1318) );
INVx1_ASAP7_75t_L g751 ( .A(n_265), .Y(n_751) );
INVx1_ASAP7_75t_L g1065 ( .A(n_267), .Y(n_1065) );
CKINVDCx5p33_ASAP7_75t_R g1588 ( .A(n_268), .Y(n_1588) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_269), .A2(n_302), .B1(n_502), .B2(n_505), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_270), .Y(n_666) );
INVx1_ASAP7_75t_L g1202 ( .A(n_271), .Y(n_1202) );
INVx1_ASAP7_75t_L g1074 ( .A(n_272), .Y(n_1074) );
INVx1_ASAP7_75t_L g774 ( .A(n_273), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_274), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g1273 ( .A(n_275), .Y(n_1273) );
INVx1_ASAP7_75t_L g1178 ( .A(n_276), .Y(n_1178) );
INVx1_ASAP7_75t_L g975 ( .A(n_277), .Y(n_975) );
OAI211xp5_ASAP7_75t_SL g982 ( .A1(n_277), .A2(n_486), .B(n_983), .C(n_985), .Y(n_982) );
XOR2x2_ASAP7_75t_L g1157 ( .A(n_279), .B(n_1158), .Y(n_1157) );
OAI211xp5_ASAP7_75t_L g646 ( .A1(n_280), .A2(n_527), .B(n_647), .C(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g661 ( .A(n_280), .Y(n_661) );
INVxp67_ASAP7_75t_SL g1125 ( .A(n_282), .Y(n_1125) );
INVx1_ASAP7_75t_L g732 ( .A(n_283), .Y(n_732) );
OAI211xp5_ASAP7_75t_L g741 ( .A1(n_283), .A2(n_596), .B(n_597), .C(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g1103 ( .A(n_284), .Y(n_1103) );
INVx1_ASAP7_75t_L g1008 ( .A(n_285), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_286), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_287), .Y(n_668) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_288), .Y(n_328) );
INVx1_ASAP7_75t_L g1533 ( .A(n_289), .Y(n_1533) );
INVx1_ASAP7_75t_L g1545 ( .A(n_290), .Y(n_1545) );
INVx1_ASAP7_75t_L g624 ( .A(n_292), .Y(n_624) );
INVx1_ASAP7_75t_L g715 ( .A(n_294), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_295), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g1605 ( .A(n_296), .Y(n_1605) );
CKINVDCx5p33_ASAP7_75t_R g871 ( .A(n_298), .Y(n_871) );
XOR2x2_ASAP7_75t_L g643 ( .A(n_301), .B(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g345 ( .A(n_303), .Y(n_345) );
INVx1_ASAP7_75t_L g381 ( .A(n_303), .Y(n_381) );
INVx1_ASAP7_75t_L g427 ( .A(n_303), .Y(n_427) );
INVx1_ASAP7_75t_L g948 ( .A(n_304), .Y(n_948) );
INVx1_ASAP7_75t_L g951 ( .A(n_306), .Y(n_951) );
INVx1_ASAP7_75t_L g626 ( .A(n_307), .Y(n_626) );
AOI21xp33_ASAP7_75t_L g1274 ( .A1(n_308), .A2(n_1145), .B(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1293 ( .A(n_308), .Y(n_1293) );
INVx1_ASAP7_75t_L g560 ( .A(n_309), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g1595 ( .A(n_310), .Y(n_1595) );
CKINVDCx5p33_ASAP7_75t_R g1260 ( .A(n_311), .Y(n_1260) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_333), .B(n_1300), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_319), .Y(n_313) );
INVx1_ASAP7_75t_L g1572 ( .A(n_314), .Y(n_1572) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g1575 ( .A(n_315), .B(n_318), .Y(n_1575) );
INVx1_ASAP7_75t_L g1616 ( .A(n_315), .Y(n_1616) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g1618 ( .A(n_318), .B(n_1616), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_323), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g470 ( .A(n_321), .B(n_471), .Y(n_470) );
AOI21xp5_ASAP7_75t_SL g1251 ( .A1(n_321), .A2(n_1252), .B(n_1265), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1571 ( .A(n_321), .B(n_1572), .Y(n_1571) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g376 ( .A(n_322), .B(n_332), .Y(n_376) );
AND2x4_ASAP7_75t_L g1276 ( .A(n_322), .B(n_331), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_323), .A2(n_436), .B1(n_774), .B2(n_775), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_323), .A2(n_436), .B1(n_1202), .B2(n_1203), .Y(n_1241) );
INVx1_ASAP7_75t_L g1524 ( .A(n_323), .Y(n_1524) );
AND2x4_ASAP7_75t_SL g1570 ( .A(n_323), .B(n_1571), .Y(n_1570) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x6_ASAP7_75t_L g324 ( .A(n_325), .B(n_330), .Y(n_324) );
OR2x6_ASAP7_75t_L g465 ( .A(n_325), .B(n_437), .Y(n_465) );
BUFx4f_ASAP7_75t_L g612 ( .A(n_325), .Y(n_612) );
INVx1_ASAP7_75t_L g859 ( .A(n_325), .Y(n_859) );
OR2x2_ASAP7_75t_L g931 ( .A(n_325), .B(n_437), .Y(n_931) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx4f_ASAP7_75t_L g350 ( .A(n_326), .Y(n_350) );
INVx3_ASAP7_75t_L g384 ( .A(n_326), .Y(n_384) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx2_ASAP7_75t_L g357 ( .A(n_328), .Y(n_357) );
INVx2_ASAP7_75t_L g363 ( .A(n_328), .Y(n_363) );
NAND2x1_ASAP7_75t_L g366 ( .A(n_328), .B(n_329), .Y(n_366) );
AND2x2_ASAP7_75t_L g439 ( .A(n_328), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g456 ( .A(n_328), .Y(n_456) );
AND2x2_ASAP7_75t_L g462 ( .A(n_328), .B(n_329), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_329), .B(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g362 ( .A(n_329), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g440 ( .A(n_329), .Y(n_440) );
BUFx2_ASAP7_75t_L g450 ( .A(n_329), .Y(n_450) );
INVx1_ASAP7_75t_L g788 ( .A(n_329), .Y(n_788) );
AND2x2_ASAP7_75t_L g802 ( .A(n_329), .B(n_357), .Y(n_802) );
OR2x6_ASAP7_75t_L g873 ( .A(n_330), .B(n_384), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g1259 ( .A1(n_330), .A2(n_1260), .B1(n_1261), .B2(n_1262), .Y(n_1259) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g460 ( .A(n_331), .Y(n_460) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_L g449 ( .A(n_332), .Y(n_449) );
AND2x4_ASAP7_75t_L g454 ( .A(n_332), .B(n_455), .Y(n_454) );
XNOR2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_1036), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_825), .B1(n_1034), .B2(n_1035), .Y(n_334) );
INVx2_ASAP7_75t_SL g1034 ( .A(n_335), .Y(n_1034) );
XOR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_576), .Y(n_335) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_512), .B(n_575), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g575 ( .A(n_338), .B(n_513), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_433), .C(n_473), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_387), .Y(n_340) );
OAI33xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_347), .A3(n_358), .B1(n_367), .B2(n_374), .B3(n_382), .Y(n_341) );
OAI33xp33_ASAP7_75t_L g562 ( .A1(n_342), .A2(n_563), .A3(n_566), .B1(n_571), .B2(n_573), .B3(n_574), .Y(n_562) );
OAI33xp33_ASAP7_75t_L g1006 ( .A1(n_342), .A2(n_573), .A3(n_1007), .B1(n_1010), .B2(n_1013), .B3(n_1016), .Y(n_1006) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g609 ( .A(n_343), .Y(n_609) );
INVx1_ASAP7_75t_L g669 ( .A(n_343), .Y(n_669) );
INVx2_ASAP7_75t_L g795 ( .A(n_343), .Y(n_795) );
INVx4_ASAP7_75t_L g1140 ( .A(n_343), .Y(n_1140) );
INVx1_ASAP7_75t_L g1547 ( .A(n_343), .Y(n_1547) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
OR2x2_ASAP7_75t_L g847 ( .A(n_344), .B(n_848), .Y(n_847) );
OR2x6_ASAP7_75t_L g1108 ( .A(n_344), .B(n_848), .Y(n_1108) );
INVx1_ASAP7_75t_L g1280 ( .A(n_344), .Y(n_1280) );
BUFx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g1099 ( .A(n_345), .Y(n_1099) );
OAI22xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_349), .B1(n_351), .B2(n_352), .Y(n_347) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_348), .A2(n_371), .B1(n_394), .B2(n_401), .Y(n_393) );
INVx2_ASAP7_75t_SL g565 ( .A(n_349), .Y(n_565) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_350), .Y(n_629) );
INVx4_ASAP7_75t_L g851 ( .A(n_350), .Y(n_851) );
OAI22xp33_ASAP7_75t_L g429 ( .A1(n_351), .A2(n_373), .B1(n_394), .B2(n_430), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_352), .A2(n_383), .B1(n_385), .B2(n_386), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_352), .A2(n_543), .B1(n_560), .B2(n_564), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_352), .A2(n_551), .B1(n_557), .B2(n_564), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_352), .A2(n_666), .B1(n_667), .B2(n_668), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g678 ( .A1(n_352), .A2(n_667), .B1(n_679), .B2(n_680), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g947 ( .A1(n_352), .A2(n_383), .B1(n_948), .B2(n_949), .Y(n_947) );
INVx6_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx5_ASAP7_75t_L g614 ( .A(n_353), .Y(n_614) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx4_ASAP7_75t_L g852 ( .A(n_354), .Y(n_852) );
INVx2_ASAP7_75t_SL g899 ( .A(n_354), .Y(n_899) );
INVx2_ASAP7_75t_L g912 ( .A(n_354), .Y(n_912) );
INVx1_ASAP7_75t_L g961 ( .A(n_354), .Y(n_961) );
INVx1_ASAP7_75t_L g1078 ( .A(n_354), .Y(n_1078) );
INVx8_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g468 ( .A(n_355), .B(n_449), .Y(n_468) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_355), .B(n_460), .Y(n_1050) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_364), .B2(n_365), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_359), .A2(n_385), .B1(n_409), .B2(n_414), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g796 ( .A1(n_360), .A2(n_527), .B1(n_757), .B2(n_764), .C(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g955 ( .A(n_360), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g1551 ( .A1(n_360), .A2(n_864), .B1(n_1535), .B2(n_1539), .Y(n_1551) );
OAI22xp5_ASAP7_75t_L g1552 ( .A1(n_360), .A2(n_864), .B1(n_1533), .B2(n_1545), .Y(n_1552) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g568 ( .A(n_361), .Y(n_568) );
INVx2_ASAP7_75t_L g903 ( .A(n_361), .Y(n_903) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g370 ( .A(n_362), .Y(n_370) );
BUFx3_ASAP7_75t_L g623 ( .A(n_362), .Y(n_623) );
INVx1_ASAP7_75t_L g673 ( .A(n_362), .Y(n_673) );
BUFx2_ASAP7_75t_L g1600 ( .A(n_362), .Y(n_1600) );
AND2x2_ASAP7_75t_L g787 ( .A(n_363), .B(n_788), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_364), .A2(n_386), .B1(n_419), .B2(n_420), .Y(n_418) );
BUFx2_ASAP7_75t_SL g372 ( .A(n_365), .Y(n_372) );
BUFx3_ASAP7_75t_L g527 ( .A(n_365), .Y(n_527) );
INVx2_ASAP7_75t_SL g620 ( .A(n_365), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_365), .A2(n_902), .B1(n_903), .B2(n_904), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_365), .A2(n_854), .B1(n_1065), .B2(n_1075), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g1599 ( .A1(n_365), .A2(n_1584), .B1(n_1595), .B2(n_1600), .Y(n_1599) );
BUFx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_366), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B1(n_372), .B2(n_373), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g950 ( .A1(n_368), .A2(n_619), .B1(n_951), .B2(n_952), .Y(n_950) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx4_ASAP7_75t_L g617 ( .A(n_369), .Y(n_617) );
INVx4_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_372), .A2(n_954), .B1(n_956), .B2(n_957), .Y(n_953) );
OAI33xp33_ASAP7_75t_L g723 ( .A1(n_374), .A2(n_608), .A3(n_724), .B1(n_725), .B2(n_726), .B3(n_727), .Y(n_723) );
OAI33xp33_ASAP7_75t_L g946 ( .A1(n_374), .A2(n_608), .A3(n_947), .B1(n_950), .B2(n_953), .B3(n_958), .Y(n_946) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_375), .Y(n_573) );
AOI33xp33_ASAP7_75t_L g1225 ( .A1(n_375), .A2(n_1226), .A3(n_1227), .B1(n_1230), .B2(n_1237), .B3(n_1238), .Y(n_1225) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
AND2x2_ASAP7_75t_SL g861 ( .A(n_376), .B(n_379), .Y(n_861) );
OAI221xp5_ASAP7_75t_L g1269 ( .A1(n_376), .A2(n_567), .B1(n_1000), .B2(n_1270), .C(n_1271), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1555 ( .A(n_376), .B(n_377), .Y(n_1555) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g389 ( .A(n_379), .B(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_379), .Y(n_511) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g472 ( .A(n_380), .Y(n_472) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_383), .A2(n_959), .B1(n_960), .B2(n_962), .Y(n_958) );
BUFx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_SL g1018 ( .A(n_384), .Y(n_1018) );
OAI33xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_393), .A3(n_408), .B1(n_418), .B2(n_422), .B3(n_429), .Y(n_387) );
OAI33xp33_ASAP7_75t_L g632 ( .A1(n_388), .A2(n_558), .A3(n_633), .B1(n_637), .B2(n_641), .B3(n_642), .Y(n_632) );
OAI33xp33_ASAP7_75t_L g703 ( .A1(n_388), .A2(n_704), .A3(n_709), .B1(n_712), .B2(n_717), .B3(n_720), .Y(n_703) );
BUFx4f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx2_ASAP7_75t_L g541 ( .A(n_389), .Y(n_541) );
BUFx8_ASAP7_75t_L g682 ( .A(n_389), .Y(n_682) );
BUFx4f_ASAP7_75t_L g749 ( .A(n_389), .Y(n_749) );
NAND2xp33_ASAP7_75t_SL g390 ( .A(n_391), .B(n_392), .Y(n_390) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_391), .Y(n_509) );
AND3x4_ASAP7_75t_L g1098 ( .A(n_391), .B(n_494), .C(n_1099), .Y(n_1098) );
INVx3_ASAP7_75t_L g425 ( .A(n_392), .Y(n_425) );
BUFx3_ASAP7_75t_L g494 ( .A(n_392), .Y(n_494) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g685 ( .A(n_396), .Y(n_685) );
INVx1_ASAP7_75t_L g695 ( .A(n_396), .Y(n_695) );
BUFx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x4_ASAP7_75t_L g477 ( .A(n_397), .B(n_425), .Y(n_477) );
OR2x4_ASAP7_75t_L g502 ( .A(n_397), .B(n_480), .Y(n_502) );
BUFx3_ASAP7_75t_L g544 ( .A(n_397), .Y(n_544) );
INVx2_ASAP7_75t_L g636 ( .A(n_397), .Y(n_636) );
BUFx4f_ASAP7_75t_L g834 ( .A(n_397), .Y(n_834) );
OR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_398), .Y(n_407) );
INVx2_ASAP7_75t_L g413 ( .A(n_398), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_398), .B(n_406), .Y(n_417) );
AND2x4_ASAP7_75t_L g488 ( .A(n_398), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g1092 ( .A(n_399), .Y(n_1092) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g412 ( .A(n_400), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g1543 ( .A1(n_401), .A2(n_1532), .B1(n_1544), .B2(n_1545), .Y(n_1543) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_403), .Y(n_770) );
OAI22xp33_ASAP7_75t_L g844 ( .A1(n_403), .A2(n_834), .B1(n_845), .B2(n_846), .Y(n_844) );
OAI22xp33_ASAP7_75t_L g921 ( .A1(n_403), .A2(n_754), .B1(n_900), .B2(n_908), .Y(n_921) );
OAI22xp33_ASAP7_75t_L g1073 ( .A1(n_403), .A2(n_834), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_403), .A2(n_754), .B1(n_1177), .B2(n_1183), .Y(n_1190) );
OAI22xp33_ASAP7_75t_L g1593 ( .A1(n_403), .A2(n_754), .B1(n_1594), .B2(n_1595), .Y(n_1593) );
BUFx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g432 ( .A(n_404), .Y(n_432) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_404), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
BUFx2_ASAP7_75t_L g498 ( .A(n_405), .Y(n_498) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g489 ( .A(n_406), .Y(n_489) );
BUFx2_ASAP7_75t_L g495 ( .A(n_407), .Y(n_495) );
INVx2_ASAP7_75t_L g884 ( .A(n_407), .Y(n_884) );
AND2x4_ASAP7_75t_L g1096 ( .A(n_407), .B(n_882), .Y(n_1096) );
BUFx3_ASAP7_75t_L g550 ( .A(n_409), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_409), .A2(n_414), .B1(n_618), .B2(n_631), .Y(n_641) );
INVx8_ASAP7_75t_L g714 ( .A(n_409), .Y(n_714) );
INVx5_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_SL g419 ( .A(n_410), .Y(n_419) );
INVx3_ASAP7_75t_L g555 ( .A(n_410), .Y(n_555) );
INVx2_ASAP7_75t_SL g758 ( .A(n_410), .Y(n_758) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_411), .Y(n_481) );
BUFx8_ASAP7_75t_L g763 ( .A(n_411), .Y(n_763) );
INVx2_ASAP7_75t_L g1030 ( .A(n_411), .Y(n_1030) );
AND2x4_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_413), .B(n_1092), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_414), .A2(n_549), .B1(n_550), .B2(n_551), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_414), .A2(n_713), .B1(n_715), .B2(n_716), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g1024 ( .A1(n_414), .A2(n_1011), .B1(n_1019), .B2(n_1025), .Y(n_1024) );
OAI221xp5_ASAP7_75t_L g1297 ( .A1(n_414), .A2(n_1268), .B1(n_1273), .B2(n_1298), .C(n_1299), .Y(n_1297) );
CKINVDCx8_ASAP7_75t_R g414 ( .A(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g760 ( .A(n_415), .Y(n_760) );
INVx3_ASAP7_75t_L g919 ( .A(n_415), .Y(n_919) );
INVx3_ASAP7_75t_L g1193 ( .A(n_415), .Y(n_1193) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g766 ( .A(n_416), .Y(n_766) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g421 ( .A(n_417), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_419), .A2(n_616), .B1(n_630), .B2(n_638), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_419), .A2(n_760), .B1(n_904), .B2(n_913), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_420), .A2(n_553), .B1(n_556), .B2(n_557), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_420), .A2(n_951), .B1(n_959), .B2(n_967), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_420), .A2(n_952), .B1(n_962), .B2(n_969), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_420), .A2(n_1012), .B1(n_1020), .B2(n_1028), .Y(n_1027) );
BUFx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OR2x6_ASAP7_75t_L g505 ( .A(n_421), .B(n_425), .Y(n_505) );
INVx1_ASAP7_75t_L g640 ( .A(n_421), .Y(n_640) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_423), .Y(n_558) );
INVx2_ASAP7_75t_L g692 ( .A(n_423), .Y(n_692) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx3_ASAP7_75t_L g719 ( .A(n_424), .Y(n_719) );
NAND3x1_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .C(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g480 ( .A(n_425), .Y(n_480) );
AND2x4_ASAP7_75t_L g487 ( .A(n_425), .B(n_488), .Y(n_487) );
NAND2x1p5_ASAP7_75t_L g848 ( .A(n_425), .B(n_428), .Y(n_848) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_430), .A2(n_544), .B1(n_560), .B2(n_561), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_430), .A2(n_611), .B1(n_624), .B2(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g708 ( .A(n_432), .Y(n_708) );
INVx1_ASAP7_75t_L g984 ( .A(n_432), .Y(n_984) );
OAI31xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_441), .A3(n_463), .B(n_469), .Y(n_433) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_436), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g1122 ( .A1(n_436), .A2(n_1123), .B1(n_1124), .B2(n_1125), .Y(n_1122) );
INVx3_ASAP7_75t_SL g1253 ( .A(n_436), .Y(n_1253) );
AND2x4_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx6f_ASAP7_75t_L g1146 ( .A(n_439), .Y(n_1146) );
INVx2_ASAP7_75t_L g1234 ( .A(n_439), .Y(n_1234) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_444), .A2(n_672), .B1(n_676), .B2(n_677), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g1013 ( .A1(n_444), .A2(n_672), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
BUFx4f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx4_ASAP7_75t_L g570 ( .A(n_445), .Y(n_570) );
BUFx4f_ASAP7_75t_L g625 ( .A(n_445), .Y(n_625) );
BUFx4f_ASAP7_75t_L g864 ( .A(n_445), .Y(n_864) );
BUFx6f_ASAP7_75t_L g907 ( .A(n_445), .Y(n_907) );
BUFx4f_ASAP7_75t_L g1184 ( .A(n_445), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_451), .B1(n_452), .B2(n_457), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_447), .A2(n_927), .B1(n_974), .B2(n_975), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1520 ( .A1(n_447), .A2(n_927), .B1(n_1521), .B2(n_1522), .Y(n_1520) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_448), .A2(n_454), .B1(n_585), .B2(n_586), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_448), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
INVx1_ASAP7_75t_L g782 ( .A(n_448), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_448), .A2(n_927), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_448), .A2(n_927), .B1(n_1163), .B2(n_1164), .Y(n_1162) );
AND2x4_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
AND2x2_ASAP7_75t_L g530 ( .A(n_449), .B(n_450), .Y(n_530) );
AND2x2_ASAP7_75t_L g785 ( .A(n_449), .B(n_786), .Y(n_785) );
O2A1O1Ixp33_ASAP7_75t_L g1254 ( .A1(n_449), .A2(n_1255), .B(n_1256), .C(n_1257), .Y(n_1254) );
INVx1_ASAP7_75t_L g1261 ( .A(n_449), .Y(n_1261) );
AND2x2_ASAP7_75t_L g925 ( .A(n_450), .B(n_460), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_451), .A2(n_491), .B1(n_496), .B2(n_499), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_452), .A2(n_520), .B1(n_530), .B2(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g650 ( .A(n_453), .Y(n_650) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g734 ( .A(n_454), .Y(n_734) );
BUFx3_ASAP7_75t_L g927 ( .A(n_454), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_454), .A2(n_925), .B1(n_1113), .B2(n_1117), .Y(n_1129) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g528 ( .A(n_459), .Y(n_528) );
INVx3_ASAP7_75t_L g647 ( .A(n_459), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g776 ( .A1(n_459), .A2(n_777), .B(n_780), .C(n_781), .Y(n_776) );
NOR3xp33_ASAP7_75t_L g1242 ( .A(n_459), .B(n_1243), .C(n_1244), .Y(n_1242) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
AND2x2_ASAP7_75t_L g866 ( .A(n_460), .B(n_867), .Y(n_866) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_461), .Y(n_779) );
BUFx3_ASAP7_75t_L g1147 ( .A(n_461), .Y(n_1147) );
BUFx3_ASAP7_75t_L g1256 ( .A(n_461), .Y(n_1256) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g868 ( .A(n_462), .Y(n_868) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g533 ( .A(n_465), .Y(n_533) );
HB1xp67_ASAP7_75t_L g1526 ( .A(n_465), .Y(n_1526) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g588 ( .A(n_467), .Y(n_588) );
INVx1_ASAP7_75t_L g1527 ( .A(n_467), .Y(n_1527) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g536 ( .A(n_468), .Y(n_536) );
INVx1_ASAP7_75t_L g792 ( .A(n_468), .Y(n_792) );
OAI31xp33_ASAP7_75t_L g523 ( .A1(n_469), .A2(n_524), .A3(n_532), .B(n_537), .Y(n_523) );
OAI31xp33_ASAP7_75t_SL g728 ( .A1(n_469), .A2(n_729), .A3(n_735), .B(n_736), .Y(n_728) );
OAI31xp33_ASAP7_75t_L g971 ( .A1(n_469), .A2(n_972), .A3(n_976), .B(n_977), .Y(n_971) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_SL g589 ( .A(n_470), .Y(n_589) );
INVx1_ASAP7_75t_L g793 ( .A(n_470), .Y(n_793) );
BUFx2_ASAP7_75t_L g875 ( .A(n_470), .Y(n_875) );
OAI31xp33_ASAP7_75t_L g1159 ( .A1(n_470), .A2(n_1160), .A3(n_1161), .B(n_1165), .Y(n_1159) );
OAI31xp33_ASAP7_75t_L g1518 ( .A1(n_470), .A2(n_1519), .A3(n_1523), .B(n_1525), .Y(n_1518) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI31xp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_482), .A3(n_500), .B(n_506), .Y(n_473) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g603 ( .A(n_477), .Y(n_603) );
INVx1_ASAP7_75t_L g740 ( .A(n_477), .Y(n_740) );
INVx2_ASAP7_75t_SL g816 ( .A(n_477), .Y(n_816) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g517 ( .A(n_479), .Y(n_517) );
INVx1_ASAP7_75t_L g604 ( .A(n_479), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_479), .A2(n_774), .B1(n_775), .B2(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g1054 ( .A(n_479), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_479), .A2(n_816), .B1(n_1202), .B2(n_1203), .Y(n_1201) );
INVx2_ASAP7_75t_L g1560 ( .A(n_479), .Y(n_1560) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
AND2x2_ASAP7_75t_L g889 ( .A(n_480), .B(n_481), .Y(n_889) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_481), .Y(n_689) );
INVx2_ASAP7_75t_L g691 ( .A(n_481), .Y(n_691) );
INVx2_ASAP7_75t_L g918 ( .A(n_481), .Y(n_918) );
INVx2_ASAP7_75t_L g969 ( .A(n_481), .Y(n_969) );
BUFx6f_ASAP7_75t_L g1026 ( .A(n_481), .Y(n_1026) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_483), .A2(n_668), .B1(n_677), .B2(n_694), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g720 ( .A1(n_483), .A2(n_634), .B1(n_721), .B2(n_722), .Y(n_720) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g596 ( .A(n_484), .Y(n_596) );
INVx1_ASAP7_75t_L g1195 ( .A(n_484), .Y(n_1195) );
INVx1_ASAP7_75t_L g1209 ( .A(n_484), .Y(n_1209) );
INVx2_ASAP7_75t_L g1285 ( .A(n_484), .Y(n_1285) );
INVx4_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g547 ( .A(n_485), .Y(n_547) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_485), .Y(n_659) );
HB1xp67_ASAP7_75t_L g965 ( .A(n_485), .Y(n_965) );
CKINVDCx8_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
CKINVDCx8_ASAP7_75t_R g597 ( .A(n_487), .Y(n_597) );
AOI211xp5_ASAP7_75t_L g809 ( .A1(n_487), .A2(n_810), .B(n_811), .C(n_812), .Y(n_809) );
NOR3xp33_ASAP7_75t_L g1204 ( .A(n_487), .B(n_1205), .C(n_1208), .Y(n_1204) );
NOR3xp33_ASAP7_75t_L g1283 ( .A(n_487), .B(n_1284), .C(n_1288), .Y(n_1283) );
BUFx3_ASAP7_75t_L g811 ( .A(n_488), .Y(n_811) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_488), .Y(n_1088) );
INVx2_ASAP7_75t_L g1115 ( .A(n_488), .Y(n_1115) );
BUFx2_ASAP7_75t_L g1170 ( .A(n_488), .Y(n_1170) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_488), .Y(n_1221) );
INVx1_ASAP7_75t_L g882 ( .A(n_489), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_491), .A2(n_496), .B1(n_520), .B2(n_521), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_491), .A2(n_496), .B1(n_974), .B2(n_986), .Y(n_985) );
BUFx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx3_ASAP7_75t_L g1563 ( .A(n_492), .Y(n_1563) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x4_ASAP7_75t_L g497 ( .A(n_493), .B(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g599 ( .A(n_493), .B(n_495), .Y(n_599) );
AND2x2_ASAP7_75t_L g885 ( .A(n_493), .B(n_498), .Y(n_885) );
AND2x4_ASAP7_75t_L g936 ( .A(n_493), .B(n_495), .Y(n_936) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g880 ( .A(n_494), .B(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g1562 ( .A1(n_496), .A2(n_1521), .B1(n_1563), .B2(n_1564), .Y(n_1562) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_497), .A2(n_585), .B1(n_599), .B2(n_600), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_497), .A2(n_599), .B1(n_649), .B2(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_497), .A2(n_599), .B1(n_731), .B2(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g814 ( .A(n_497), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_497), .A2(n_599), .B1(n_995), .B2(n_996), .Y(n_994) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_SL g818 ( .A(n_502), .Y(n_818) );
BUFx2_ASAP7_75t_L g980 ( .A(n_502), .Y(n_980) );
BUFx2_ASAP7_75t_L g1206 ( .A(n_502), .Y(n_1206) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g593 ( .A(n_505), .Y(n_593) );
INVx2_ASAP7_75t_L g819 ( .A(n_505), .Y(n_819) );
BUFx3_ASAP7_75t_L g981 ( .A(n_505), .Y(n_981) );
OAI31xp33_ASAP7_75t_L g515 ( .A1(n_506), .A2(n_516), .A3(n_518), .B(n_522), .Y(n_515) );
OAI31xp33_ASAP7_75t_L g978 ( .A1(n_506), .A2(n_979), .A3(n_982), .B(n_987), .Y(n_978) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g1281 ( .A1(n_507), .A2(n_1282), .B(n_1291), .Y(n_1281) );
OAI31xp33_ASAP7_75t_L g1557 ( .A1(n_507), .A2(n_1558), .A3(n_1561), .B(n_1565), .Y(n_1557) );
AND2x2_ASAP7_75t_SL g507 ( .A(n_508), .B(n_510), .Y(n_507) );
AND2x2_ASAP7_75t_L g605 ( .A(n_508), .B(n_510), .Y(n_605) );
AND2x4_ASAP7_75t_L g821 ( .A(n_508), .B(n_510), .Y(n_821) );
AND2x2_ASAP7_75t_L g890 ( .A(n_508), .B(n_510), .Y(n_890) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_508), .B(n_510), .Y(n_1120) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .C(n_539), .Y(n_514) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OAI221xp5_ASAP7_75t_L g803 ( .A1(n_527), .A2(n_755), .B1(n_771), .B2(n_804), .C(n_806), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_530), .A2(n_649), .B1(n_650), .B2(n_651), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_530), .A2(n_733), .B1(n_870), .B2(n_871), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_530), .A2(n_650), .B1(n_995), .B2(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_562), .Y(n_539) );
OAI33xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .A3(n_548), .B1(n_552), .B2(n_558), .B3(n_559), .Y(n_540) );
OAI33xp33_ASAP7_75t_L g963 ( .A1(n_541), .A2(n_558), .A3(n_964), .B1(n_966), .B2(n_968), .B3(n_970), .Y(n_963) );
OAI33xp33_ASAP7_75t_L g1021 ( .A1(n_541), .A2(n_692), .A3(n_1022), .B1(n_1024), .B2(n_1027), .B3(n_1031), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g1291 ( .A1(n_541), .A2(n_558), .B1(n_1292), .B2(n_1297), .Y(n_1291) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g964 ( .A1(n_544), .A2(n_948), .B1(n_956), .B2(n_965), .Y(n_964) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_544), .A2(n_707), .B1(n_949), .B2(n_957), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_545), .A2(n_561), .B1(n_567), .B2(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g686 ( .A(n_547), .Y(n_686) );
INVx3_ASAP7_75t_L g1585 ( .A(n_547), .Y(n_1585) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_549), .A2(n_556), .B1(n_567), .B2(n_569), .Y(n_566) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI22xp33_ASAP7_75t_SL g709 ( .A1(n_555), .A2(n_638), .B1(n_710), .B2(n_711), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_555), .A2(n_765), .B1(n_842), .B2(n_843), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g1191 ( .A1(n_555), .A2(n_919), .B1(n_1180), .B2(n_1187), .Y(n_1191) );
INVx1_ASAP7_75t_L g1224 ( .A(n_558), .Y(n_1224) );
OAI22xp5_ASAP7_75t_L g1548 ( .A1(n_564), .A2(n_1531), .B1(n_1544), .B2(n_1549), .Y(n_1548) );
OAI22xp5_ASAP7_75t_L g1556 ( .A1(n_564), .A2(n_1537), .B1(n_1540), .B2(n_1549), .Y(n_1556) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx4_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g572 ( .A(n_570), .Y(n_572) );
INVx2_ASAP7_75t_L g855 ( .A(n_570), .Y(n_855) );
INVx1_ASAP7_75t_L g1000 ( .A(n_570), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_572), .A2(n_671), .B1(n_672), .B2(n_674), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_572), .A2(n_617), .B1(n_710), .B2(n_715), .Y(n_725) );
OAI33xp33_ASAP7_75t_L g607 ( .A1(n_573), .A2(n_608), .A3(n_610), .B1(n_615), .B2(n_621), .B3(n_627), .Y(n_607) );
OAI33xp33_ASAP7_75t_L g664 ( .A1(n_573), .A2(n_665), .A3(n_669), .B1(n_670), .B2(n_675), .B3(n_678), .Y(n_664) );
OAI22xp5_ASAP7_75t_SL g794 ( .A1(n_573), .A2(n_795), .B1(n_796), .B2(n_803), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_697), .B1(n_698), .B2(n_824), .Y(n_576) );
INVx1_ASAP7_75t_L g824 ( .A(n_577), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B1(n_643), .B2(n_696), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_590), .C(n_606), .Y(n_580) );
OAI31xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .A3(n_587), .B(n_589), .Y(n_581) );
OAI31xp33_ASAP7_75t_L g645 ( .A1(n_589), .A2(n_646), .A3(n_652), .B(n_653), .Y(n_645) );
OAI31xp33_ASAP7_75t_L g998 ( .A1(n_589), .A2(n_999), .A3(n_1003), .B(n_1004), .Y(n_998) );
OAI31xp33_ASAP7_75t_SL g1043 ( .A1(n_589), .A2(n_1044), .A3(n_1049), .B(n_1051), .Y(n_1043) );
OAI31xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_594), .A3(n_601), .B(n_605), .Y(n_590) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_596), .A2(n_613), .B1(n_626), .B2(n_634), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g1055 ( .A(n_597), .B(n_1056), .C(n_1058), .Y(n_1055) );
NAND3xp33_ASAP7_75t_SL g1111 ( .A(n_597), .B(n_1112), .C(n_1116), .Y(n_1111) );
NAND3xp33_ASAP7_75t_SL g1168 ( .A(n_597), .B(n_1169), .C(n_1171), .Y(n_1168) );
INVx1_ASAP7_75t_L g813 ( .A(n_599), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_599), .A2(n_885), .B1(n_1047), .B2(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g1289 ( .A1(n_603), .A2(n_889), .B1(n_1260), .B2(n_1290), .Y(n_1289) );
OAI31xp33_ASAP7_75t_L g654 ( .A1(n_605), .A2(n_655), .A3(n_656), .B(n_662), .Y(n_654) );
OAI31xp33_ASAP7_75t_L g737 ( .A1(n_605), .A2(n_738), .A3(n_741), .B(n_744), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_632), .Y(n_606) );
INVx1_ASAP7_75t_L g1226 ( .A(n_608), .Y(n_1226) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI33xp33_ASAP7_75t_L g896 ( .A1(n_609), .A2(n_897), .A3(n_901), .B1(n_905), .B2(n_909), .B3(n_914), .Y(n_896) );
OAI33xp33_ASAP7_75t_L g1175 ( .A1(n_609), .A2(n_914), .A3(n_1176), .B1(n_1179), .B2(n_1182), .B3(n_1186), .Y(n_1175) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g724 ( .A1(n_612), .A2(n_614), .B1(n_705), .B2(n_721), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_612), .A2(n_614), .B1(n_1267), .B2(n_1268), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_614), .A2(n_628), .B1(n_630), .B2(n_631), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_614), .A2(n_628), .B1(n_711), .B2(n_716), .Y(n_727) );
OAI22xp33_ASAP7_75t_L g1007 ( .A1(n_614), .A2(n_667), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_614), .A2(n_1017), .B1(n_1019), .B2(n_1020), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_617), .A2(n_625), .B1(n_706), .B2(n_722), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_619), .A2(n_672), .B1(n_1011), .B2(n_1012), .Y(n_1010) );
INVx5_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_625), .B2(n_626), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g805 ( .A(n_623), .Y(n_805) );
OAI211xp5_ASAP7_75t_SL g1272 ( .A1(n_625), .A2(n_1273), .B(n_1274), .C(n_1277), .Y(n_1272) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx3_ASAP7_75t_L g667 ( .A(n_629), .Y(n_667) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_634), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_704) );
BUFx4f_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_SL g754 ( .A(n_636), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_638), .A2(n_671), .B1(n_679), .B2(n_688), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_638), .A2(n_674), .B1(n_680), .B2(n_691), .Y(n_690) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g839 ( .A(n_640), .Y(n_839) );
INVx1_ASAP7_75t_L g696 ( .A(n_643), .Y(n_696) );
NAND3xp33_ASAP7_75t_SL g644 ( .A(n_645), .B(n_654), .C(n_663), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g1530 ( .A1(n_657), .A2(n_1531), .B1(n_1532), .B2(n_1533), .Y(n_1530) );
INVx2_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_659), .A2(n_751), .B1(n_752), .B2(n_755), .Y(n_750) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_659), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_659), .A2(n_754), .B1(n_898), .B2(n_906), .Y(n_916) );
OAI22xp33_ASAP7_75t_L g1031 ( .A1(n_659), .A2(n_684), .B1(n_1009), .B2(n_1015), .Y(n_1031) );
OAI22xp33_ASAP7_75t_L g1063 ( .A1(n_659), .A2(n_834), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
NOR2xp33_ASAP7_75t_SL g663 ( .A(n_664), .B(n_681), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_666), .A2(n_676), .B1(n_684), .B2(n_686), .Y(n_683) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g854 ( .A(n_673), .Y(n_854) );
OAI33xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .A3(n_687), .B1(n_690), .B2(n_692), .B3(n_693), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_684), .A2(n_1008), .B1(n_1014), .B2(n_1023), .Y(n_1022) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g967 ( .A(n_689), .Y(n_967) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_745), .B1(n_822), .B2(n_823), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_700), .Y(n_822) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_728), .C(n_737), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_723), .Y(n_702) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g1536 ( .A(n_714), .Y(n_1536) );
OAI33xp33_ASAP7_75t_L g747 ( .A1(n_717), .A2(n_748), .A3(n_750), .B1(n_756), .B2(n_761), .B3(n_768), .Y(n_747) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
BUFx2_ASAP7_75t_L g1542 ( .A(n_719), .Y(n_1542) );
AOI22xp5_ASAP7_75t_L g1604 ( .A1(n_733), .A2(n_925), .B1(n_1605), .B2(n_1606), .Y(n_1604) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g823 ( .A(n_745), .Y(n_823) );
NOR4xp25_ASAP7_75t_L g746 ( .A(n_747), .B(n_772), .C(n_794), .D(n_808), .Y(n_746) );
OAI33xp33_ASAP7_75t_L g1529 ( .A1(n_748), .A2(n_1530), .A3(n_1534), .B1(n_1538), .B2(n_1541), .B3(n_1543), .Y(n_1529) );
BUFx3_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI33xp33_ASAP7_75t_L g831 ( .A1(n_749), .A2(n_832), .A3(n_836), .B1(n_841), .B2(n_844), .B3(n_847), .Y(n_831) );
OAI33xp33_ASAP7_75t_L g915 ( .A1(n_749), .A2(n_847), .A3(n_916), .B1(n_917), .B2(n_920), .B3(n_921), .Y(n_915) );
OAI33xp33_ASAP7_75t_L g1062 ( .A1(n_749), .A2(n_847), .A3(n_1063), .B1(n_1066), .B2(n_1070), .B3(n_1073), .Y(n_1062) );
OAI33xp33_ASAP7_75t_L g1189 ( .A1(n_749), .A2(n_847), .A3(n_1190), .B1(n_1191), .B2(n_1192), .B3(n_1194), .Y(n_1189) );
OAI33xp33_ASAP7_75t_L g1581 ( .A1(n_749), .A2(n_847), .A3(n_1582), .B1(n_1586), .B2(n_1589), .B3(n_1593), .Y(n_1581) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g1532 ( .A(n_753), .Y(n_1532) );
INVx2_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
OAI22xp33_ASAP7_75t_L g768 ( .A1(n_754), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B1(n_759), .B2(n_760), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g1534 ( .A1(n_760), .A2(n_1535), .B1(n_1536), .B2(n_1537), .Y(n_1534) );
OAI22xp5_ASAP7_75t_L g1538 ( .A1(n_760), .A2(n_1068), .B1(n_1539), .B2(n_1540), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_764), .B1(n_765), .B2(n_767), .Y(n_761) );
INVx2_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_SL g838 ( .A(n_763), .Y(n_838) );
INVx3_ASAP7_75t_L g1068 ( .A(n_763), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_765), .A2(n_838), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
BUFx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AOI31xp33_ASAP7_75t_SL g772 ( .A1(n_773), .A2(n_776), .A3(n_783), .B(n_793), .Y(n_772) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B1(n_789), .B2(n_790), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_784), .A2(n_789), .B1(n_818), .B2(n_819), .Y(n_817) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_786), .Y(n_807) );
INVx3_ASAP7_75t_L g1151 ( .A(n_786), .Y(n_1151) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx3_ASAP7_75t_L g799 ( .A(n_787), .Y(n_799) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_SL g1263 ( .A(n_792), .B(n_1264), .Y(n_1263) );
AO21x1_ASAP7_75t_L g1121 ( .A1(n_793), .A2(n_1122), .B(n_1126), .Y(n_1121) );
AO21x1_ASAP7_75t_L g1240 ( .A1(n_793), .A2(n_1241), .B(n_1242), .Y(n_1240) );
OAI33xp33_ASAP7_75t_L g849 ( .A1(n_795), .A2(n_850), .A3(n_853), .B1(n_856), .B2(n_857), .B3(n_860), .Y(n_849) );
OAI33xp33_ASAP7_75t_L g1076 ( .A1(n_795), .A2(n_860), .A3(n_1077), .B1(n_1079), .B2(n_1080), .B3(n_1081), .Y(n_1076) );
OAI33xp33_ASAP7_75t_L g1596 ( .A1(n_795), .A2(n_914), .A3(n_1597), .B1(n_1598), .B2(n_1599), .B3(n_1601), .Y(n_1596) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g1142 ( .A(n_799), .Y(n_1142) );
INVx1_ASAP7_75t_L g1228 ( .A(n_799), .Y(n_1228) );
INVx2_ASAP7_75t_SL g1239 ( .A(n_799), .Y(n_1239) );
INVx2_ASAP7_75t_L g1278 ( .A(n_799), .Y(n_1278) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
BUFx3_ASAP7_75t_L g1143 ( .A(n_802), .Y(n_1143) );
INVx2_ASAP7_75t_L g1153 ( .A(n_802), .Y(n_1153) );
INVx3_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AOI31xp33_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_815), .A3(n_817), .B(n_820), .Y(n_808) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_811), .Y(n_1059) );
INVx1_ASAP7_75t_L g1102 ( .A(n_811), .Y(n_1102) );
INVx2_ASAP7_75t_SL g1559 ( .A(n_816), .Y(n_1559) );
INVx1_ASAP7_75t_L g1566 ( .A(n_818), .Y(n_1566) );
INVx2_ASAP7_75t_L g1207 ( .A(n_819), .Y(n_1207) );
AO21x1_ASAP7_75t_L g1200 ( .A1(n_820), .A2(n_1201), .B(n_1204), .Y(n_1200) );
CKINVDCx14_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
OAI31xp33_ASAP7_75t_L g991 ( .A1(n_821), .A2(n_992), .A3(n_993), .B(n_997), .Y(n_991) );
INVx1_ASAP7_75t_L g1035 ( .A(n_825), .Y(n_1035) );
XOR2x1_ASAP7_75t_L g825 ( .A(n_826), .B(n_940), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_891), .B1(n_892), .B2(n_939), .Y(n_826) );
INVx1_ASAP7_75t_L g939 ( .A(n_827), .Y(n_939) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
NAND3xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_862), .C(n_876), .Y(n_829) );
NOR2xp33_ASAP7_75t_SL g830 ( .A(n_831), .B(n_849), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_833), .A2(n_845), .B1(n_851), .B2(n_852), .Y(n_850) );
OAI22xp33_ASAP7_75t_L g1194 ( .A1(n_834), .A2(n_1178), .B1(n_1185), .B2(n_1195), .Y(n_1194) );
OAI22xp5_ASAP7_75t_L g1582 ( .A1(n_834), .A2(n_1583), .B1(n_1584), .B2(n_1585), .Y(n_1582) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_835), .A2(n_846), .B1(n_854), .B2(n_855), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B1(n_839), .B2(n_840), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_837), .A2(n_842), .B1(n_854), .B2(n_855), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_839), .A2(n_1067), .B1(n_1068), .B2(n_1069), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g1589 ( .A1(n_839), .A2(n_1590), .B1(n_1591), .B2(n_1592), .Y(n_1589) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_840), .A2(n_843), .B1(n_852), .B2(n_858), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_851), .A2(n_898), .B1(n_899), .B2(n_900), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_851), .A2(n_910), .B1(n_911), .B2(n_913), .Y(n_909) );
OAI22xp33_ASAP7_75t_L g1077 ( .A1(n_851), .A2(n_1064), .B1(n_1074), .B2(n_1078), .Y(n_1077) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_851), .A2(n_911), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
OAI22xp5_ASAP7_75t_L g1186 ( .A1(n_851), .A2(n_899), .B1(n_1187), .B2(n_1188), .Y(n_1186) );
OAI22xp5_ASAP7_75t_L g1597 ( .A1(n_851), .A2(n_911), .B1(n_1583), .B2(n_1594), .Y(n_1597) );
OAI22xp5_ASAP7_75t_L g1601 ( .A1(n_851), .A2(n_852), .B1(n_1588), .B2(n_1592), .Y(n_1601) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_852), .A2(n_858), .B1(n_1069), .B2(n_1072), .Y(n_1081) );
INVx2_ASAP7_75t_L g1550 ( .A(n_852), .Y(n_1550) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_854), .A2(n_855), .B1(n_1067), .B2(n_1071), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1598 ( .A1(n_855), .A2(n_903), .B1(n_1587), .B2(n_1590), .Y(n_1598) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx2_ASAP7_75t_L g914 ( .A(n_861), .Y(n_914) );
AOI33xp33_ASAP7_75t_L g1138 ( .A1(n_861), .A2(n_1139), .A3(n_1141), .B1(n_1144), .B2(n_1148), .B3(n_1149), .Y(n_1138) );
OAI31xp33_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_872), .A3(n_874), .B(n_875), .Y(n_862) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g1133 ( .A(n_866), .Y(n_1133) );
INVx1_ASAP7_75t_L g1132 ( .A(n_867), .Y(n_1132) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
BUFx2_ASAP7_75t_L g1236 ( .A(n_868), .Y(n_1236) );
AOI32xp33_ASAP7_75t_L g879 ( .A1(n_871), .A2(n_880), .A3(n_883), .B1(n_885), .B2(n_886), .Y(n_879) );
INVx1_ASAP7_75t_L g1124 ( .A(n_873), .Y(n_1124) );
OAI31xp33_ASAP7_75t_L g922 ( .A1(n_875), .A2(n_923), .A3(n_929), .B(n_930), .Y(n_922) );
OAI31xp33_ASAP7_75t_L g1602 ( .A1(n_875), .A2(n_1603), .A3(n_1607), .B(n_1608), .Y(n_1602) );
OAI31xp33_ASAP7_75t_SL g876 ( .A1(n_877), .A2(n_878), .A3(n_887), .B(n_890), .Y(n_876) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx3_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g935 ( .A1(n_885), .A2(n_926), .B1(n_936), .B2(n_937), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_885), .A2(n_936), .B1(n_1117), .B2(n_1118), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_885), .A2(n_936), .B1(n_1163), .B2(n_1172), .Y(n_1171) );
INVxp67_ASAP7_75t_L g1287 ( .A(n_885), .Y(n_1287) );
AOI22xp33_ASAP7_75t_SL g1612 ( .A1(n_885), .A2(n_936), .B1(n_1605), .B2(n_1613), .Y(n_1612) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
OAI31xp33_ASAP7_75t_SL g932 ( .A1(n_890), .A2(n_933), .A3(n_934), .B(n_938), .Y(n_932) );
OAI31xp33_ASAP7_75t_L g1052 ( .A1(n_890), .A2(n_1053), .A3(n_1055), .B(n_1060), .Y(n_1052) );
OAI31xp33_ASAP7_75t_SL g1609 ( .A1(n_890), .A2(n_1610), .A3(n_1611), .B(n_1614), .Y(n_1609) );
INVxp67_ASAP7_75t_SL g891 ( .A(n_892), .Y(n_891) );
HB1xp67_ASAP7_75t_SL g892 ( .A(n_893), .Y(n_892) );
AND3x1_ASAP7_75t_L g894 ( .A(n_895), .B(n_922), .C(n_932), .Y(n_894) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_915), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_902), .A2(n_910), .B1(n_918), .B2(n_919), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_903), .A2(n_906), .B1(n_907), .B2(n_908), .Y(n_905) );
OAI22xp5_ASAP7_75t_L g1179 ( .A1(n_903), .A2(n_907), .B1(n_1180), .B2(n_1181), .Y(n_1179) );
OAI22xp5_ASAP7_75t_L g1182 ( .A1(n_903), .A2(n_1183), .B1(n_1184), .B2(n_1185), .Y(n_1182) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_907), .Y(n_1045) );
BUFx6f_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g1192 ( .A1(n_918), .A2(n_1181), .B1(n_1188), .B2(n_1193), .Y(n_1192) );
OAI22xp5_ASAP7_75t_L g1586 ( .A1(n_918), .A2(n_919), .B1(n_1587), .B2(n_1588), .Y(n_1586) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_925), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_924) );
INVx1_ASAP7_75t_L g1258 ( .A(n_925), .Y(n_1258) );
INVx1_ASAP7_75t_L g1286 ( .A(n_936), .Y(n_1286) );
INVx2_ASAP7_75t_SL g940 ( .A(n_941), .Y(n_940) );
OA22x2_ASAP7_75t_L g941 ( .A1(n_942), .A2(n_943), .B1(n_988), .B2(n_989), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
NAND3xp33_ASAP7_75t_L g944 ( .A(n_945), .B(n_971), .C(n_978), .Y(n_944) );
NOR2xp33_ASAP7_75t_SL g945 ( .A(n_946), .B(n_963), .Y(n_945) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
BUFx3_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVxp67_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g1023 ( .A(n_984), .Y(n_1023) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1032 ( .A(n_990), .Y(n_1032) );
NAND3xp33_ASAP7_75t_L g990 ( .A(n_991), .B(n_998), .C(n_1005), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1021), .Y(n_1005) );
INVx2_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
OAI211xp5_ASAP7_75t_L g1292 ( .A1(n_1025), .A2(n_1293), .B(n_1294), .C(n_1295), .Y(n_1292) );
INVx2_ASAP7_75t_SL g1025 ( .A(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx2_ASAP7_75t_L g1591 ( .A(n_1029), .Y(n_1591) );
INVx3_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
BUFx2_ASAP7_75t_L g1217 ( .A(n_1030), .Y(n_1217) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1030), .Y(n_1223) );
BUFx2_ASAP7_75t_L g1298 ( .A(n_1030), .Y(n_1298) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1038), .B1(n_1247), .B2(n_1248), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
XNOR2xp5_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1082), .Y(n_1039) );
INVx2_ASAP7_75t_SL g1040 ( .A(n_1041), .Y(n_1040) );
NAND3xp33_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1052), .C(n_1061), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1048), .B(n_1059), .Y(n_1058) );
NOR2xp33_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1076), .Y(n_1061) );
AOI22xp5_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1196), .B1(n_1245), .B2(n_1246), .Y(n_1082) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1083), .Y(n_1246) );
XNOR2x1_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1157), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1134), .Y(n_1084) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1086), .Y(n_1136) );
AOI21xp5_ASAP7_75t_L g1086 ( .A1(n_1087), .A2(n_1093), .B(n_1100), .Y(n_1086) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx8_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
BUFx3_ASAP7_75t_L g1105 ( .A(n_1091), .Y(n_1105) );
INVx2_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1095), .Y(n_1218) );
INVx5_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
BUFx2_ASAP7_75t_L g1296 ( .A(n_1096), .Y(n_1296) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
BUFx3_ASAP7_75t_L g1211 ( .A(n_1098), .Y(n_1211) );
OAI221xp5_ASAP7_75t_L g1101 ( .A1(n_1102), .A2(n_1103), .B1(n_1104), .B2(n_1106), .C(n_1107), .Y(n_1101) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1104), .Y(n_1214) );
INVx2_ASAP7_75t_SL g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1109), .B(n_1121), .Y(n_1135) );
OAI31xp33_ASAP7_75t_SL g1109 ( .A1(n_1110), .A2(n_1111), .A3(n_1119), .B(n_1120), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .Y(n_1112) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1118), .B(n_1131), .Y(n_1130) );
OAI31xp33_ASAP7_75t_SL g1166 ( .A1(n_1120), .A2(n_1167), .A3(n_1168), .B(n_1173), .Y(n_1166) );
NOR2xp33_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1128), .Y(n_1126) );
NAND3xp33_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1130), .C(n_1133), .Y(n_1128) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
OAI31xp33_ASAP7_75t_L g1134 ( .A1(n_1135), .A2(n_1136), .A3(n_1137), .B(n_1154), .Y(n_1134) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1138), .Y(n_1156) );
INVx2_ASAP7_75t_SL g1139 ( .A(n_1140), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_1143), .Y(n_1229) );
BUFx6f_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1156), .Y(n_1154) );
NAND3xp33_ASAP7_75t_SL g1158 ( .A(n_1159), .B(n_1166), .C(n_1174), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1164), .B(n_1170), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1189), .Y(n_1174) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1198), .Y(n_1245) );
NAND4xp25_ASAP7_75t_SL g1199 ( .A(n_1200), .B(n_1210), .C(n_1225), .D(n_1240), .Y(n_1199) );
AOI33xp33_ASAP7_75t_L g1210 ( .A1(n_1211), .A2(n_1212), .A3(n_1215), .B1(n_1219), .B2(n_1222), .B3(n_1224), .Y(n_1210) );
BUFx2_ASAP7_75t_SL g1213 ( .A(n_1214), .Y(n_1213) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
BUFx2_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx2_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
HB1xp67_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
OAI21xp5_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1279), .B(n_1281), .Y(n_1250) );
OAI21xp5_ASAP7_75t_L g1265 ( .A1(n_1266), .A2(n_1269), .B(n_1272), .Y(n_1265) );
INVx2_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
BUFx2_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
NAND2xp5_ASAP7_75t_SL g1282 ( .A(n_1283), .B(n_1289), .Y(n_1282) );
OAI221xp5_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1508), .B1(n_1512), .B2(n_1568), .C(n_1573), .Y(n_1300) );
AOI211xp5_ASAP7_75t_L g1301 ( .A1(n_1302), .A2(n_1422), .B(n_1468), .C(n_1492), .Y(n_1301) );
OAI211xp5_ASAP7_75t_L g1302 ( .A1(n_1303), .A2(n_1319), .B(n_1364), .C(n_1410), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1442 ( .A(n_1303), .B(n_1443), .Y(n_1442) );
OAI211xp5_ASAP7_75t_L g1492 ( .A1(n_1303), .A2(n_1493), .B(n_1495), .C(n_1501), .Y(n_1492) );
INVx2_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
OAI221xp5_ASAP7_75t_L g1394 ( .A1(n_1304), .A2(n_1395), .B1(n_1401), .B2(n_1404), .C(n_1406), .Y(n_1394) );
OAI32xp33_ASAP7_75t_L g1460 ( .A1(n_1304), .A2(n_1365), .A3(n_1382), .B1(n_1417), .B2(n_1461), .Y(n_1460) );
OAI221xp5_ASAP7_75t_L g1468 ( .A1(n_1304), .A2(n_1393), .B1(n_1469), .B2(n_1476), .C(n_1478), .Y(n_1468) );
INVx3_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx3_ASAP7_75t_L g1388 ( .A(n_1305), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1305), .B(n_1392), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1305), .B(n_1338), .Y(n_1405) );
OR2x2_ASAP7_75t_L g1427 ( .A(n_1305), .B(n_1360), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1305), .B(n_1351), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1305), .B(n_1376), .Y(n_1484) );
NAND2xp5_ASAP7_75t_L g1491 ( .A(n_1305), .B(n_1360), .Y(n_1491) );
NOR2xp33_ASAP7_75t_L g1496 ( .A(n_1305), .B(n_1497), .Y(n_1496) );
AND2x4_ASAP7_75t_SL g1305 ( .A(n_1306), .B(n_1313), .Y(n_1305) );
AND2x6_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1309), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1308), .B(n_1312), .Y(n_1311) );
AND2x4_ASAP7_75t_L g1314 ( .A(n_1308), .B(n_1315), .Y(n_1314) );
AND2x6_ASAP7_75t_L g1317 ( .A(n_1308), .B(n_1318), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1308), .B(n_1312), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1308), .B(n_1312), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1310), .B(n_1316), .Y(n_1315) );
HB1xp67_ASAP7_75t_L g1511 ( .A(n_1311), .Y(n_1511) );
OAI21xp5_ASAP7_75t_L g1615 ( .A1(n_1312), .A2(n_1616), .B(n_1617), .Y(n_1615) );
AOI221xp5_ASAP7_75t_L g1319 ( .A1(n_1320), .A2(n_1331), .B1(n_1342), .B2(n_1359), .C(n_1361), .Y(n_1319) );
A2O1A1Ixp33_ASAP7_75t_SL g1389 ( .A1(n_1320), .A2(n_1370), .B(n_1390), .C(n_1391), .Y(n_1389) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1320), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1327), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
OR2x2_ASAP7_75t_L g1382 ( .A(n_1322), .B(n_1327), .Y(n_1382) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1346 ( .A(n_1323), .B(n_1347), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1323), .B(n_1347), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1323), .B(n_1348), .Y(n_1373) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1323), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1397 ( .A(n_1323), .B(n_1327), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1325), .Y(n_1323) );
NOR2xp33_ASAP7_75t_L g1344 ( .A(n_1327), .B(n_1334), .Y(n_1344) );
CKINVDCx5p33_ASAP7_75t_R g1358 ( .A(n_1327), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1327), .B(n_1334), .Y(n_1363) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_1327), .B(n_1357), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1327), .B(n_1373), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1327), .B(n_1385), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1474 ( .A(n_1327), .B(n_1475), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1330), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1328), .B(n_1330), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1332), .B(n_1337), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1332), .B(n_1384), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1332), .B(n_1397), .Y(n_1396) );
OR2x2_ASAP7_75t_L g1437 ( .A(n_1332), .B(n_1400), .Y(n_1437) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1332), .B(n_1376), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1332), .B(n_1365), .Y(n_1502) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1333), .B(n_1356), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1333), .B(n_1362), .Y(n_1411) );
NOR2xp33_ASAP7_75t_L g1415 ( .A(n_1333), .B(n_1382), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1333), .B(n_1365), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1333), .B(n_1429), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1333), .B(n_1372), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_1333), .B(n_1367), .Y(n_1440) );
INVx3_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx2_ASAP7_75t_L g1370 ( .A(n_1334), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_1334), .B(n_1338), .Y(n_1455) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1334), .B(n_1367), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1336), .Y(n_1334) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1338), .Y(n_1412) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1338), .B(n_1477), .Y(n_1476) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
OR2x2_ASAP7_75t_L g1359 ( .A(n_1339), .B(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1339), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1339), .B(n_1360), .Y(n_1376) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1339), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1341), .Y(n_1339) );
OAI32xp33_ASAP7_75t_L g1342 ( .A1(n_1343), .A2(n_1345), .A3(n_1351), .B1(n_1352), .B2(n_1355), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1344), .B(n_1362), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1345), .B(n_1403), .Y(n_1402) );
NAND2xp5_ASAP7_75t_SL g1417 ( .A(n_1345), .B(n_1370), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1345), .B(n_1358), .Y(n_1459) );
OAI21xp5_ASAP7_75t_L g1464 ( .A1(n_1345), .A2(n_1465), .B(n_1467), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1345), .B(n_1363), .Y(n_1471) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1347), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1347), .B(n_1385), .Y(n_1384) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1348), .Y(n_1475) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1349), .B(n_1350), .Y(n_1348) );
OAI21xp33_ASAP7_75t_L g1413 ( .A1(n_1351), .A2(n_1414), .B(n_1416), .Y(n_1413) );
AOI221xp5_ASAP7_75t_L g1501 ( .A1(n_1351), .A2(n_1383), .B1(n_1502), .B2(n_1503), .C(n_1504), .Y(n_1501) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g1395 ( .A1(n_1352), .A2(n_1396), .B1(n_1398), .B2(n_1399), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1352), .B(n_1367), .Y(n_1398) );
CKINVDCx6p67_ASAP7_75t_R g1446 ( .A(n_1352), .Y(n_1446) );
AND2x4_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1354), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1353), .B(n_1354), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1358), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1358), .B(n_1373), .Y(n_1372) );
OR2x2_ASAP7_75t_L g1377 ( .A(n_1358), .B(n_1378), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1358), .B(n_1384), .Y(n_1383) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_1358), .B(n_1417), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1358), .B(n_1481), .Y(n_1480) );
OR2x2_ASAP7_75t_L g1387 ( .A(n_1359), .B(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1359), .Y(n_1462) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1360), .B(n_1367), .Y(n_1366) );
AOI21xp33_ASAP7_75t_L g1435 ( .A1(n_1360), .A2(n_1406), .B(n_1436), .Y(n_1435) );
NAND2xp5_ASAP7_75t_SL g1451 ( .A(n_1360), .B(n_1452), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1360), .B(n_1388), .Y(n_1507) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1361), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1494 ( .A(n_1361), .B(n_1392), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1503 ( .A(n_1361), .B(n_1393), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1363), .Y(n_1361) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1362), .Y(n_1378) );
AOI211xp5_ASAP7_75t_L g1364 ( .A1(n_1365), .A2(n_1368), .B(n_1374), .C(n_1394), .Y(n_1364) );
INVx2_ASAP7_75t_SL g1365 ( .A(n_1366), .Y(n_1365) );
NOR2xp33_ASAP7_75t_L g1449 ( .A(n_1366), .B(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1371), .Y(n_1369) );
INVx2_ASAP7_75t_L g1381 ( .A(n_1370), .Y(n_1381) );
NAND2xp5_ASAP7_75t_SL g1434 ( .A(n_1370), .B(n_1398), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1370), .B(n_1454), .Y(n_1488) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1373), .Y(n_1483) );
OAI211xp5_ASAP7_75t_L g1374 ( .A1(n_1375), .A2(n_1377), .B(n_1379), .C(n_1389), .Y(n_1374) );
CKINVDCx14_ASAP7_75t_R g1375 ( .A(n_1376), .Y(n_1375) );
NOR2xp33_ASAP7_75t_L g1424 ( .A(n_1377), .B(n_1387), .Y(n_1424) );
OR2x2_ASAP7_75t_L g1466 ( .A(n_1378), .B(n_1403), .Y(n_1466) );
OAI21xp5_ASAP7_75t_L g1379 ( .A1(n_1380), .A2(n_1383), .B(n_1386), .Y(n_1379) );
NOR2xp33_ASAP7_75t_L g1380 ( .A(n_1381), .B(n_1382), .Y(n_1380) );
AOI311xp33_ASAP7_75t_L g1456 ( .A1(n_1381), .A2(n_1426), .A3(n_1457), .B(n_1460), .C(n_1463), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1381), .B(n_1383), .Y(n_1490) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1383), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1384), .B(n_1403), .Y(n_1429) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1384), .Y(n_1482) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1388), .B(n_1462), .Y(n_1461) );
AOI221xp5_ASAP7_75t_L g1430 ( .A1(n_1391), .A2(n_1431), .B1(n_1433), .B2(n_1442), .C(n_1444), .Y(n_1430) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1392), .Y(n_1418) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
AOI21xp5_ASAP7_75t_L g1504 ( .A1(n_1401), .A2(n_1505), .B(n_1506), .Y(n_1504) );
CKINVDCx5p33_ASAP7_75t_R g1401 ( .A(n_1402), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1403), .B(n_1411), .Y(n_1479) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1406), .Y(n_1443) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1408), .B(n_1409), .Y(n_1407) );
AOI221xp5_ASAP7_75t_L g1410 ( .A1(n_1411), .A2(n_1412), .B1(n_1413), .B2(n_1418), .C(n_1419), .Y(n_1410) );
INVxp33_ASAP7_75t_SL g1414 ( .A(n_1415), .Y(n_1414) );
OAI31xp33_ASAP7_75t_L g1486 ( .A1(n_1418), .A2(n_1436), .A3(n_1465), .B(n_1487), .Y(n_1486) );
NOR2xp33_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1421), .Y(n_1419) );
OAI211xp5_ASAP7_75t_L g1433 ( .A1(n_1420), .A2(n_1434), .B(n_1435), .C(n_1438), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1420), .B(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1421), .Y(n_1498) );
NAND3xp33_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1430), .C(n_1456), .Y(n_1422) );
NOR2xp33_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1425), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1428), .Y(n_1425) );
AOI22xp33_ASAP7_75t_SL g1469 ( .A1(n_1426), .A2(n_1470), .B1(n_1472), .B2(n_1473), .Y(n_1469) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1429), .Y(n_1500) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_1439), .B(n_1441), .Y(n_1438) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
OAI211xp5_ASAP7_75t_L g1444 ( .A1(n_1445), .A2(n_1447), .B(n_1448), .C(n_1451), .Y(n_1444) );
CKINVDCx6p67_ASAP7_75t_R g1445 ( .A(n_1446), .Y(n_1445) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVxp33_ASAP7_75t_SL g1505 ( .A(n_1452), .Y(n_1505) );
NOR2xp33_ASAP7_75t_L g1452 ( .A(n_1453), .B(n_1455), .Y(n_1452) );
CKINVDCx14_ASAP7_75t_R g1453 ( .A(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVxp67_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1466), .B(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
O2A1O1Ixp33_ASAP7_75t_L g1478 ( .A1(n_1479), .A2(n_1480), .B(n_1484), .C(n_1485), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1481 ( .A(n_1482), .B(n_1483), .Y(n_1481) );
AOI21xp5_ASAP7_75t_L g1485 ( .A1(n_1486), .A2(n_1489), .B(n_1491), .Y(n_1485) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
OAI21xp33_ASAP7_75t_L g1495 ( .A1(n_1496), .A2(n_1498), .B(n_1499), .Y(n_1495) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
CKINVDCx20_ASAP7_75t_R g1508 ( .A(n_1509), .Y(n_1508) );
CKINVDCx20_ASAP7_75t_R g1509 ( .A(n_1510), .Y(n_1509) );
INVx4_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
HB1xp67_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
NAND3xp33_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1528), .C(n_1557), .Y(n_1517) );
NOR2xp33_ASAP7_75t_SL g1528 ( .A(n_1529), .B(n_1546), .Y(n_1528) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
OAI33xp33_ASAP7_75t_L g1546 ( .A1(n_1547), .A2(n_1548), .A3(n_1551), .B1(n_1552), .B2(n_1553), .B3(n_1556), .Y(n_1546) );
INVx2_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
INVx2_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVx2_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
BUFx3_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
BUFx3_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVxp33_ASAP7_75t_SL g1576 ( .A(n_1577), .Y(n_1576) );
HB1xp67_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
AND3x1_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1602), .C(n_1609), .Y(n_1579) );
NOR2xp33_ASAP7_75t_SL g1580 ( .A(n_1581), .B(n_1596), .Y(n_1580) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
endmodule