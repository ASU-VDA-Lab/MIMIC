module fake_jpeg_7802_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_0),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

CKINVDCx10_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_56),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_65),
.Y(n_69)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_45),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_46),
.B1(n_48),
.B2(n_53),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_67),
.A2(n_83),
.B1(n_86),
.B2(n_16),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_47),
.B(n_49),
.C(n_55),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_50),
.B1(n_43),
.B2(n_52),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_75),
.B1(n_17),
.B2(n_19),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_23),
.B1(n_37),
.B2(n_36),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_1),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_2),
.B1(n_3),
.B2(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_2),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_3),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_92),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_25),
.CON(n_102),
.SN(n_102)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_80),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_101),
.C(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_103),
.C(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_112),
.B(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_99),
.B(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_116),
.B(n_93),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_102),
.C(n_94),
.Y(n_118)
);

OAI221xp5_ASAP7_75t_SL g119 ( 
.A1(n_118),
.A2(n_100),
.B1(n_106),
.B2(n_96),
.C(n_29),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_104),
.B(n_95),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_69),
.Y(n_121)
);


endmodule