module real_jpeg_26945_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

INVx11_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_65),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_1),
.A2(n_25),
.B1(n_30),
.B2(n_65),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_65),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_68),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_2),
.A2(n_25),
.B1(n_30),
.B2(n_68),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_4),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_78),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_4),
.A2(n_25),
.B1(n_30),
.B2(n_78),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_6),
.A2(n_25),
.B1(n_30),
.B2(n_48),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_6),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_113)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_7),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_7),
.A2(n_57),
.B(n_58),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_143),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_7),
.B(n_38),
.Y(n_204)
);

A2O1A1O1Ixp25_ASAP7_75t_L g206 ( 
.A1(n_7),
.A2(n_38),
.B(n_42),
.C(n_204),
.D(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_7),
.B(n_72),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_7),
.A2(n_24),
.B(n_217),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g244 ( 
.A1(n_7),
.A2(n_59),
.B(n_71),
.C(n_156),
.D(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_7),
.B(n_59),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_9),
.A2(n_25),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_9),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_10),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_99),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_99),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_10),
.A2(n_25),
.B1(n_30),
.B2(n_99),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_11),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_11),
.A2(n_25),
.B1(n_30),
.B2(n_40),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_12),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_12),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_86)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_13),
.A2(n_25),
.B1(n_30),
.B2(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_13),
.B(n_25),
.Y(n_205)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_20),
.B(n_105),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.C(n_90),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_21),
.B(n_82),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_50),
.B1(n_51),
.B2(n_81),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_36),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_24),
.A2(n_34),
.B(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_24),
.A2(n_28),
.B1(n_29),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_24),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_24),
.A2(n_89),
.B1(n_149),
.B2(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_24),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_24),
.B(n_219),
.Y(n_232)
);

NAND2x1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_28),
.B(n_143),
.Y(n_236)
);

AOI32xp33_ASAP7_75t_L g203 ( 
.A1(n_30),
.A2(n_39),
.A3(n_44),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_30),
.B(n_236),
.Y(n_235)
);

INVx5_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_33),
.B(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_33),
.A2(n_232),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_37),
.A2(n_41),
.B1(n_49),
.B2(n_96),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_43),
.Y(n_45)
);

AOI32xp33_ASAP7_75t_L g252 ( 
.A1(n_38),
.A2(n_58),
.A3(n_245),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_39),
.B(n_76),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_41),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_42),
.A2(n_46),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_42),
.A2(n_46),
.B1(n_86),
.B2(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_42),
.B(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_42),
.A2(n_46),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_49),
.A2(n_96),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_49),
.B(n_172),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_49),
.A2(n_170),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_49),
.B(n_143),
.Y(n_229)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_69),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_52),
.B(n_69),
.C(n_81),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_63),
.B(n_66),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_54),
.A2(n_55),
.B1(n_64),
.B2(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_54),
.B(n_67),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_54),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_60),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_56),
.A2(n_61),
.B(n_143),
.C(n_144),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_59),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_66),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_70),
.A2(n_153),
.B(n_155),
.Y(n_152)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_72),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_71),
.A2(n_72),
.B1(n_154),
.B2(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_76),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_79),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_79),
.B(n_104),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_79),
.A2(n_102),
.B(n_178),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_80),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_88),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_88),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_89),
.A2(n_224),
.B(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_90),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.C(n_100),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_92),
.B(n_95),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_94),
.A2(n_147),
.B1(n_148),
.B2(n_150),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_133),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_98),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_125),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_115),
.B1(n_116),
.B2(n_124),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B(n_114),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_111),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_122),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_122),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_120),
.B(n_143),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_159),
.B(n_274),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_157),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_130),
.B(n_157),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.C(n_135),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_131),
.B(n_134),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_135),
.A2(n_136),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_151),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_138),
.B1(n_151),
.B2(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_147),
.A2(n_150),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_196),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_182),
.B(n_195),
.Y(n_161)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_162),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_179),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_179),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.C(n_176),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_169),
.B1(n_176),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_183),
.B(n_185),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_190),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_186),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_189),
.B(n_190),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.C(n_194),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_191),
.B(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_192),
.B(n_194),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_193),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_272),
.C(n_273),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_267),
.B(n_271),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_256),
.B(n_266),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_240),
.B(n_255),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_220),
.B(n_239),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_202),
.B(n_208),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_206),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_213),
.C(n_215),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_214),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_216),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_227),
.B(n_238),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_226),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_233),
.B(n_237),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_241),
.B(n_242),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_249),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_246),
.C(n_249),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_248),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_252),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_262),
.C(n_263),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);


endmodule