module fake_netlist_1_667_n_654 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_654);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_654;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_476;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_163;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_24), .Y(n_75) );
BUFx5_ASAP7_75t_L g76 ( .A(n_54), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_62), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_41), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_30), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_44), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_29), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_2), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_20), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_49), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_46), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_9), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_36), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_69), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_45), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_12), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_47), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_52), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_13), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_43), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_42), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_34), .Y(n_97) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_28), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_1), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_4), .Y(n_100) );
INVx3_ASAP7_75t_L g101 ( .A(n_6), .Y(n_101) );
INVx3_ASAP7_75t_L g102 ( .A(n_19), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_1), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_51), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_31), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_38), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_64), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_59), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_4), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_11), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_68), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_3), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_37), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_2), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_40), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_76), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_101), .B(n_0), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_106), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_98), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_90), .B(n_3), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_101), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_101), .B(n_5), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_102), .B(n_5), .Y(n_128) );
NOR2xp33_ASAP7_75t_SL g129 ( .A(n_87), .B(n_27), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_98), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_102), .Y(n_131) );
INVxp33_ASAP7_75t_SL g132 ( .A(n_116), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_76), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_102), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_75), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_76), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_75), .Y(n_137) );
INVxp67_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_82), .B(n_6), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_83), .B(n_7), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_83), .B(n_7), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_77), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_94), .B(n_8), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_76), .B(n_8), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_77), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_76), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_78), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_76), .Y(n_148) );
NOR2x1_ASAP7_75t_L g149 ( .A(n_96), .B(n_10), .Y(n_149) );
INVxp67_ASAP7_75t_L g150 ( .A(n_94), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_76), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_98), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_78), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_80), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_80), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_81), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_105), .B(n_10), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_81), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_84), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_76), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_124), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_121), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_122), .B(n_112), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_123), .B(n_104), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_121), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_121), .Y(n_167) );
NAND3x1_ASAP7_75t_L g168 ( .A(n_149), .B(n_117), .C(n_111), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_133), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_123), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_122), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_133), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_122), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_122), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_138), .B(n_120), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_127), .B(n_117), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_136), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_124), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_138), .B(n_108), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_148), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_151), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_127), .B(n_114), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_127), .B(n_114), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_150), .B(n_79), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_150), .B(n_109), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_126), .B(n_110), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_125), .B(n_111), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_139), .A2(n_113), .B1(n_99), .B2(n_103), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_125), .B(n_113), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_127), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_128), .B(n_119), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_135), .B(n_79), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_126), .B(n_89), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_151), .Y(n_203) );
AND2x6_ASAP7_75t_L g204 ( .A(n_139), .B(n_118), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_151), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_139), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_131), .B(n_89), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_139), .B(n_100), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_135), .B(n_86), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_140), .B(n_85), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_140), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_161), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_124), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_137), .B(n_118), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_153), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_140), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_170), .B(n_140), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_204), .A2(n_141), .B1(n_143), .B2(n_145), .Y(n_221) );
INVx3_ASAP7_75t_SL g222 ( .A(n_200), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_204), .B(n_153), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_204), .B(n_153), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_174), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_198), .B(n_141), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_174), .Y(n_227) );
AND2x6_ASAP7_75t_L g228 ( .A(n_199), .B(n_141), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_171), .A2(n_144), .B(n_159), .Y(n_229) );
OR2x2_ASAP7_75t_SL g230 ( .A(n_172), .B(n_128), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_170), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_178), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_206), .A2(n_129), .B1(n_141), .B2(n_143), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_178), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_178), .Y(n_235) );
AOI221xp5_ASAP7_75t_SL g236 ( .A1(n_197), .A2(n_160), .B1(n_159), .B2(n_137), .C(n_142), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_178), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_204), .B(n_158), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_165), .B(n_160), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_171), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_191), .Y(n_241) );
OR2x6_ASAP7_75t_L g242 ( .A(n_196), .B(n_149), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_200), .B(n_142), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_206), .A2(n_154), .B1(n_145), .B2(n_156), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_191), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_204), .B(n_158), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_212), .B(n_129), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_191), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_191), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_164), .Y(n_250) );
AOI21xp33_ASAP7_75t_L g251 ( .A1(n_166), .A2(n_156), .B(n_155), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_212), .B(n_155), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_204), .B(n_158), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_204), .B(n_158), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_164), .B(n_154), .Y(n_255) );
CKINVDCx11_ASAP7_75t_R g256 ( .A(n_192), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_192), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_196), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_212), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_198), .B(n_147), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_209), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_193), .B(n_147), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_164), .B(n_134), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_164), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_192), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_164), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_192), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_164), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_217), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_164), .B(n_134), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_217), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_171), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_209), .B(n_131), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_208), .B(n_157), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_171), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_211), .A2(n_97), .B1(n_95), .B2(n_85), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_211), .Y(n_277) );
AOI21x1_ASAP7_75t_L g278 ( .A1(n_218), .A2(n_88), .B(n_91), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_208), .B(n_88), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_218), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_269), .Y(n_281) );
AOI221xp5_ASAP7_75t_L g282 ( .A1(n_258), .A2(n_195), .B1(n_186), .B2(n_177), .C(n_194), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_271), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_250), .B(n_226), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_264), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_240), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_280), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_243), .B(n_208), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_264), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_236), .B(n_207), .C(n_202), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_222), .B(n_201), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_230), .B(n_208), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_277), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_272), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_231), .Y(n_295) );
OR2x6_ASAP7_75t_L g296 ( .A(n_264), .B(n_211), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_275), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_221), .A2(n_211), .B1(n_212), .B2(n_219), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_250), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_232), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_234), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_259), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_235), .Y(n_303) );
OR2x6_ASAP7_75t_L g304 ( .A(n_266), .B(n_219), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_250), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_260), .B(n_219), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_237), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_277), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_277), .Y(n_309) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_278), .A2(n_93), .B(n_92), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_250), .B(n_219), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_220), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_256), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_225), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_241), .Y(n_315) );
AOI222xp33_ASAP7_75t_L g316 ( .A1(n_261), .A2(n_216), .B1(n_176), .B2(n_93), .C1(n_91), .C2(n_92), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_220), .Y(n_317) );
NOR2xp33_ASAP7_75t_SL g318 ( .A(n_268), .B(n_176), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_225), .Y(n_319) );
INVx1_ASAP7_75t_SL g320 ( .A(n_260), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_225), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_226), .B(n_176), .Y(n_322) );
AOI21xp33_ASAP7_75t_L g323 ( .A1(n_244), .A2(n_176), .B(n_168), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_259), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_244), .Y(n_325) );
INVx4_ASAP7_75t_L g326 ( .A(n_228), .Y(n_326) );
NAND2x1_ASAP7_75t_SL g327 ( .A(n_233), .B(n_112), .Y(n_327) );
CKINVDCx6p67_ASAP7_75t_R g328 ( .A(n_313), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_281), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_325), .A2(n_274), .B1(n_242), .B2(n_249), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_292), .A2(n_274), .B1(n_242), .B2(n_248), .Y(n_331) );
OAI22xp5_ASAP7_75t_SL g332 ( .A1(n_295), .A2(n_242), .B1(n_276), .B2(n_239), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_281), .Y(n_333) );
INVx6_ASAP7_75t_L g334 ( .A(n_284), .Y(n_334) );
OR2x6_ASAP7_75t_L g335 ( .A(n_296), .B(n_279), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_320), .A2(n_265), .B1(n_257), .B2(n_245), .Y(n_336) );
AOI22xp33_ASAP7_75t_SL g337 ( .A1(n_312), .A2(n_279), .B1(n_228), .B2(n_268), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_291), .B(n_273), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_291), .Y(n_339) );
AOI22xp33_ASAP7_75t_SL g340 ( .A1(n_317), .A2(n_228), .B1(n_273), .B2(n_262), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_283), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_306), .B(n_267), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_283), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_287), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_322), .A2(n_228), .B1(n_227), .B2(n_255), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_287), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_319), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_288), .A2(n_247), .B(n_252), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_296), .A2(n_255), .B1(n_223), .B2(n_246), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_296), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_300), .Y(n_351) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_296), .A2(n_246), .B1(n_223), .B2(n_254), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_300), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_306), .A2(n_270), .B1(n_263), .B2(n_254), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_296), .A2(n_238), .B1(n_224), .B2(n_253), .Y(n_355) );
AO21x2_ASAP7_75t_L g356 ( .A1(n_310), .A2(n_251), .B(n_229), .Y(n_356) );
AO31x2_ASAP7_75t_L g357 ( .A1(n_326), .A2(n_115), .A3(n_107), .B(n_238), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_335), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_333), .A2(n_290), .B1(n_326), .B2(n_323), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_332), .A2(n_282), .B1(n_290), .B2(n_322), .C(n_303), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_335), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_333), .A2(n_326), .B1(n_298), .B2(n_301), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_346), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_348), .A2(n_318), .B(n_310), .Y(n_364) );
OAI221xp5_ASAP7_75t_L g365 ( .A1(n_330), .A2(n_327), .B1(n_316), .B2(n_301), .C(n_303), .Y(n_365) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_331), .A2(n_327), .B(n_251), .C(n_307), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_338), .A2(n_322), .B1(n_284), .B2(n_326), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_335), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_340), .A2(n_322), .B1(n_284), .B2(n_309), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_335), .A2(n_168), .B1(n_315), .B2(n_307), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_346), .B(n_315), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_329), .A2(n_263), .B(n_270), .C(n_253), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_329), .B(n_284), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_343), .A2(n_309), .B1(n_324), .B2(n_308), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_343), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_344), .B(n_294), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_344), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_341), .B(n_294), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_350), .A2(n_324), .B1(n_293), .B2(n_308), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_351), .B(n_297), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g382 ( .A1(n_336), .A2(n_115), .B(n_308), .C(n_293), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g383 ( .A1(n_328), .A2(n_304), .B1(n_224), .B2(n_297), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_371), .A2(n_328), .B1(n_350), .B2(n_351), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_369), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_364), .A2(n_356), .B(n_310), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_363), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_363), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_376), .B(n_353), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_376), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g391 ( .A1(n_360), .A2(n_337), .B1(n_345), .B2(n_342), .C(n_354), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_377), .B(n_357), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_377), .B(n_357), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_365), .A2(n_352), .B1(n_334), .B2(n_347), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_365), .A2(n_334), .B1(n_347), .B2(n_304), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_363), .B(n_357), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_372), .B(n_357), .Y(n_397) );
NAND3xp33_ASAP7_75t_L g398 ( .A(n_366), .B(n_98), .C(n_152), .Y(n_398) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_383), .A2(n_342), .B(n_355), .C(n_349), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_371), .A2(n_334), .B1(n_324), .B2(n_293), .C(n_308), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
CKINVDCx11_ASAP7_75t_R g402 ( .A(n_361), .Y(n_402) );
OAI222xp33_ASAP7_75t_L g403 ( .A1(n_361), .A2(n_107), .B1(n_304), .B2(n_286), .C1(n_357), .C2(n_293), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_368), .A2(n_334), .B1(n_314), .B2(n_319), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_378), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_358), .B(n_314), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_368), .A2(n_304), .B1(n_314), .B2(n_286), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_374), .A2(n_356), .B1(n_324), .B2(n_302), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_372), .B(n_356), .Y(n_409) );
AND2x4_ASAP7_75t_SL g410 ( .A(n_374), .B(n_314), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_374), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_378), .B(n_314), .Y(n_412) );
NAND4xp25_ASAP7_75t_SL g413 ( .A(n_370), .B(n_11), .C(n_12), .D(n_13), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_381), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_379), .B(n_321), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_358), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_381), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_413), .A2(n_359), .B(n_362), .Y(n_418) );
OAI33xp33_ASAP7_75t_L g419 ( .A1(n_384), .A2(n_359), .A3(n_362), .B1(n_16), .B2(n_17), .B3(n_18), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_409), .B(n_374), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_385), .A2(n_358), .B1(n_367), .B2(n_375), .C(n_373), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_409), .B(n_358), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_405), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_405), .Y(n_424) );
CKINVDCx14_ASAP7_75t_R g425 ( .A(n_402), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_401), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_405), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_392), .B(n_382), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_390), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_414), .B(n_380), .Y(n_431) );
NOR2xp67_ASAP7_75t_L g432 ( .A(n_398), .B(n_21), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_392), .B(n_98), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_393), .B(n_14), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_415), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_398), .A2(n_285), .B(n_304), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_388), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_387), .B(n_50), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_414), .B(n_14), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_417), .B(n_15), .Y(n_440) );
AO22x1_ASAP7_75t_L g441 ( .A1(n_395), .A2(n_289), .B1(n_299), .B2(n_311), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_393), .B(n_15), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_397), .B(n_16), .Y(n_443) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_408), .B(n_152), .C(n_124), .Y(n_444) );
INVx4_ASAP7_75t_L g445 ( .A(n_410), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_390), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_387), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_396), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_397), .B(n_17), .Y(n_449) );
OAI332xp33_ASAP7_75t_L g450 ( .A1(n_394), .A2(n_18), .A3(n_19), .B1(n_20), .B2(n_302), .B3(n_215), .C1(n_210), .C2(n_190), .Y(n_450) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_386), .A2(n_166), .B(n_215), .Y(n_451) );
NAND4xp25_ASAP7_75t_L g452 ( .A(n_395), .B(n_311), .C(n_188), .D(n_184), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_396), .B(n_152), .Y(n_453) );
OAI211xp5_ASAP7_75t_L g454 ( .A1(n_399), .A2(n_130), .B(n_124), .C(n_152), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_388), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_412), .B(n_152), .Y(n_457) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_388), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_412), .B(n_152), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_388), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_399), .B(n_311), .C(n_188), .D(n_184), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g462 ( .A1(n_394), .A2(n_124), .B(n_130), .C(n_311), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_417), .B(n_130), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_407), .A2(n_285), .B(n_289), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_391), .A2(n_130), .B1(n_175), .B2(n_179), .C(n_180), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_427), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_422), .B(n_388), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_435), .B(n_389), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_422), .B(n_388), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_430), .Y(n_470) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_434), .B(n_416), .Y(n_471) );
NAND4xp25_ASAP7_75t_L g472 ( .A(n_434), .B(n_416), .C(n_411), .D(n_400), .Y(n_472) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_456), .Y(n_473) );
OAI221xp5_ASAP7_75t_L g474 ( .A1(n_461), .A2(n_411), .B1(n_404), .B2(n_130), .C(n_299), .Y(n_474) );
OAI322xp33_ASAP7_75t_L g475 ( .A1(n_425), .A2(n_130), .A3(n_411), .B1(n_214), .B2(n_162), .C1(n_183), .C2(n_403), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_443), .B(n_411), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_443), .B(n_406), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_430), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_448), .B(n_406), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_449), .B(n_406), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_448), .B(n_406), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_449), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_420), .B(n_410), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g484 ( .A(n_450), .B(n_169), .C(n_175), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_446), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_446), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_420), .B(n_410), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_433), .B(n_22), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_433), .B(n_23), .Y(n_490) );
NAND4xp25_ASAP7_75t_L g491 ( .A(n_462), .B(n_169), .C(n_179), .D(n_210), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_423), .B(n_25), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_424), .Y(n_493) );
NAND2x1p5_ASAP7_75t_L g494 ( .A(n_445), .B(n_285), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_424), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_442), .B(n_26), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_428), .Y(n_497) );
NAND2xp33_ASAP7_75t_L g498 ( .A(n_442), .B(n_285), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_428), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_453), .B(n_32), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_453), .B(n_33), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g502 ( .A(n_419), .B(n_180), .C(n_189), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g503 ( .A1(n_439), .A2(n_35), .B(n_39), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_431), .B(n_48), .Y(n_504) );
AO211x2_ASAP7_75t_L g505 ( .A1(n_452), .A2(n_53), .B(n_55), .C(n_56), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_426), .B(n_57), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_426), .B(n_58), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_447), .B(n_60), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_454), .A2(n_189), .B(n_190), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_447), .B(n_61), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_460), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_463), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_440), .B(n_63), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_462), .A2(n_182), .B(n_213), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_437), .B(n_455), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_429), .Y(n_516) );
AOI33xp33_ASAP7_75t_L g517 ( .A1(n_421), .A2(n_182), .A3(n_213), .B1(n_205), .B2(n_203), .B3(n_187), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_429), .B(n_65), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_437), .B(n_66), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_457), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_516), .B(n_418), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_466), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_473), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_472), .B(n_441), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_470), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_478), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_479), .B(n_445), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_468), .B(n_457), .Y(n_528) );
NAND4xp25_ASAP7_75t_L g529 ( .A(n_482), .B(n_465), .C(n_436), .D(n_445), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_485), .B(n_459), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_477), .B(n_455), .Y(n_531) );
AOI211xp5_ASAP7_75t_L g532 ( .A1(n_474), .A2(n_441), .B(n_432), .C(n_459), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_486), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_487), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_493), .Y(n_535) );
NOR3xp33_ASAP7_75t_L g536 ( .A(n_475), .B(n_444), .C(n_432), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_467), .B(n_460), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_495), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_483), .B(n_458), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_497), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_499), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_480), .B(n_451), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_493), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_481), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_467), .B(n_451), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_476), .B(n_451), .Y(n_546) );
BUFx3_ASAP7_75t_L g547 ( .A(n_494), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_481), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_515), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_471), .B(n_438), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_498), .A2(n_438), .B(n_464), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_483), .Y(n_552) );
NAND4xp25_ASAP7_75t_L g553 ( .A(n_518), .B(n_438), .C(n_185), .D(n_187), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_511), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_488), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_469), .B(n_438), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_512), .B(n_72), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_471), .B(n_520), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_515), .Y(n_559) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_491), .B(n_173), .C(n_205), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_518), .B(n_73), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_488), .B(n_162), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_469), .B(n_162), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_511), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_517), .B(n_162), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_498), .A2(n_285), .B(n_305), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_517), .B(n_162), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_492), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_524), .A2(n_505), .B1(n_513), .B2(n_496), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_524), .B(n_494), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_521), .B(n_484), .C(n_490), .D(n_489), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_523), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_552), .B(n_519), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_555), .B(n_519), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_525), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_529), .A2(n_505), .B1(n_489), .B2(n_490), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_549), .B(n_500), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_526), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_553), .A2(n_522), .B1(n_545), .B2(n_561), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_533), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_534), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_543), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_538), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_540), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_544), .B(n_501), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_549), .B(n_501), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_554), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_541), .Y(n_588) );
XOR2x2_ASAP7_75t_L g589 ( .A(n_561), .B(n_500), .Y(n_589) );
XOR2x2_ASAP7_75t_L g590 ( .A(n_527), .B(n_502), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_548), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_559), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_531), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_528), .B(n_510), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_545), .B(n_507), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_558), .B(n_504), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_535), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_542), .B(n_506), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_535), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_568), .A2(n_503), .B1(n_506), .B2(n_514), .C(n_508), .Y(n_600) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_536), .A2(n_509), .B(n_510), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_562), .B(n_508), .C(n_167), .Y(n_602) );
AOI322xp5_ASAP7_75t_L g603 ( .A1(n_527), .A2(n_183), .A3(n_214), .B1(n_305), .B2(n_181), .C1(n_173), .C2(n_185), .Y(n_603) );
OAI211xp5_ASAP7_75t_SL g604 ( .A1(n_532), .A2(n_163), .B(n_167), .C(n_181), .Y(n_604) );
OAI21xp33_ASAP7_75t_L g605 ( .A1(n_546), .A2(n_183), .B(n_214), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_537), .B(n_183), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_530), .A2(n_554), .B1(n_537), .B2(n_539), .C(n_527), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_564), .B(n_183), .Y(n_608) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_547), .A2(n_305), .B(n_214), .C(n_203), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_550), .A2(n_305), .B1(n_214), .B2(n_163), .Y(n_610) );
INVxp67_ASAP7_75t_SL g611 ( .A(n_554), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_556), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_556), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_547), .B(n_563), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_551), .B(n_557), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_567), .Y(n_616) );
AOI21xp33_ASAP7_75t_L g617 ( .A1(n_565), .A2(n_566), .B(n_536), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_560), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_560), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_521), .B(n_516), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_522), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_583), .Y(n_622) );
NAND4xp25_ASAP7_75t_SL g623 ( .A(n_607), .B(n_579), .C(n_576), .D(n_569), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_570), .A2(n_571), .B1(n_621), .B2(n_611), .Y(n_624) );
OAI211xp5_ASAP7_75t_SL g625 ( .A1(n_576), .A2(n_570), .B(n_617), .C(n_616), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_617), .A2(n_604), .B(n_596), .C(n_615), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_572), .Y(n_627) );
NAND3x1_ASAP7_75t_L g628 ( .A(n_602), .B(n_601), .C(n_596), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_590), .A2(n_593), .B1(n_618), .B2(n_619), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_590), .A2(n_589), .B1(n_620), .B2(n_577), .Y(n_630) );
AOI211xp5_ASAP7_75t_L g631 ( .A1(n_600), .A2(n_610), .B(n_587), .C(n_614), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_589), .A2(n_586), .B1(n_591), .B2(n_573), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_588), .Y(n_633) );
XOR2xp5_ASAP7_75t_L g634 ( .A(n_614), .B(n_594), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_630), .A2(n_582), .B1(n_587), .B2(n_578), .Y(n_635) );
AO21x1_ASAP7_75t_L g636 ( .A1(n_624), .A2(n_610), .B(n_575), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_622), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g638 ( .A1(n_623), .A2(n_605), .B(n_582), .C(n_609), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_629), .B(n_613), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_626), .B(n_592), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_632), .A2(n_612), .B1(n_585), .B2(n_595), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_637), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_639), .B(n_627), .Y(n_643) );
NAND5xp2_ASAP7_75t_L g644 ( .A(n_638), .B(n_631), .C(n_628), .D(n_603), .E(n_625), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_640), .B(n_633), .Y(n_645) );
NAND4xp25_ASAP7_75t_L g646 ( .A(n_644), .B(n_635), .C(n_636), .D(n_606), .Y(n_646) );
OR4x2_ASAP7_75t_L g647 ( .A(n_643), .B(n_635), .C(n_634), .D(n_641), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_643), .B(n_580), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_648), .B(n_645), .Y(n_649) );
OA21x2_ASAP7_75t_L g650 ( .A1(n_646), .A2(n_642), .B(n_608), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_650), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_649), .B1(n_647), .B2(n_581), .Y(n_652) );
XNOR2xp5_ASAP7_75t_L g653 ( .A(n_652), .B(n_584), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_597), .B1(n_599), .B2(n_574), .C(n_598), .Y(n_654) );
endmodule