module real_aes_6810_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_404;
wire n_147;
wire n_288;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp5_ASAP7_75t_SL g445 ( .A1(n_0), .A2(n_68), .B1(n_446), .B2(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g140 ( .A(n_1), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_2), .A2(n_34), .B1(n_106), .B2(n_158), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_3), .B(n_109), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_4), .Y(n_460) );
AND2x6_ASAP7_75t_L g111 ( .A(n_5), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g498 ( .A(n_5), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_5), .B(n_504), .Y(n_503) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_6), .Y(n_402) );
AO22x2_ASAP7_75t_L g420 ( .A1(n_7), .A2(n_30), .B1(n_421), .B2(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g132 ( .A(n_8), .Y(n_132) );
INVx1_ASAP7_75t_L g93 ( .A(n_9), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_10), .B(n_99), .Y(n_152) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_11), .A2(n_60), .B1(n_474), .B2(n_477), .Y(n_473) );
XOR2xp5_ASAP7_75t_L g512 ( .A(n_12), .B(n_410), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g88 ( .A(n_13), .B(n_89), .Y(n_88) );
AO32x2_ASAP7_75t_L g169 ( .A1(n_14), .A2(n_109), .A3(n_110), .B1(n_129), .B2(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_15), .B(n_106), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_16), .A2(n_398), .B1(n_405), .B2(n_406), .Y(n_397) );
INVx1_ASAP7_75t_L g405 ( .A(n_16), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_17), .B(n_89), .Y(n_142) );
AO22x2_ASAP7_75t_L g424 ( .A1(n_18), .A2(n_33), .B1(n_421), .B2(n_425), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_19), .A2(n_42), .B1(n_106), .B2(n_158), .Y(n_172) );
AOI22xp33_ASAP7_75t_SL g166 ( .A1(n_20), .A2(n_63), .B1(n_99), .B2(n_106), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_21), .B(n_106), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_22), .A2(n_48), .B1(n_453), .B2(n_455), .Y(n_452) );
BUFx6f_ASAP7_75t_L g97 ( .A(n_23), .Y(n_97) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_24), .B(n_148), .Y(n_206) );
AOI22xp5_ASAP7_75t_SL g437 ( .A1(n_25), .A2(n_47), .B1(n_438), .B2(n_442), .Y(n_437) );
AOI22xp5_ASAP7_75t_SL g413 ( .A1(n_26), .A2(n_38), .B1(n_414), .B2(n_431), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_27), .A2(n_62), .B1(n_482), .B2(n_485), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_28), .B(n_148), .Y(n_185) );
INVx2_ASAP7_75t_L g101 ( .A(n_29), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_31), .B(n_106), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_32), .B(n_148), .Y(n_160) );
OAI221xp5_ASAP7_75t_L g490 ( .A1(n_33), .A2(n_46), .B1(n_58), .B2(n_491), .C(n_492), .Y(n_490) );
INVxp67_ASAP7_75t_L g493 ( .A(n_33), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_35), .A2(n_55), .B1(n_465), .B2(n_470), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g119 ( .A(n_36), .B(n_106), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_37), .A2(n_71), .B1(n_158), .B2(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_39), .B(n_106), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_40), .B(n_106), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_41), .B(n_124), .Y(n_123) );
AOI22xp33_ASAP7_75t_SL g105 ( .A1(n_43), .A2(n_49), .B1(n_99), .B2(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_44), .B(n_106), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_45), .B(n_106), .Y(n_205) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_45), .Y(n_501) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_46), .A2(n_66), .B1(n_421), .B2(n_425), .Y(n_428) );
INVxp67_ASAP7_75t_L g494 ( .A(n_46), .Y(n_494) );
INVx1_ASAP7_75t_L g112 ( .A(n_50), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_51), .B(n_106), .Y(n_141) );
OAI22xp5_ASAP7_75t_SL g401 ( .A1(n_51), .A2(n_402), .B1(n_403), .B2(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_51), .Y(n_404) );
INVx1_ASAP7_75t_L g92 ( .A(n_52), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_53), .Y(n_491) );
AO32x2_ASAP7_75t_L g162 ( .A1(n_54), .A2(n_109), .A3(n_110), .B1(n_163), .B2(n_167), .Y(n_162) );
INVx1_ASAP7_75t_L g204 ( .A(n_56), .Y(n_204) );
INVx1_ASAP7_75t_L g180 ( .A(n_57), .Y(n_180) );
AO22x2_ASAP7_75t_L g430 ( .A1(n_58), .A2(n_73), .B1(n_421), .B2(n_422), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_59), .B(n_99), .Y(n_181) );
INVx1_ASAP7_75t_L g409 ( .A(n_61), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_64), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_65), .B(n_99), .Y(n_184) );
INVx2_ASAP7_75t_L g90 ( .A(n_67), .Y(n_90) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_69), .A2(n_399), .B1(n_400), .B2(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_69), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_70), .B(n_99), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g98 ( .A1(n_72), .A2(n_76), .B1(n_99), .B2(n_100), .Y(n_98) );
INVx1_ASAP7_75t_L g421 ( .A(n_74), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_74), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_75), .B(n_99), .Y(n_202) );
AOI221xp5_ASAP7_75t_SL g77 ( .A1(n_78), .A2(n_388), .B1(n_396), .B2(n_487), .C(n_499), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
AND2x2_ASAP7_75t_SL g82 ( .A(n_83), .B(n_322), .Y(n_82) );
NOR5xp2_ASAP7_75t_L g83 ( .A(n_84), .B(n_235), .C(n_281), .D(n_294), .E(n_306), .Y(n_83) );
OAI211xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_143), .B(n_189), .C(n_216), .Y(n_84) );
INVx1_ASAP7_75t_SL g317 ( .A(n_85), .Y(n_317) );
OR2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_113), .Y(n_85) );
AND2x2_ASAP7_75t_L g241 ( .A(n_86), .B(n_114), .Y(n_241) );
AND2x2_ASAP7_75t_L g269 ( .A(n_86), .B(n_215), .Y(n_269) );
AND2x2_ASAP7_75t_L g277 ( .A(n_86), .B(n_220), .Y(n_277) );
INVx3_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g207 ( .A(n_87), .B(n_115), .Y(n_207) );
INVx2_ASAP7_75t_L g219 ( .A(n_87), .Y(n_219) );
AND2x2_ASAP7_75t_L g344 ( .A(n_87), .B(n_286), .Y(n_344) );
OR2x2_ASAP7_75t_L g346 ( .A(n_87), .B(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_94), .Y(n_87) );
INVx1_ASAP7_75t_L g213 ( .A(n_88), .Y(n_213) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_89), .Y(n_109) );
INVx1_ASAP7_75t_L g129 ( .A(n_89), .Y(n_129) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_91), .Y(n_89) );
AND2x2_ASAP7_75t_SL g148 ( .A(n_90), .B(n_91), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g91 ( .A(n_92), .B(n_93), .Y(n_91) );
NAND3xp33_ASAP7_75t_L g94 ( .A(n_95), .B(n_108), .C(n_110), .Y(n_94) );
AO21x1_ASAP7_75t_L g212 ( .A1(n_95), .A2(n_108), .B(n_213), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g95 ( .A1(n_96), .A2(n_98), .B1(n_102), .B2(n_105), .Y(n_95) );
INVx2_ASAP7_75t_L g159 ( .A(n_96), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g163 ( .A1(n_96), .A2(n_104), .B1(n_164), .B2(n_166), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_96), .A2(n_102), .B1(n_171), .B2(n_172), .Y(n_170) );
BUFx6f_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx3_ASAP7_75t_L g104 ( .A(n_97), .Y(n_104) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_97), .Y(n_137) );
INVx1_ASAP7_75t_L g154 ( .A(n_97), .Y(n_154) );
INVx2_ASAP7_75t_L g133 ( .A(n_99), .Y(n_133) );
INVx3_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g107 ( .A(n_101), .Y(n_107) );
INVx1_ASAP7_75t_L g125 ( .A(n_101), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_102), .A2(n_122), .B(n_123), .Y(n_121) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_102), .A2(n_139), .B(n_140), .C(n_141), .Y(n_138) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_103), .A2(n_119), .B(n_120), .Y(n_118) );
O2A1O1Ixp5_ASAP7_75t_SL g178 ( .A1(n_103), .A2(n_179), .B(n_180), .C(n_181), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_103), .A2(n_201), .B(n_202), .Y(n_200) );
INVx5_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx3_ASAP7_75t_L g179 ( .A(n_106), .Y(n_179) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g158 ( .A(n_107), .Y(n_158) );
BUFx3_ASAP7_75t_L g165 ( .A(n_107), .Y(n_165) );
INVx4_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_109), .A2(n_117), .B(n_126), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_110), .A2(n_200), .B(n_203), .Y(n_199) );
BUFx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_111), .A2(n_118), .B(n_121), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g130 ( .A1(n_111), .A2(n_131), .B(n_138), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g149 ( .A1(n_111), .A2(n_150), .B(n_155), .Y(n_149) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_111), .A2(n_178), .B(n_182), .Y(n_177) );
INVx4_ASAP7_75t_SL g395 ( .A(n_111), .Y(n_395) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_112), .Y(n_496) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g257 ( .A(n_114), .B(n_229), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_114), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g371 ( .A(n_114), .B(n_211), .Y(n_371) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_127), .Y(n_114) );
AND2x2_ASAP7_75t_L g214 ( .A(n_115), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g261 ( .A(n_115), .Y(n_261) );
AND2x2_ASAP7_75t_L g286 ( .A(n_115), .B(n_198), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_115), .B(n_319), .Y(n_356) );
INVx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g220 ( .A(n_116), .B(n_198), .Y(n_220) );
AND2x2_ASAP7_75t_L g234 ( .A(n_116), .B(n_197), .Y(n_234) );
AND2x2_ASAP7_75t_L g251 ( .A(n_116), .B(n_127), .Y(n_251) );
AND2x2_ASAP7_75t_L g308 ( .A(n_116), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_116), .B(n_215), .Y(n_321) );
AND2x2_ASAP7_75t_L g373 ( .A(n_116), .B(n_298), .Y(n_373) );
INVx2_ASAP7_75t_L g139 ( .A(n_124), .Y(n_139) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g196 ( .A(n_127), .B(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g215 ( .A(n_127), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_127), .B(n_198), .Y(n_292) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_130), .B(n_142), .Y(n_127) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_128), .A2(n_199), .B(n_206), .Y(n_198) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_134), .C(n_135), .Y(n_131) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_136), .A2(n_183), .B(n_184), .Y(n_182) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g393 ( .A(n_137), .Y(n_393) );
O2A1O1Ixp5_ASAP7_75t_L g203 ( .A1(n_139), .A2(n_159), .B(n_204), .C(n_205), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_139), .B(n_395), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_139), .B(n_509), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_173), .B(n_186), .Y(n_143) );
INVx1_ASAP7_75t_SL g305 ( .A(n_144), .Y(n_305) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_161), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_SL g193 ( .A(n_146), .B(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
INVx1_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
AND2x2_ASAP7_75t_L g246 ( .A(n_147), .B(n_168), .Y(n_246) );
AND2x2_ASAP7_75t_L g280 ( .A(n_147), .B(n_169), .Y(n_280) );
OR2x2_ASAP7_75t_L g299 ( .A(n_147), .B(n_175), .Y(n_299) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_147), .Y(n_313) );
AND2x2_ASAP7_75t_L g326 ( .A(n_147), .B(n_327), .Y(n_326) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_160), .Y(n_147) );
INVx2_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_148), .A2(n_177), .B(n_185), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_159), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_161), .A2(n_248), .B1(n_249), .B2(n_258), .Y(n_247) );
AND2x2_ASAP7_75t_L g331 ( .A(n_161), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_168), .Y(n_161) );
INVx1_ASAP7_75t_L g192 ( .A(n_162), .Y(n_192) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_162), .Y(n_229) );
INVx1_ASAP7_75t_L g240 ( .A(n_162), .Y(n_240) );
AND2x2_ASAP7_75t_L g255 ( .A(n_162), .B(n_169), .Y(n_255) );
OR2x2_ASAP7_75t_L g209 ( .A(n_168), .B(n_194), .Y(n_209) );
AND2x2_ASAP7_75t_L g239 ( .A(n_168), .B(n_240), .Y(n_239) );
NOR2xp67_ASAP7_75t_L g327 ( .A(n_168), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g187 ( .A(n_169), .B(n_188), .Y(n_187) );
BUFx2_ASAP7_75t_L g296 ( .A(n_169), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_173), .B(n_312), .Y(n_311) );
BUFx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g274 ( .A(n_174), .B(n_240), .Y(n_274) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g186 ( .A(n_175), .B(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g245 ( .A(n_175), .Y(n_245) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g194 ( .A(n_176), .Y(n_194) );
OR2x2_ASAP7_75t_L g224 ( .A(n_176), .B(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_176), .Y(n_279) );
AOI32xp33_ASAP7_75t_L g316 ( .A1(n_186), .A2(n_246), .A3(n_317), .B1(n_318), .B2(n_320), .Y(n_316) );
AND2x2_ASAP7_75t_L g242 ( .A(n_187), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_187), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_187), .B(n_274), .Y(n_360) );
INVx1_ASAP7_75t_L g365 ( .A(n_187), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_195), .B1(n_208), .B2(n_210), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_193), .Y(n_190) );
AND2x2_ASAP7_75t_L g295 ( .A(n_191), .B(n_296), .Y(n_295) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_192), .B(n_194), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_193), .A2(n_217), .B1(n_221), .B2(n_231), .Y(n_216) );
AND2x2_ASAP7_75t_L g238 ( .A(n_193), .B(n_239), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_193), .A2(n_207), .B(n_255), .C(n_290), .Y(n_289) );
OAI332xp33_ASAP7_75t_L g294 ( .A1(n_193), .A2(n_295), .A3(n_297), .B1(n_299), .B2(n_300), .B3(n_302), .C1(n_303), .C2(n_305), .Y(n_294) );
INVx2_ASAP7_75t_L g335 ( .A(n_193), .Y(n_335) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_194), .Y(n_253) );
INVx1_ASAP7_75t_L g328 ( .A(n_194), .Y(n_328) );
AND2x2_ASAP7_75t_L g382 ( .A(n_194), .B(n_246), .Y(n_382) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_207), .Y(n_195) );
AND2x2_ASAP7_75t_L g262 ( .A(n_197), .B(n_212), .Y(n_262) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g211 ( .A(n_198), .B(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g310 ( .A(n_198), .B(n_212), .Y(n_310) );
INVx1_ASAP7_75t_L g319 ( .A(n_198), .Y(n_319) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_204), .Y(n_511) );
INVx1_ASAP7_75t_L g293 ( .A(n_207), .Y(n_293) );
INVxp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g377 ( .A(n_209), .B(n_229), .Y(n_377) );
INVx1_ASAP7_75t_SL g288 ( .A(n_210), .Y(n_288) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_214), .Y(n_210) );
AND2x2_ASAP7_75t_L g315 ( .A(n_211), .B(n_273), .Y(n_315) );
INVx1_ASAP7_75t_L g334 ( .A(n_211), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_211), .B(n_301), .Y(n_336) );
INVx1_ASAP7_75t_L g233 ( .A(n_212), .Y(n_233) );
AND2x2_ASAP7_75t_L g237 ( .A(n_214), .B(n_218), .Y(n_237) );
AND2x2_ASAP7_75t_L g304 ( .A(n_214), .B(n_262), .Y(n_304) );
INVx2_ASAP7_75t_L g347 ( .A(n_214), .Y(n_347) );
INVx2_ASAP7_75t_L g230 ( .A(n_215), .Y(n_230) );
AND2x2_ASAP7_75t_L g232 ( .A(n_215), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
INVx1_ASAP7_75t_L g248 ( .A(n_218), .Y(n_248) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_219), .B(n_292), .Y(n_298) );
OR2x2_ASAP7_75t_L g362 ( .A(n_219), .B(n_321), .Y(n_362) );
INVx1_ASAP7_75t_L g386 ( .A(n_219), .Y(n_386) );
INVx1_ASAP7_75t_L g342 ( .A(n_220), .Y(n_342) );
AND2x2_ASAP7_75t_L g387 ( .A(n_220), .B(n_230), .Y(n_387) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_226), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_224), .A2(n_250), .B1(n_252), .B2(n_256), .Y(n_249) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OAI322xp33_ASAP7_75t_SL g333 ( .A1(n_227), .A2(n_334), .A3(n_335), .B1(n_336), .B2(n_337), .C1(n_340), .C2(n_342), .Y(n_333) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
AND2x2_ASAP7_75t_L g330 ( .A(n_228), .B(n_246), .Y(n_330) );
OR2x2_ASAP7_75t_L g364 ( .A(n_228), .B(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g367 ( .A(n_228), .B(n_299), .Y(n_367) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g312 ( .A(n_229), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g368 ( .A(n_229), .B(n_299), .Y(n_368) );
INVx3_ASAP7_75t_L g301 ( .A(n_230), .Y(n_301) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g357 ( .A(n_232), .Y(n_357) );
AOI222xp33_ASAP7_75t_L g236 ( .A1(n_234), .A2(n_237), .B1(n_238), .B2(n_241), .C1(n_242), .C2(n_244), .Y(n_236) );
INVx1_ASAP7_75t_L g267 ( .A(n_234), .Y(n_267) );
NAND3xp33_ASAP7_75t_SL g235 ( .A(n_236), .B(n_247), .C(n_264), .Y(n_235) );
AND2x2_ASAP7_75t_L g352 ( .A(n_239), .B(n_253), .Y(n_352) );
BUFx2_ASAP7_75t_L g243 ( .A(n_240), .Y(n_243) );
INVx1_ASAP7_75t_L g284 ( .A(n_240), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_241), .A2(n_277), .B1(n_330), .B2(n_331), .C(n_333), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_243), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_246), .Y(n_270) );
AND2x2_ASAP7_75t_L g283 ( .A(n_246), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_251), .B(n_262), .Y(n_263) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
OAI21xp33_ASAP7_75t_L g258 ( .A1(n_253), .A2(n_259), .B(n_263), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_253), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g350 ( .A(n_255), .B(n_332), .Y(n_350) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g273 ( .A(n_261), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_262), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g379 ( .A(n_262), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_270), .B1(n_271), .B2(n_274), .C(n_275), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_266), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g375 ( .A(n_274), .B(n_280), .Y(n_375) );
INVxp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OAI31xp33_ASAP7_75t_SL g343 ( .A1(n_278), .A2(n_317), .A3(n_344), .B(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g332 ( .A(n_279), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_280), .B(n_284), .Y(n_383) );
OAI221xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_285), .B1(n_287), .B2(n_288), .C(n_289), .Y(n_281) );
INVx1_ASAP7_75t_L g287 ( .A(n_283), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_286), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g302 ( .A(n_295), .Y(n_302) );
INVx2_ASAP7_75t_L g338 ( .A(n_296), .Y(n_338) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g324 ( .A(n_301), .B(n_310), .Y(n_324) );
A2O1A1Ixp33_ASAP7_75t_L g374 ( .A1(n_301), .A2(n_318), .B(n_375), .C(n_376), .Y(n_374) );
OAI221xp5_ASAP7_75t_SL g306 ( .A1(n_302), .A2(n_307), .B1(n_311), .B2(n_314), .C(n_316), .Y(n_306) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_L g369 ( .A1(n_305), .A2(n_370), .B(n_372), .C(n_374), .Y(n_369) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g358 ( .A1(n_308), .A2(n_359), .B1(n_361), .B2(n_363), .C(n_366), .Y(n_358) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
NOR4xp25_ASAP7_75t_L g322 ( .A(n_323), .B(n_348), .C(n_369), .D(n_380), .Y(n_322) );
OAI211xp5_ASAP7_75t_SL g323 ( .A1(n_324), .A2(n_325), .B(n_329), .C(n_343), .Y(n_323) );
INVx1_ASAP7_75t_SL g378 ( .A(n_330), .Y(n_378) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_SL g341 ( .A(n_339), .Y(n_341) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_346), .A2(n_355), .B1(n_367), .B2(n_368), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B(n_353), .C(n_358), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI31xp33_ASAP7_75t_L g380 ( .A1(n_351), .A2(n_381), .A3(n_383), .B(n_384), .Y(n_380) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_389), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_394), .Y(n_390) );
INVx1_ASAP7_75t_L g509 ( .A(n_391), .Y(n_509) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
XOR2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_407), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_398), .Y(n_406) );
CKINVDCx16_ASAP7_75t_R g400 ( .A(n_401), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_402), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B1(n_411), .B2(n_486), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_408), .Y(n_486) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_410), .A2(n_411), .B1(n_501), .B2(n_502), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND4xp75_ASAP7_75t_SL g412 ( .A(n_413), .B(n_437), .C(n_444), .D(n_458), .Y(n_412) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx11_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x6_ASAP7_75t_L g416 ( .A(n_417), .B(n_426), .Y(n_416) );
AND2x4_ASAP7_75t_L g484 ( .A(n_417), .B(n_457), .Y(n_484) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_424), .Y(n_418) );
AND2x2_ASAP7_75t_L g436 ( .A(n_419), .B(n_424), .Y(n_436) );
AND2x2_ASAP7_75t_L g440 ( .A(n_419), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g463 ( .A(n_420), .B(n_424), .Y(n_463) );
AND2x2_ASAP7_75t_L g469 ( .A(n_420), .B(n_428), .Y(n_469) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_423), .Y(n_425) );
INVx2_ASAP7_75t_L g441 ( .A(n_424), .Y(n_441) );
INVx1_ASAP7_75t_L g480 ( .A(n_424), .Y(n_480) );
AND2x2_ASAP7_75t_L g439 ( .A(n_426), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g443 ( .A(n_426), .B(n_436), .Y(n_443) );
AND2x6_ASAP7_75t_L g462 ( .A(n_426), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
AND2x2_ASAP7_75t_L g457 ( .A(n_427), .B(n_430), .Y(n_457) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g434 ( .A(n_428), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_428), .B(n_430), .Y(n_449) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g435 ( .A(n_430), .Y(n_435) );
INVx1_ASAP7_75t_L g468 ( .A(n_430), .Y(n_468) );
INVx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx8_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
AND2x2_ASAP7_75t_L g454 ( .A(n_434), .B(n_440), .Y(n_454) );
INVx1_ASAP7_75t_L g471 ( .A(n_435), .Y(n_471) );
AND2x6_ASAP7_75t_L g485 ( .A(n_436), .B(n_457), .Y(n_485) );
BUFx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g447 ( .A(n_440), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g456 ( .A(n_440), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g451 ( .A(n_441), .Y(n_451) );
AND2x2_ASAP7_75t_L g476 ( .A(n_441), .B(n_468), .Y(n_476) );
BUFx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_452), .Y(n_444) );
BUFx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g450 ( .A(n_448), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_472), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_464), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g470 ( .A(n_463), .B(n_471), .Y(n_470) );
BUFx12f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g475 ( .A(n_469), .B(n_476), .Y(n_475) );
AND2x4_ASAP7_75t_L g478 ( .A(n_469), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_481), .Y(n_472) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx5_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx4_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
AND3x1_ASAP7_75t_SL g489 ( .A(n_490), .B(n_495), .C(n_497), .Y(n_489) );
INVxp67_ASAP7_75t_L g504 ( .A(n_490), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx1_ASAP7_75t_SL g505 ( .A(n_495), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_495), .A2(n_508), .B(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g516 ( .A(n_495), .Y(n_516) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_496), .B(n_498), .Y(n_510) );
OR2x2_ASAP7_75t_SL g515 ( .A(n_497), .B(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
OAI322xp33_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_503), .A3(n_505), .B1(n_506), .B2(n_511), .C1(n_512), .C2(n_513), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_501), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
endmodule