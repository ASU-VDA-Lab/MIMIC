module real_aes_2629_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_0), .B(n_133), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_1), .A2(n_142), .B(n_147), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_2), .B(n_447), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_3), .A2(n_4), .B1(n_802), .B2(n_803), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_3), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_4), .Y(n_802) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_5), .B(n_149), .Y(n_188) );
INVx1_ASAP7_75t_L g140 ( .A(n_6), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_7), .B(n_149), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_8), .B(n_158), .Y(n_516) );
INVx1_ASAP7_75t_L g499 ( .A(n_9), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_10), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_11), .Y(n_474) );
NAND2xp33_ASAP7_75t_L g231 ( .A(n_12), .B(n_151), .Y(n_231) );
INVx2_ASAP7_75t_L g130 ( .A(n_13), .Y(n_130) );
AOI221x1_ASAP7_75t_L g173 ( .A1(n_14), .A2(n_28), .B1(n_133), .B2(n_142), .C(n_174), .Y(n_173) );
OAI22xp5_ASAP7_75t_SL g799 ( .A1(n_15), .A2(n_800), .B1(n_801), .B2(n_804), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_15), .Y(n_804) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_16), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_17), .B(n_133), .Y(n_227) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_18), .A2(n_225), .B(n_226), .Y(n_224) );
INVx1_ASAP7_75t_L g524 ( .A(n_19), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_20), .B(n_153), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_21), .A2(n_81), .B1(n_439), .B2(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_21), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_22), .B(n_149), .Y(n_162) );
AO21x1_ASAP7_75t_L g183 ( .A1(n_23), .A2(n_133), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g114 ( .A(n_24), .Y(n_114) );
INVx1_ASAP7_75t_L g522 ( .A(n_25), .Y(n_522) );
INVx1_ASAP7_75t_SL g510 ( .A(n_26), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_27), .B(n_134), .Y(n_565) );
NAND2x1_ASAP7_75t_L g205 ( .A(n_29), .B(n_149), .Y(n_205) );
AOI33xp33_ASAP7_75t_L g545 ( .A1(n_30), .A2(n_54), .A3(n_464), .B1(n_479), .B2(n_546), .B3(n_547), .Y(n_545) );
NAND2x1_ASAP7_75t_L g238 ( .A(n_31), .B(n_151), .Y(n_238) );
INVx1_ASAP7_75t_L g467 ( .A(n_32), .Y(n_467) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_33), .A2(n_88), .B(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g155 ( .A(n_33), .B(n_88), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_34), .B(n_482), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_35), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_36), .B(n_149), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_37), .B(n_151), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_38), .A2(n_142), .B(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g139 ( .A(n_39), .B(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g143 ( .A(n_39), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g478 ( .A(n_39), .Y(n_478) );
OR2x6_ASAP7_75t_L g112 ( .A(n_40), .B(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_41), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_42), .B(n_133), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_43), .B(n_482), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_44), .A2(n_128), .B1(n_158), .B2(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_45), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_46), .B(n_134), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_47), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_48), .B(n_151), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_49), .B(n_225), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_50), .B(n_134), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_51), .A2(n_142), .B(n_237), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_52), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_53), .B(n_151), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_55), .B(n_134), .Y(n_493) );
INVx1_ASAP7_75t_L g136 ( .A(n_56), .Y(n_136) );
INVx1_ASAP7_75t_L g146 ( .A(n_56), .Y(n_146) );
AND2x2_ASAP7_75t_L g494 ( .A(n_57), .B(n_153), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_58), .A2(n_76), .B1(n_476), .B2(n_482), .C(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_59), .B(n_482), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_60), .B(n_149), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_61), .B(n_128), .Y(n_480) );
AOI21xp5_ASAP7_75t_SL g532 ( .A1(n_62), .A2(n_476), .B(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_63), .A2(n_142), .B(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g519 ( .A(n_64), .Y(n_519) );
AO21x1_ASAP7_75t_L g185 ( .A1(n_65), .A2(n_142), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_66), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g492 ( .A(n_67), .Y(n_492) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_68), .A2(n_103), .B1(n_444), .B2(n_449), .C1(n_819), .C2(n_825), .Y(n_102) );
XNOR2x1_ASAP7_75t_L g116 ( .A(n_68), .B(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_69), .B(n_133), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_70), .A2(n_476), .B(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_71), .Y(n_806) );
AND2x2_ASAP7_75t_L g199 ( .A(n_72), .B(n_154), .Y(n_199) );
INVx1_ASAP7_75t_L g138 ( .A(n_73), .Y(n_138) );
INVx1_ASAP7_75t_L g144 ( .A(n_73), .Y(n_144) );
AND2x2_ASAP7_75t_L g242 ( .A(n_74), .B(n_127), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_75), .B(n_482), .Y(n_548) );
AND2x2_ASAP7_75t_L g512 ( .A(n_77), .B(n_127), .Y(n_512) );
INVx1_ASAP7_75t_L g520 ( .A(n_78), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_79), .A2(n_476), .B(n_509), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_80), .A2(n_476), .B(n_540), .C(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g440 ( .A(n_81), .Y(n_440) );
INVx1_ASAP7_75t_L g115 ( .A(n_82), .Y(n_115) );
AND2x2_ASAP7_75t_L g126 ( .A(n_83), .B(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_84), .B(n_133), .Y(n_164) );
AND2x2_ASAP7_75t_SL g530 ( .A(n_85), .B(n_127), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_86), .A2(n_476), .B1(n_543), .B2(n_544), .Y(n_542) );
AND2x2_ASAP7_75t_L g184 ( .A(n_87), .B(n_158), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_89), .B(n_151), .Y(n_163) );
AND2x2_ASAP7_75t_L g208 ( .A(n_90), .B(n_127), .Y(n_208) );
INVx1_ASAP7_75t_L g534 ( .A(n_91), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_92), .B(n_149), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_93), .A2(n_142), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_94), .B(n_151), .Y(n_175) );
AND2x2_ASAP7_75t_L g549 ( .A(n_95), .B(n_127), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_96), .B(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_97), .A2(n_462), .B(n_466), .C(n_469), .Y(n_461) );
BUFx2_ASAP7_75t_L g448 ( .A(n_98), .Y(n_448) );
BUFx2_ASAP7_75t_SL g831 ( .A(n_98), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_99), .A2(n_142), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_100), .B(n_134), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_101), .B(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI21x1_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_116), .B(n_441), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g443 ( .A(n_109), .Y(n_443) );
BUFx2_ASAP7_75t_L g824 ( .A(n_109), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x6_ASAP7_75t_SL g796 ( .A(n_110), .B(n_111), .Y(n_796) );
AND2x6_ASAP7_75t_SL g798 ( .A(n_110), .B(n_112), .Y(n_798) );
OR2x2_ASAP7_75t_L g809 ( .A(n_110), .B(n_112), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
XOR2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_438), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_118), .A2(n_452), .B1(n_794), .B2(n_797), .Y(n_451) );
INVx3_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g814 ( .A(n_119), .Y(n_814) );
NOR2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_325), .Y(n_119) );
AO211x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_167), .B(n_218), .C(n_293), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
AND3x2_ASAP7_75t_L g374 ( .A(n_123), .B(n_255), .C(n_271), .Y(n_374) );
AND2x4_ASAP7_75t_L g377 ( .A(n_123), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_156), .Y(n_123) );
NAND2x1p5_ASAP7_75t_L g232 ( .A(n_124), .B(n_233), .Y(n_232) );
INVx4_ASAP7_75t_L g286 ( .A(n_124), .Y(n_286) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_124), .B(n_280), .Y(n_371) );
AND2x2_ASAP7_75t_L g414 ( .A(n_124), .B(n_234), .Y(n_414) );
INVx5_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g263 ( .A(n_125), .Y(n_263) );
AND2x2_ASAP7_75t_L g282 ( .A(n_125), .B(n_224), .Y(n_282) );
AND2x2_ASAP7_75t_L g300 ( .A(n_125), .B(n_234), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_125), .B(n_233), .Y(n_360) );
NOR2x1_ASAP7_75t_SL g387 ( .A(n_125), .B(n_156), .Y(n_387) );
OR2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_131), .Y(n_125) );
INVx3_ASAP7_75t_L g198 ( .A(n_127), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_127), .A2(n_198), .B1(n_461), .B2(n_470), .Y(n_460) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_128), .B(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx4f_ASAP7_75t_L g225 ( .A(n_129), .Y(n_225) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_130), .B(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g158 ( .A(n_130), .B(n_155), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_141), .B(n_153), .Y(n_131) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_139), .Y(n_133) );
INVx1_ASAP7_75t_L g468 ( .A(n_134), .Y(n_468) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
AND2x6_ASAP7_75t_L g151 ( .A(n_135), .B(n_144), .Y(n_151) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g149 ( .A(n_137), .B(n_146), .Y(n_149) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx5_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_139), .Y(n_469) );
AND2x2_ASAP7_75t_L g145 ( .A(n_140), .B(n_146), .Y(n_145) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_140), .Y(n_484) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
BUFx3_ASAP7_75t_L g485 ( .A(n_143), .Y(n_485) );
INVx2_ASAP7_75t_L g465 ( .A(n_144), .Y(n_465) );
AND2x4_ASAP7_75t_L g476 ( .A(n_145), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g464 ( .A(n_146), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_150), .B(n_152), .Y(n_147) );
INVxp67_ASAP7_75t_L g525 ( .A(n_149), .Y(n_525) );
INVxp67_ASAP7_75t_L g523 ( .A(n_151), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_152), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_152), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_152), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_152), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_152), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_152), .A2(n_230), .B(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_152), .A2(n_238), .B(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_152), .A2(n_463), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g498 ( .A1(n_152), .A2(n_463), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_SL g509 ( .A1(n_152), .A2(n_463), .B(n_510), .C(n_511), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_152), .B(n_158), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_152), .A2(n_463), .B(n_534), .C(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g543 ( .A(n_152), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_152), .A2(n_565), .B(n_566), .Y(n_564) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_153), .A2(n_173), .B(n_177), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_153), .Y(n_241) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_153), .A2(n_173), .B(n_177), .Y(n_246) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_156), .B(n_224), .Y(n_223) );
AO21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_165), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_157), .B(n_166), .Y(n_165) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_157), .A2(n_159), .B(n_165), .Y(n_259) );
INVx1_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_158), .B(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_158), .A2(n_227), .B(n_228), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_158), .A2(n_532), .B(n_536), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
AO21x1_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_200), .B(n_209), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp33_ASAP7_75t_L g268 ( .A1(n_169), .A2(n_269), .B1(n_273), .B2(n_274), .Y(n_268) );
OR2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_178), .Y(n_169) );
AND2x2_ASAP7_75t_L g329 ( .A(n_170), .B(n_215), .Y(n_329) );
BUFx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x4_ASAP7_75t_L g262 ( .A(n_171), .B(n_245), .Y(n_262) );
AND2x2_ASAP7_75t_L g334 ( .A(n_171), .B(n_217), .Y(n_334) );
AND2x2_ASAP7_75t_L g353 ( .A(n_171), .B(n_319), .Y(n_353) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g210 ( .A(n_172), .Y(n_210) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_172), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_178), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g313 ( .A(n_179), .B(n_212), .Y(n_313) );
AND2x4_ASAP7_75t_L g179 ( .A(n_180), .B(n_191), .Y(n_179) );
AND2x2_ASAP7_75t_L g215 ( .A(n_180), .B(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g250 ( .A(n_180), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_SL g310 ( .A(n_180), .B(n_246), .Y(n_310) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx2_ASAP7_75t_L g403 ( .A(n_181), .Y(n_403) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g245 ( .A(n_182), .Y(n_245) );
OAI21x1_ASAP7_75t_SL g182 ( .A1(n_183), .A2(n_185), .B(n_189), .Y(n_182) );
INVx1_ASAP7_75t_L g190 ( .A(n_184), .Y(n_190) );
INVx2_ASAP7_75t_L g251 ( .A(n_191), .Y(n_251) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_191), .Y(n_351) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_198), .B(n_199), .Y(n_191) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_192), .A2(n_198), .B(n_199), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_193), .B(n_197), .Y(n_192) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_198), .A2(n_202), .B(n_208), .Y(n_201) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_198), .A2(n_202), .B(n_208), .Y(n_214) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_198), .A2(n_488), .B(n_494), .Y(n_487) );
AO21x2_ASAP7_75t_L g581 ( .A1(n_198), .A2(n_488), .B(n_494), .Y(n_581) );
INVx2_ASAP7_75t_L g247 ( .A(n_200), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_200), .B(n_379), .Y(n_405) );
AND2x2_ASAP7_75t_L g424 ( .A(n_200), .B(n_414), .Y(n_424) );
BUFx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x4_ASAP7_75t_SL g292 ( .A(n_201), .B(n_251), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_207), .Y(n_202) );
AND2x2_ASAP7_75t_SL g209 ( .A(n_210), .B(n_211), .Y(n_209) );
AND2x2_ASAP7_75t_L g291 ( .A(n_210), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_210), .B(n_261), .Y(n_296) );
INVx1_ASAP7_75t_SL g423 ( .A(n_210), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_211), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_215), .Y(n_211) );
INVx1_ASAP7_75t_L g249 ( .A(n_212), .Y(n_249) );
AND2x2_ASAP7_75t_L g435 ( .A(n_212), .B(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g311 ( .A(n_213), .B(n_216), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_213), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g365 ( .A(n_213), .B(n_217), .Y(n_365) );
AND2x2_ASAP7_75t_L g396 ( .A(n_213), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g261 ( .A(n_214), .B(n_217), .Y(n_261) );
INVxp67_ASAP7_75t_L g278 ( .A(n_214), .Y(n_278) );
BUFx3_ASAP7_75t_L g319 ( .A(n_214), .Y(n_319) );
AND2x2_ASAP7_75t_L g339 ( .A(n_215), .B(n_340), .Y(n_339) );
NAND2xp33_ASAP7_75t_L g352 ( .A(n_215), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_216), .B(n_245), .Y(n_308) );
AND2x2_ASAP7_75t_L g397 ( .A(n_216), .B(n_246), .Y(n_397) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g324 ( .A(n_217), .B(n_246), .Y(n_324) );
OR3x1_ASAP7_75t_L g218 ( .A(n_219), .B(n_268), .C(n_283), .Y(n_218) );
OAI321xp33_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_232), .A3(n_243), .B1(n_248), .B2(n_252), .C(n_260), .Y(n_219) );
INVx1_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_223), .Y(n_299) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_223), .Y(n_317) );
OR2x2_ASAP7_75t_L g321 ( .A(n_223), .B(n_232), .Y(n_321) );
BUFx3_ASAP7_75t_L g255 ( .A(n_224), .Y(n_255) );
AND2x2_ASAP7_75t_L g272 ( .A(n_224), .B(n_258), .Y(n_272) );
INVx1_ASAP7_75t_L g289 ( .A(n_224), .Y(n_289) );
INVx2_ASAP7_75t_L g305 ( .A(n_224), .Y(n_305) );
OR2x2_ASAP7_75t_L g344 ( .A(n_224), .B(n_233), .Y(n_344) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_225), .A2(n_497), .B(n_501), .Y(n_496) );
INVx2_ASAP7_75t_SL g540 ( .A(n_225), .Y(n_540) );
INVx2_ASAP7_75t_L g332 ( .A(n_232), .Y(n_332) );
AND2x2_ASAP7_75t_L g256 ( .A(n_233), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g271 ( .A(n_233), .Y(n_271) );
AND2x4_ASAP7_75t_L g280 ( .A(n_233), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_233), .B(n_257), .Y(n_303) );
AND2x2_ASAP7_75t_L g410 ( .A(n_233), .B(n_305), .Y(n_410) );
INVx4_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_234), .Y(n_369) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_241), .B(n_242), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_240), .Y(n_235) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_241), .A2(n_506), .B(n_512), .Y(n_505) );
INVx1_ASAP7_75t_L g297 ( .A(n_243), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_244), .B(n_247), .Y(n_243) );
AND2x2_ASAP7_75t_L g384 ( .A(n_244), .B(n_311), .Y(n_384) );
INVx1_ASAP7_75t_SL g401 ( .A(n_244), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_244), .B(n_377), .Y(n_430) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
OR2x2_ASAP7_75t_L g273 ( .A(n_245), .B(n_246), .Y(n_273) );
AND2x2_ASAP7_75t_L g366 ( .A(n_247), .B(n_262), .Y(n_366) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_251), .B(n_262), .Y(n_389) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_253), .A2(n_402), .B1(n_407), .B2(n_409), .Y(n_406) );
AND2x4_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
AND2x2_ASAP7_75t_L g331 ( .A(n_254), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g426 ( .A(n_254), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g382 ( .A(n_255), .B(n_300), .Y(n_382) );
AND2x4_ASAP7_75t_L g336 ( .A(n_256), .B(n_282), .Y(n_336) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_258), .Y(n_434) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g267 ( .A(n_259), .Y(n_267) );
INVx1_ASAP7_75t_L g281 ( .A(n_259), .Y(n_281) );
NAND4xp25_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .C(n_263), .D(n_264), .Y(n_260) );
AND2x2_ASAP7_75t_L g418 ( .A(n_261), .B(n_403), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_261), .B(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_262), .B(n_338), .Y(n_337) );
OAI322xp33_ASAP7_75t_L g345 ( .A1(n_262), .A2(n_346), .A3(n_350), .B1(n_352), .B2(n_354), .C1(n_356), .C2(n_361), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_262), .B(n_311), .Y(n_361) );
INVx1_ASAP7_75t_L g429 ( .A(n_262), .Y(n_429) );
INVx2_ASAP7_75t_L g275 ( .A(n_263), .Y(n_275) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_266), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_267), .B(n_286), .Y(n_343) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_270), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
AND2x2_ASAP7_75t_L g388 ( .A(n_271), .B(n_299), .Y(n_388) );
AOI31xp33_ASAP7_75t_L g274 ( .A1(n_272), .A2(n_275), .A3(n_276), .B(n_279), .Y(n_274) );
AND2x2_ASAP7_75t_L g285 ( .A(n_272), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g413 ( .A(n_272), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_272), .B(n_300), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_272), .Y(n_421) );
INVx1_ASAP7_75t_SL g379 ( .A(n_273), .Y(n_379) );
NAND3xp33_ASAP7_75t_SL g407 ( .A(n_273), .B(n_401), .C(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g307 ( .A(n_278), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
AND2x2_ASAP7_75t_L g288 ( .A(n_280), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g349 ( .A(n_280), .Y(n_349) );
AOI322xp5_ASAP7_75t_L g431 ( .A1(n_280), .A2(n_310), .A3(n_313), .B1(n_432), .B2(n_433), .C1(n_435), .C2(n_437), .Y(n_431) );
AND2x2_ASAP7_75t_L g437 ( .A(n_280), .B(n_286), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_287), .B(n_290), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_286), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g432 ( .A(n_286), .B(n_319), .Y(n_432) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g358 ( .A(n_289), .Y(n_358) );
AND2x2_ASAP7_75t_L g386 ( .A(n_289), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g433 ( .A(n_289), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g338 ( .A(n_292), .Y(n_338) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
O2A1O1Ixp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_297), .B(n_298), .C(n_301), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x2_ASAP7_75t_L g355 ( .A(n_300), .B(n_305), .Y(n_355) );
OAI211xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_306), .B(n_312), .C(n_314), .Y(n_301) );
OAI221xp5_ASAP7_75t_L g327 ( .A1(n_302), .A2(n_328), .B1(n_330), .B2(n_333), .C(n_335), .Y(n_327) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g347 ( .A(n_304), .Y(n_347) );
OR2x2_ASAP7_75t_L g367 ( .A(n_304), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g412 ( .A(n_307), .Y(n_412) );
INVx1_ASAP7_75t_L g436 ( .A(n_308), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g318 ( .A(n_310), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_310), .B(n_380), .Y(n_392) );
INVx1_ASAP7_75t_L g372 ( .A(n_311), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B1(n_320), .B2(n_322), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_SL g380 ( .A(n_319), .Y(n_380) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND4xp75_ASAP7_75t_L g325 ( .A(n_326), .B(n_362), .C(n_390), .D(n_415), .Y(n_325) );
NOR2xp67_ASAP7_75t_L g326 ( .A(n_327), .B(n_345), .Y(n_326) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_SL g402 ( .A(n_334), .B(n_403), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_339), .B2(n_341), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_338), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx2_ASAP7_75t_L g378 ( .A(n_344), .Y(n_378) );
OR2x2_ASAP7_75t_L g393 ( .A(n_344), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g408 ( .A(n_353), .Y(n_408) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
OAI21xp5_ASAP7_75t_SL g399 ( .A1(n_355), .A2(n_400), .B(n_402), .Y(n_399) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_363), .B(n_375), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_367), .B1(n_370), .B2(n_372), .C(n_373), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_365), .A2(n_412), .B(n_413), .Y(n_411) );
INVx3_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OAI322xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .A3(n_380), .B1(n_381), .B2(n_383), .C1(n_385), .C2(n_389), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVx1_ASAP7_75t_L g398 ( .A(n_386), .Y(n_398) );
INVx1_ASAP7_75t_L g394 ( .A(n_387), .Y(n_394) );
AND2x2_ASAP7_75t_L g409 ( .A(n_387), .B(n_410), .Y(n_409) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_391), .B(n_404), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_395), .B2(n_398), .C(n_399), .Y(n_391) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OAI211xp5_ASAP7_75t_SL g404 ( .A1(n_398), .A2(n_405), .B(n_406), .C(n_411), .Y(n_404) );
INVx2_ASAP7_75t_SL g427 ( .A(n_414), .Y(n_427) );
NOR2x1_ASAP7_75t_L g415 ( .A(n_416), .B(n_425), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_421), .B2(n_422), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
OAI211xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_428), .B(n_430), .C(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g832 ( .A(n_443), .Y(n_832) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_SL g445 ( .A(n_446), .B(n_448), .Y(n_445) );
INVx2_ASAP7_75t_L g823 ( .A(n_446), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_446), .A2(n_829), .B(n_832), .Y(n_828) );
NAND2xp5_ASAP7_75t_SL g822 ( .A(n_448), .B(n_823), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_810), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_799), .B(n_805), .Y(n_450) );
INVxp67_ASAP7_75t_SL g812 ( .A(n_452), .Y(n_812) );
NAND3x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_673), .C(n_740), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_633), .Y(n_453) );
NOR3x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_584), .C(n_613), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_502), .B1(n_537), .B2(n_552), .C(n_569), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_SL g747 ( .A1(n_456), .A2(n_514), .B(n_748), .C(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_457), .A2(n_719), .B1(n_722), .B2(n_724), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_457), .B(n_538), .Y(n_793) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_486), .Y(n_457) );
BUFx2_ASAP7_75t_L g712 ( .A(n_458), .Y(n_712) );
INVx1_ASAP7_75t_SL g725 ( .A(n_458), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_458), .B(n_580), .Y(n_767) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g550 ( .A(n_459), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g595 ( .A(n_459), .B(n_496), .Y(n_595) );
INVx1_ASAP7_75t_L g606 ( .A(n_459), .Y(n_606) );
INVx2_ASAP7_75t_L g610 ( .A(n_459), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_459), .B(n_581), .Y(n_737) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .Y(n_459) );
INVxp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_463), .A2(n_468), .B1(n_519), .B2(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g567 ( .A(n_463), .Y(n_567) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
AND2x2_ASAP7_75t_L g483 ( .A(n_464), .B(n_484), .Y(n_483) );
INVxp33_ASAP7_75t_L g546 ( .A(n_464), .Y(n_546) );
INVx3_ASAP7_75t_L g479 ( .A(n_465), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_475), .B1(n_480), .B2(n_481), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVxp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2x1p5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g547 ( .A(n_479), .Y(n_547) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
INVx1_ASAP7_75t_L g560 ( .A(n_483), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_485), .Y(n_561) );
AND2x2_ASAP7_75t_L g686 ( .A(n_486), .B(n_687), .Y(n_686) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_487), .B(n_495), .Y(n_486) );
INVx2_ASAP7_75t_L g589 ( .A(n_487), .Y(n_589) );
AND2x2_ASAP7_75t_L g609 ( .A(n_487), .B(n_610), .Y(n_609) );
NOR2xp67_ASAP7_75t_L g734 ( .A(n_487), .B(n_610), .Y(n_734) );
AND2x2_ASAP7_75t_L g759 ( .A(n_487), .B(n_602), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g551 ( .A(n_496), .Y(n_551) );
INVx1_ASAP7_75t_L g573 ( .A(n_496), .Y(n_573) );
INVxp67_ASAP7_75t_L g612 ( .A(n_496), .Y(n_612) );
AND2x4_ASAP7_75t_L g652 ( .A(n_496), .B(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_496), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_496), .B(n_603), .Y(n_738) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_513), .Y(n_503) );
AND2x2_ASAP7_75t_L g626 ( .A(n_504), .B(n_598), .Y(n_626) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_505), .Y(n_554) );
AND2x2_ASAP7_75t_L g582 ( .A(n_505), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g593 ( .A(n_505), .Y(n_593) );
INVx1_ASAP7_75t_L g617 ( .A(n_505), .Y(n_617) );
AND2x2_ASAP7_75t_L g620 ( .A(n_505), .B(n_515), .Y(n_620) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_505), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
NOR2x1_ASAP7_75t_L g513 ( .A(n_514), .B(n_527), .Y(n_513) );
AND2x2_ASAP7_75t_L g607 ( .A(n_514), .B(n_529), .Y(n_607) );
NAND2x1_ASAP7_75t_L g640 ( .A(n_514), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g743 ( .A(n_514), .Y(n_743) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx3_ASAP7_75t_L g583 ( .A(n_515), .Y(n_583) );
AND2x2_ASAP7_75t_L g598 ( .A(n_515), .B(n_557), .Y(n_598) );
NOR2x1_ASAP7_75t_SL g667 ( .A(n_515), .B(n_529), .Y(n_667) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_521), .B(n_526), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_524), .B2(n_525), .Y(n_521) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_527), .B(n_691), .Y(n_704) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g629 ( .A(n_528), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g568 ( .A(n_529), .Y(n_568) );
AND2x4_ASAP7_75t_L g575 ( .A(n_529), .B(n_576), .Y(n_575) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_529), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_529), .B(n_592), .Y(n_692) );
AND2x2_ASAP7_75t_L g720 ( .A(n_529), .B(n_557), .Y(n_720) );
OR2x6_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
NAND2x1_ASAP7_75t_SL g537 ( .A(n_538), .B(n_550), .Y(n_537) );
OR2x2_ASAP7_75t_L g748 ( .A(n_538), .B(n_660), .Y(n_748) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_L g588 ( .A(n_539), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g653 ( .A(n_539), .Y(n_653) );
AND2x2_ASAP7_75t_L g687 ( .A(n_539), .B(n_610), .Y(n_687) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B(n_549), .Y(n_539) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_540), .A2(n_541), .B(n_549), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_542), .B(n_548), .Y(n_541) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx3_ASAP7_75t_L g660 ( .A(n_550), .Y(n_660) );
AND2x2_ASAP7_75t_L g668 ( .A(n_550), .B(n_601), .Y(n_668) );
AND2x2_ASAP7_75t_L g785 ( .A(n_550), .B(n_588), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
BUFx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g739 ( .A(n_554), .B(n_680), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_554), .B(n_579), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_555), .A2(n_616), .B(n_619), .Y(n_615) );
AND2x2_ASAP7_75t_L g685 ( .A(n_555), .B(n_591), .Y(n_685) );
INVx2_ASAP7_75t_SL g772 ( .A(n_555), .Y(n_772) );
AND2x4_ASAP7_75t_SL g555 ( .A(n_556), .B(n_568), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g576 ( .A(n_557), .Y(n_576) );
INVx2_ASAP7_75t_L g623 ( .A(n_557), .Y(n_623) );
AND2x4_ASAP7_75t_L g630 ( .A(n_557), .B(n_583), .Y(n_630) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_563), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .C(n_562), .Y(n_559) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_568), .Y(n_586) );
AND2x4_ASAP7_75t_L g662 ( .A(n_568), .B(n_576), .Y(n_662) );
OR2x2_ASAP7_75t_L g788 ( .A(n_568), .B(n_789), .Y(n_788) );
NAND4xp25_ASAP7_75t_L g569 ( .A(n_570), .B(n_574), .C(n_577), .D(n_582), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g635 ( .A(n_571), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g732 ( .A(n_571), .Y(n_732) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g632 ( .A(n_572), .B(n_580), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_572), .B(n_637), .Y(n_766) );
BUFx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_575), .B(n_591), .Y(n_644) );
INVx2_ASAP7_75t_L g746 ( .A(n_575), .Y(n_746) );
AND2x2_ASAP7_75t_SL g756 ( .A(n_575), .B(n_616), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_575), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g648 ( .A(n_579), .B(n_595), .Y(n_648) );
AND2x2_ASAP7_75t_L g716 ( .A(n_579), .B(n_652), .Y(n_716) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g601 ( .A(n_580), .B(n_602), .Y(n_601) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_581), .Y(n_655) );
AND2x2_ASAP7_75t_L g706 ( .A(n_581), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_581), .B(n_603), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_582), .B(n_746), .Y(n_753) );
INVx1_ASAP7_75t_SL g789 ( .A(n_582), .Y(n_789) );
INVx1_ASAP7_75t_L g618 ( .A(n_583), .Y(n_618) );
AND2x2_ASAP7_75t_L g680 ( .A(n_583), .B(n_623), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_594), .B(n_596), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
AND2x2_ASAP7_75t_L g646 ( .A(n_588), .B(n_595), .Y(n_646) );
AND2x2_ASAP7_75t_L g754 ( .A(n_588), .B(n_605), .Y(n_754) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g628 ( .A(n_591), .Y(n_628) );
AND2x2_ASAP7_75t_L g661 ( .A(n_591), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g666 ( .A(n_591), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_591), .B(n_630), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g765 ( .A(n_591), .B(n_766), .C(n_767), .Y(n_765) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVxp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_600), .B1(n_607), .B2(n_608), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g691 ( .A(n_598), .Y(n_691) );
AND2x2_ASAP7_75t_L g625 ( .A(n_599), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g647 ( .A(n_599), .B(n_620), .Y(n_647) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_599), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
INVx1_ASAP7_75t_L g658 ( .A(n_601), .Y(n_658) );
AND2x2_ASAP7_75t_L g611 ( .A(n_602), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g637 ( .A(n_602), .Y(n_637) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g700 ( .A(n_606), .B(n_652), .Y(n_700) );
INVx1_ASAP7_75t_L g758 ( .A(n_606), .Y(n_758) );
INVx1_ASAP7_75t_L g614 ( .A(n_608), .Y(n_614) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_609), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g745 ( .A(n_609), .B(n_652), .Y(n_745) );
AND2x2_ASAP7_75t_L g711 ( .A(n_611), .B(n_712), .Y(n_711) );
NAND2x1p5_ASAP7_75t_L g779 ( .A(n_611), .B(n_780), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B(n_624), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_616), .B(n_651), .Y(n_650) );
AND2x4_ASAP7_75t_L g672 ( .A(n_616), .B(n_621), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_616), .B(n_662), .Y(n_723) );
AND2x4_ASAP7_75t_SL g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_617), .B(n_680), .Y(n_710) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_617), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_619), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_645) );
AND2x2_ASAP7_75t_SL g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_620), .B(n_662), .Y(n_681) );
INVx1_ASAP7_75t_L g782 ( .A(n_620), .Y(n_782) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B(n_631), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_626), .B(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g763 ( .A(n_629), .Y(n_763) );
INVx4_ASAP7_75t_L g665 ( .A(n_630), .Y(n_665) );
INVxp33_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g693 ( .A(n_632), .B(n_694), .Y(n_693) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_634), .B(n_649), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .B(n_645), .Y(n_634) );
INVx1_ASAP7_75t_L g683 ( .A(n_636), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_643), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g688 ( .A(n_640), .Y(n_688) );
INVx1_ASAP7_75t_L g721 ( .A(n_641), .Y(n_721) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_646), .A2(n_685), .B1(n_686), .B2(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g698 ( .A(n_647), .Y(n_698) );
NAND4xp25_ASAP7_75t_SL g649 ( .A(n_650), .B(n_656), .C(n_663), .D(n_669), .Y(n_649) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g671 ( .A(n_652), .Y(n_671) );
AND2x2_ASAP7_75t_L g783 ( .A(n_652), .B(n_780), .Y(n_783) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_661), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g790 ( .A(n_660), .B(n_727), .Y(n_790) );
INVx1_ASAP7_75t_L g787 ( .A(n_661), .Y(n_787) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_662), .Y(n_696) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B(n_668), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_701), .Y(n_673) );
NOR3xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_689), .C(n_697), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_682), .B(n_684), .Y(n_675) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_679), .A2(n_711), .B1(n_714), .B2(n_716), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_682), .A2(n_690), .B1(n_693), .B2(n_695), .Y(n_689) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g694 ( .A(n_687), .Y(n_694) );
AND2x4_ASAP7_75t_L g705 ( .A(n_687), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_692), .Y(n_792) );
AOI31xp33_ASAP7_75t_L g791 ( .A1(n_695), .A2(n_768), .A3(n_792), .B(n_793), .Y(n_791) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_717), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_703), .B(n_713), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_708), .B2(n_711), .Y(n_703) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_707), .Y(n_771) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_715), .B(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_718), .B(n_728), .Y(n_717) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
AND2x2_ASAP7_75t_L g729 ( .A(n_720), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g768 ( .A(n_720), .Y(n_768) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_720), .A2(n_778), .B1(n_781), .B2(n_783), .Y(n_777) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_725), .B(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B1(n_735), .B2(n_739), .Y(n_728) );
NOR2xp33_ASAP7_75t_SL g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVxp67_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
OR2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
INVx2_ASAP7_75t_SL g780 ( .A(n_737), .Y(n_780) );
INVx2_ASAP7_75t_L g761 ( .A(n_738), .Y(n_761) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_775), .Y(n_740) );
AOI211xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_747), .B(n_750), .C(n_764), .Y(n_741) );
OAI21xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B(n_746), .Y(n_742) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g749 ( .A(n_746), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_751), .B(n_755), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B1(n_760), .B2(n_762), .Y(n_755) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
AND2x2_ASAP7_75t_L g760 ( .A(n_758), .B(n_761), .Y(n_760) );
AO22x1_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_768), .B1(n_769), .B2(n_773), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NOR3xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_786), .C(n_791), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_777), .B(n_784), .Y(n_776) );
INVx3_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AOI21xp33_ASAP7_75t_R g786 ( .A1(n_787), .A2(n_788), .B(n_790), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_795), .Y(n_813) );
CKINVDCx11_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
CKINVDCx11_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_798), .Y(n_817) );
INVxp33_ASAP7_75t_L g818 ( .A(n_799), .Y(n_818) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx1_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g810 ( .A(n_811), .B(n_818), .Y(n_810) );
OAI22x1_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_813), .B1(n_814), .B2(n_815), .Y(n_811) );
CKINVDCx11_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
INVx3_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
BUFx4f_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_824), .Y(n_820) );
INVxp67_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_SL g827 ( .A(n_828), .Y(n_827) );
CKINVDCx11_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
CKINVDCx8_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
endmodule