module fake_netlist_1_6177_n_689 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_689);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_689;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_627;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_54), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_19), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_66), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_60), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_73), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_49), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_0), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_35), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_57), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_3), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_37), .Y(n_87) );
INVx3_ASAP7_75t_L g88 ( .A(n_21), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_44), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_72), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_33), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_50), .Y(n_92) );
BUFx3_ASAP7_75t_L g93 ( .A(n_7), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_13), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_58), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_74), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_68), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_5), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_38), .Y(n_99) );
NOR2xp67_ASAP7_75t_L g100 ( .A(n_3), .B(n_8), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_34), .Y(n_101) );
NOR2xp67_ASAP7_75t_L g102 ( .A(n_29), .B(n_26), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_5), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_64), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_76), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_24), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_62), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_6), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_23), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_15), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_56), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_47), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_75), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_25), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_12), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_69), .Y(n_117) );
INVxp33_ASAP7_75t_L g118 ( .A(n_48), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_36), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_12), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_11), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_7), .Y(n_122) );
BUFx10_ASAP7_75t_L g123 ( .A(n_32), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_123), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_121), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_88), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_104), .B(n_0), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_88), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_123), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_104), .B(n_1), .Y(n_132) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_78), .A2(n_31), .B(n_70), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_80), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g135 ( .A1(n_108), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_80), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_97), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_81), .B(n_39), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_85), .B(n_2), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_81), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_89), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_97), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_89), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_123), .Y(n_146) );
NAND2xp33_ASAP7_75t_R g147 ( .A(n_113), .B(n_40), .Y(n_147) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_90), .A2(n_30), .B(n_67), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_77), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_93), .B(n_4), .Y(n_150) );
INVx2_ASAP7_75t_SL g151 ( .A(n_95), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_95), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_99), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_99), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_101), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_105), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_105), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_86), .B(n_6), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_116), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_86), .B(n_8), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g161 ( .A1(n_83), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_161) );
CKINVDCx16_ASAP7_75t_R g162 ( .A(n_109), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_106), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_106), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_150), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_124), .B(n_107), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_127), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_124), .B(n_82), .Y(n_169) );
AO22x2_ASAP7_75t_L g170 ( .A1(n_150), .A2(n_117), .B1(n_119), .B2(n_120), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_150), .A2(n_103), .B1(n_120), .B2(n_94), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_124), .B(n_118), .Y(n_172) );
INVx5_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_128), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_127), .Y(n_176) );
INVx1_ASAP7_75t_SL g177 ( .A(n_125), .Y(n_177) );
INVx1_ASAP7_75t_SL g178 ( .A(n_155), .Y(n_178) );
OR2x6_ASAP7_75t_L g179 ( .A(n_161), .B(n_100), .Y(n_179) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_128), .B(n_117), .Y(n_180) );
NAND3xp33_ASAP7_75t_L g181 ( .A(n_132), .B(n_122), .C(n_111), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_127), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_124), .B(n_84), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_132), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_131), .B(n_98), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_131), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_127), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_127), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_129), .Y(n_192) );
OR2x2_ASAP7_75t_L g193 ( .A(n_139), .B(n_122), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_127), .Y(n_195) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_162), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_152), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_130), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_131), .B(n_103), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_131), .B(n_79), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_139), .B(n_111), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_130), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_130), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_146), .B(n_94), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_146), .B(n_116), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_146), .B(n_110), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_146), .B(n_87), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_129), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_162), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_130), .Y(n_211) );
NAND2x1_ASAP7_75t_L g212 ( .A(n_138), .B(n_119), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_130), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_130), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_152), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_129), .Y(n_216) );
OR2x2_ASAP7_75t_L g217 ( .A(n_164), .B(n_110), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_144), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_152), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_149), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_137), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_126), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_144), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_126), .B(n_96), .Y(n_224) );
OR2x2_ASAP7_75t_SL g225 ( .A(n_148), .B(n_9), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_134), .B(n_115), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_198), .Y(n_227) );
OR2x6_ASAP7_75t_L g228 ( .A(n_180), .B(n_135), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_186), .Y(n_229) );
AND2x6_ASAP7_75t_SL g230 ( .A(n_179), .B(n_158), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_199), .Y(n_231) );
INVxp33_ASAP7_75t_L g232 ( .A(n_187), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_198), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_222), .Y(n_234) );
OR2x2_ASAP7_75t_L g235 ( .A(n_193), .B(n_160), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_206), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_180), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_171), .A2(n_143), .B1(n_163), .B2(n_134), .Y(n_238) );
NOR2x2_ASAP7_75t_L g239 ( .A(n_179), .B(n_135), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_166), .B(n_136), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_170), .A2(n_161), .B1(n_147), .B2(n_151), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_174), .B(n_151), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_180), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_170), .A2(n_151), .B1(n_164), .B2(n_136), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_170), .A2(n_138), .B1(n_141), .B2(n_163), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_206), .Y(n_246) );
INVx1_ASAP7_75t_SL g247 ( .A(n_174), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_175), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_220), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_184), .B(n_141), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_221), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_170), .A2(n_143), .B1(n_140), .B2(n_157), .Y(n_252) );
BUFx8_ASAP7_75t_L g253 ( .A(n_182), .Y(n_253) );
INVx1_ASAP7_75t_SL g254 ( .A(n_193), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_224), .B(n_140), .Y(n_255) );
INVx4_ASAP7_75t_L g256 ( .A(n_175), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_168), .B(n_160), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_199), .Y(n_258) );
AND2x4_ASAP7_75t_SL g259 ( .A(n_210), .B(n_157), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_168), .B(n_158), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_199), .B(n_159), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_204), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_201), .A2(n_144), .B(n_156), .C(n_154), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_221), .Y(n_264) );
BUFx4f_ASAP7_75t_L g265 ( .A(n_204), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_224), .B(n_138), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_204), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_201), .B(n_138), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_175), .B(n_138), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_169), .B(n_156), .Y(n_270) );
NAND2x1p5_ASAP7_75t_L g271 ( .A(n_217), .B(n_159), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_188), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_172), .A2(n_156), .B1(n_154), .B2(n_153), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_207), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_218), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_188), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_181), .A2(n_154), .B1(n_153), .B2(n_142), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_207), .B(n_153), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_192), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_217), .Y(n_280) );
AND2x6_ASAP7_75t_L g281 ( .A(n_165), .B(n_142), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_168), .B(n_159), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_205), .A2(n_142), .B1(n_137), .B2(n_159), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_226), .B(n_137), .Y(n_284) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_179), .A2(n_148), .B1(n_133), .B2(n_114), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_179), .A2(n_112), .B1(n_92), .B2(n_91), .Y(n_286) );
AO22x1_ASAP7_75t_L g287 ( .A1(n_220), .A2(n_177), .B1(n_178), .B2(n_205), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_205), .A2(n_148), .B1(n_133), .B2(n_102), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_173), .B(n_148), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_209), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_216), .Y(n_291) );
NOR2xp33_ASAP7_75t_SL g292 ( .A(n_249), .B(n_196), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_254), .B(n_208), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_254), .B(n_235), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_275), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_278), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_253), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_237), .A2(n_225), .B1(n_200), .B2(n_212), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_278), .Y(n_299) );
INVx2_ASAP7_75t_SL g300 ( .A(n_265), .Y(n_300) );
AND2x2_ASAP7_75t_SL g301 ( .A(n_245), .B(n_148), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_247), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_253), .Y(n_304) );
BUFx12f_ASAP7_75t_L g305 ( .A(n_230), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_263), .A2(n_212), .B(n_223), .C(n_173), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_280), .B(n_173), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_244), .A2(n_173), .B1(n_210), .B2(n_133), .Y(n_308) );
AND2x6_ASAP7_75t_L g309 ( .A(n_252), .B(n_231), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_251), .Y(n_310) );
OAI22xp5_ASAP7_75t_SL g311 ( .A1(n_228), .A2(n_225), .B1(n_133), .B2(n_173), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_290), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_271), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_232), .B(n_202), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_264), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_247), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_291), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_243), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_269), .A2(n_195), .B(n_214), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_279), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_248), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_248), .Y(n_322) );
INVxp67_ASAP7_75t_SL g323 ( .A(n_265), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_258), .Y(n_324) );
O2A1O1Ixp33_ASAP7_75t_SL g325 ( .A1(n_285), .A2(n_185), .B(n_195), .C(n_214), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_256), .Y(n_326) );
NAND2x1_ASAP7_75t_SL g327 ( .A(n_241), .B(n_215), .Y(n_327) );
OR2x6_ASAP7_75t_L g328 ( .A(n_228), .B(n_167), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_256), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_289), .A2(n_213), .B(n_211), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_227), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_259), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_263), .A2(n_215), .B(n_190), .C(n_194), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_234), .A2(n_267), .B1(n_229), .B2(n_274), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_242), .B(n_202), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_268), .A2(n_211), .B1(n_213), .B2(n_185), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_267), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_242), .B(n_197), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_281), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_282), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_310), .Y(n_342) );
OA21x2_ASAP7_75t_L g343 ( .A1(n_330), .A2(n_288), .B(n_269), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_296), .B(n_268), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_294), .A2(n_228), .B1(n_236), .B2(n_246), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_301), .A2(n_285), .B(n_266), .Y(n_347) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_294), .A2(n_239), .B1(n_238), .B2(n_255), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_298), .A2(n_284), .B(n_238), .C(n_270), .Y(n_349) );
INVx4_ASAP7_75t_L g350 ( .A(n_295), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_310), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_301), .A2(n_266), .B(n_260), .Y(n_352) );
AOI21x1_ASAP7_75t_L g353 ( .A1(n_330), .A2(n_284), .B(n_219), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_308), .B(n_273), .C(n_287), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_301), .A2(n_257), .B(n_283), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_309), .A2(n_250), .B1(n_240), .B2(n_261), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_316), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_332), .B(n_286), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_296), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_327), .A2(n_277), .B(n_276), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_299), .B(n_255), .Y(n_361) );
AO21x2_ASAP7_75t_L g362 ( .A1(n_325), .A2(n_219), .B(n_272), .Y(n_362) );
OA21x2_ASAP7_75t_L g363 ( .A1(n_308), .A2(n_233), .B(n_282), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_309), .A2(n_261), .B1(n_281), .B2(n_276), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_299), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_302), .B(n_281), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_312), .B(n_281), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_311), .A2(n_190), .B(n_215), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_312), .B(n_281), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_315), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_332), .B(n_10), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_342), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_361), .B(n_293), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_361), .B(n_317), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_359), .B(n_293), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_358), .B(n_292), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g377 ( .A1(n_349), .A2(n_327), .B(n_333), .C(n_317), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g378 ( .A1(n_344), .A2(n_304), .B1(n_328), .B2(n_297), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_348), .A2(n_346), .B1(n_335), .B2(n_356), .C(n_344), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_348), .B(n_305), .Y(n_380) );
AO22x1_ASAP7_75t_L g381 ( .A1(n_347), .A2(n_304), .B1(n_309), .B2(n_313), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_371), .A2(n_334), .B1(n_341), .B2(n_300), .C(n_323), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_349), .A2(n_334), .B1(n_341), .B2(n_300), .C(n_307), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_359), .B(n_302), .Y(n_384) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_366), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_365), .B(n_313), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_365), .B(n_320), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_368), .A2(n_319), .B(n_306), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_357), .A2(n_309), .B1(n_328), .B2(n_305), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_342), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_357), .A2(n_309), .B1(n_328), .B2(n_340), .Y(n_391) );
OAI21xp33_ASAP7_75t_L g392 ( .A1(n_354), .A2(n_328), .B(n_320), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_345), .B(n_315), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_356), .B(n_324), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_366), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_351), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_374), .B(n_351), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_374), .B(n_347), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_395), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_385), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_393), .B(n_345), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_387), .B(n_370), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_385), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_397), .B(n_350), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_398), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_372), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_372), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_387), .B(n_370), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_397), .B(n_350), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_393), .B(n_370), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_390), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_395), .B(n_369), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
NOR2x1_ASAP7_75t_R g417 ( .A(n_385), .B(n_350), .Y(n_417) );
NOR2x1_ASAP7_75t_L g418 ( .A(n_396), .B(n_350), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_397), .B(n_369), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_396), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_384), .B(n_369), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_379), .A2(n_309), .B1(n_363), .B2(n_354), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_380), .A2(n_309), .B1(n_363), .B2(n_364), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_390), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_384), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_373), .B(n_363), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_375), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_375), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_394), .B(n_363), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_386), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_377), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_389), .B(n_363), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_381), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_407), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_414), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_428), .B(n_376), .Y(n_437) );
BUFx12f_ASAP7_75t_L g438 ( .A(n_402), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_401), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_413), .B(n_391), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_408), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_408), .B(n_429), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_399), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_428), .B(n_378), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_429), .B(n_392), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_414), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_422), .A2(n_366), .B(n_382), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_401), .Y(n_448) );
AOI33xp33_ASAP7_75t_L g449 ( .A1(n_423), .A2(n_383), .A3(n_366), .B1(n_307), .B2(n_17), .B3(n_16), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_402), .B(n_392), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_399), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_420), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_413), .B(n_352), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_404), .B(n_352), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_420), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_422), .A2(n_368), .B(n_388), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_404), .B(n_411), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_402), .B(n_295), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_432), .A2(n_355), .B1(n_367), .B2(n_295), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_424), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_424), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_407), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_409), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_411), .B(n_362), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_427), .A2(n_324), .B1(n_367), .B2(n_314), .C(n_355), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_427), .B(n_318), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_417), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_432), .A2(n_295), .B1(n_340), .B2(n_318), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_427), .B(n_318), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_418), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_409), .Y(n_473) );
INVx4_ASAP7_75t_L g474 ( .A(n_405), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_425), .A2(n_295), .B1(n_318), .B2(n_338), .Y(n_475) );
AOI21xp33_ASAP7_75t_L g476 ( .A1(n_417), .A2(n_362), .B(n_360), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_430), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_403), .A2(n_318), .B1(n_321), .B2(n_326), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_426), .B(n_362), .Y(n_479) );
OAI222xp33_ASAP7_75t_L g480 ( .A1(n_434), .A2(n_353), .B1(n_321), .B2(n_326), .C1(n_17), .C2(n_16), .Y(n_480) );
INVxp67_ASAP7_75t_SL g481 ( .A(n_409), .Y(n_481) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_426), .A2(n_353), .B(n_362), .Y(n_482) );
NOR2xp67_ASAP7_75t_L g483 ( .A(n_433), .B(n_14), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_403), .B(n_343), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_400), .B(n_343), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_439), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_439), .B(n_434), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_435), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_448), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_458), .B(n_433), .Y(n_490) );
AND3x1_ASAP7_75t_L g491 ( .A(n_437), .B(n_433), .C(n_421), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_442), .B(n_441), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_458), .B(n_410), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_443), .B(n_430), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_438), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_466), .B(n_410), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_441), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_442), .B(n_410), .Y(n_498) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_474), .B(n_405), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_466), .B(n_416), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_448), .B(n_416), .Y(n_501) );
NAND4xp25_ASAP7_75t_L g502 ( .A(n_449), .B(n_421), .C(n_400), .D(n_405), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_452), .B(n_416), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_435), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_452), .B(n_415), .Y(n_505) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_474), .B(n_430), .Y(n_506) );
NOR2x1_ASAP7_75t_SL g507 ( .A(n_438), .B(n_425), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_474), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_451), .B(n_425), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_444), .B(n_415), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_436), .B(n_425), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_455), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_455), .B(n_425), .Y(n_513) );
AOI221x1_ASAP7_75t_L g514 ( .A1(n_476), .A2(n_412), .B1(n_406), .B2(n_431), .C(n_419), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g515 ( .A(n_447), .B(n_419), .C(n_406), .D(n_412), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_481), .B(n_425), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_464), .B(n_431), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_464), .B(n_431), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_456), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_436), .B(n_419), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_465), .B(n_431), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_446), .B(n_419), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_446), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_465), .B(n_431), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_462), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_477), .B(n_431), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_462), .B(n_412), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_469), .A2(n_412), .B1(n_406), .B2(n_341), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_463), .B(n_406), .Y(n_529) );
NAND2x1p5_ASAP7_75t_SL g530 ( .A(n_450), .B(n_331), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_463), .B(n_14), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_456), .B(n_343), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_454), .B(n_15), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_460), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_445), .B(n_343), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_440), .B(n_338), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_473), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_473), .B(n_343), .Y(n_538) );
AOI211x1_ASAP7_75t_L g539 ( .A1(n_480), .A2(n_336), .B(n_339), .C(n_337), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_468), .Y(n_540) );
NAND2xp33_ASAP7_75t_SL g541 ( .A(n_460), .B(n_329), .Y(n_541) );
AND2x4_ASAP7_75t_SL g542 ( .A(n_440), .B(n_322), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_459), .B(n_472), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_482), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_505), .B(n_484), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_505), .B(n_479), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_525), .B(n_479), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_495), .B(n_472), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_486), .B(n_445), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_493), .B(n_454), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_489), .B(n_485), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_512), .B(n_485), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_492), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_493), .Y(n_555) );
NOR2xp67_ASAP7_75t_L g556 ( .A(n_515), .B(n_483), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_494), .B(n_471), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_498), .B(n_453), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_497), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_487), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_487), .Y(n_561) );
NAND3xp33_ASAP7_75t_L g562 ( .A(n_534), .B(n_457), .C(n_470), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_487), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_510), .B(n_453), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_508), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_490), .B(n_461), .Y(n_566) );
NAND4xp25_ASAP7_75t_L g567 ( .A(n_502), .B(n_467), .C(n_478), .D(n_475), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_529), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_508), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_490), .B(n_482), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_529), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_540), .B(n_482), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_527), .B(n_360), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_527), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_498), .B(n_360), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_523), .B(n_18), .Y(n_576) );
NAND2x1p5_ASAP7_75t_L g577 ( .A(n_499), .B(n_329), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_496), .B(n_20), .Y(n_578) );
NAND3xp33_ASAP7_75t_SL g579 ( .A(n_531), .B(n_322), .C(n_331), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_506), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_496), .B(n_22), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_501), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_509), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_501), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_503), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_500), .B(n_27), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_503), .B(n_203), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_531), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_500), .B(n_203), .Y(n_589) );
XNOR2x2_ASAP7_75t_L g590 ( .A(n_543), .B(n_28), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_509), .B(n_41), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_523), .B(n_203), .Y(n_592) );
INVx2_ASAP7_75t_SL g593 ( .A(n_520), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_513), .B(n_203), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_513), .B(n_203), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_536), .A2(n_189), .B1(n_176), .B2(n_191), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_588), .A2(n_491), .B1(n_533), .B2(n_539), .C(n_526), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_551), .B(n_542), .Y(n_598) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_579), .B(n_522), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_546), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_554), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_555), .B(n_520), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_568), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_593), .B(n_542), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_571), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_562), .B(n_514), .C(n_544), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_574), .Y(n_607) );
AOI31xp33_ASAP7_75t_L g608 ( .A1(n_565), .A2(n_541), .A3(n_522), .B(n_528), .Y(n_608) );
OAI211xp5_ASAP7_75t_L g609 ( .A1(n_556), .A2(n_541), .B(n_511), .C(n_535), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_558), .B(n_511), .Y(n_610) );
NAND3xp33_ASAP7_75t_SL g611 ( .A(n_577), .B(n_530), .C(n_516), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_569), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_567), .A2(n_526), .B1(n_517), .B2(n_518), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_577), .A2(n_516), .B1(n_504), .B2(n_537), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_559), .B(n_521), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_582), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_550), .B(n_518), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_584), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_549), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_576), .A2(n_507), .B(n_521), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_560), .A2(n_517), .B(n_524), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_585), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_561), .B(n_524), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_550), .B(n_544), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g625 ( .A1(n_563), .A2(n_535), .B(n_537), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_583), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_557), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_547), .B(n_519), .Y(n_628) );
OAI21xp33_ASAP7_75t_SL g629 ( .A1(n_580), .A2(n_519), .B(n_504), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_547), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_576), .A2(n_488), .B(n_530), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_570), .B(n_488), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_608), .A2(n_572), .B(n_548), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_617), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_608), .A2(n_545), .B1(n_564), .B2(n_566), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_630), .B(n_545), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_597), .A2(n_548), .B1(n_553), .B2(n_552), .C(n_589), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_619), .B(n_553), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_617), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_627), .B(n_552), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_628), .Y(n_641) );
OAI21xp33_ASAP7_75t_L g642 ( .A1(n_613), .A2(n_573), .B(n_589), .Y(n_642) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_606), .A2(n_591), .B(n_595), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_616), .Y(n_644) );
AO22x2_ASAP7_75t_L g645 ( .A1(n_600), .A2(n_575), .B1(n_586), .B2(n_578), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_612), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_618), .B(n_595), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_622), .B(n_594), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_607), .Y(n_649) );
OAI321xp33_ASAP7_75t_L g650 ( .A1(n_609), .A2(n_581), .A3(n_596), .B1(n_590), .B2(n_594), .C(n_592), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_610), .Y(n_651) );
INVx1_ASAP7_75t_SL g652 ( .A(n_598), .Y(n_652) );
NAND4xp25_ASAP7_75t_SL g653 ( .A(n_629), .B(n_592), .C(n_587), .D(n_538), .Y(n_653) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_611), .B(n_587), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_635), .A2(n_597), .B(n_601), .C(n_599), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_637), .A2(n_631), .B(n_614), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_638), .A2(n_603), .B1(n_605), .B2(n_625), .C(n_621), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_634), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_653), .A2(n_624), .B1(n_614), .B2(n_615), .C(n_623), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g660 ( .A(n_652), .Y(n_660) );
AOI322xp5_ASAP7_75t_L g661 ( .A1(n_640), .A2(n_632), .A3(n_623), .B1(n_626), .B2(n_604), .C1(n_624), .C2(n_538), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_639), .B(n_602), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_645), .A2(n_620), .B1(n_631), .B2(n_532), .Y(n_663) );
AOI221xp5_ASAP7_75t_SL g664 ( .A1(n_633), .A2(n_532), .B1(n_167), .B2(n_191), .C(n_189), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_650), .A2(n_197), .B(n_194), .Y(n_665) );
A2O1A1Ixp33_ASAP7_75t_SL g666 ( .A1(n_643), .A2(n_197), .B(n_194), .C(n_190), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_644), .Y(n_667) );
XNOR2x1_ASAP7_75t_L g668 ( .A(n_660), .B(n_645), .Y(n_668) );
NOR4xp25_ASAP7_75t_L g669 ( .A(n_655), .B(n_642), .C(n_646), .D(n_649), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_656), .A2(n_641), .B1(n_651), .B2(n_648), .C(n_647), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_667), .B(n_646), .Y(n_671) );
O2A1O1Ixp5_ASAP7_75t_L g672 ( .A1(n_658), .A2(n_636), .B(n_654), .C(n_45), .Y(n_672) );
OAI211xp5_ASAP7_75t_SL g673 ( .A1(n_663), .A2(n_42), .B(n_43), .C(n_46), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_667), .B(n_51), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_659), .A2(n_191), .B1(n_189), .B2(n_183), .C(n_176), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_671), .Y(n_676) );
NAND5xp2_ASAP7_75t_L g677 ( .A(n_675), .B(n_664), .C(n_661), .D(n_657), .E(n_665), .Y(n_677) );
OAI21xp33_ASAP7_75t_SL g678 ( .A1(n_669), .A2(n_662), .B(n_666), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g679 ( .A(n_672), .B(n_52), .C(n_53), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_678), .A2(n_668), .B1(n_670), .B2(n_673), .C(n_674), .Y(n_680) );
OA22x2_ASAP7_75t_SL g681 ( .A1(n_676), .A2(n_55), .B1(n_59), .B2(n_61), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_679), .B(n_176), .C(n_189), .Y(n_682) );
OA22x2_ASAP7_75t_L g683 ( .A1(n_680), .A2(n_677), .B1(n_65), .B2(n_71), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_682), .A2(n_681), .B1(n_167), .B2(n_176), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_683), .A2(n_167), .B1(n_176), .B2(n_183), .C(n_189), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_685), .Y(n_686) );
XNOR2xp5_ASAP7_75t_L g687 ( .A(n_686), .B(n_684), .Y(n_687) );
AOI22x1_ASAP7_75t_L g688 ( .A1(n_687), .A2(n_167), .B1(n_183), .B2(n_191), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_688), .A2(n_63), .B1(n_183), .B2(n_191), .C(n_680), .Y(n_689) );
endmodule