module real_aes_9931_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g150 ( .A(n_0), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g510 ( .A(n_1), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_2), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_3), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_4), .B(n_529), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_5), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_6), .B(n_180), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_7), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_8), .B(n_143), .Y(n_142) );
NOR2xp67_ASAP7_75t_L g107 ( .A(n_9), .B(n_91), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_10), .B(n_136), .Y(n_213) );
INVx1_ASAP7_75t_L g862 ( .A(n_11), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_11), .B(n_863), .Y(n_870) );
AOI21xp33_ASAP7_75t_SL g873 ( .A1(n_12), .A2(n_871), .B(n_874), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_13), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_14), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_15), .B(n_143), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_16), .B(n_199), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_17), .B(n_267), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_18), .B(n_161), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_19), .B(n_143), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_20), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_21), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_22), .B(n_136), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_23), .B(n_180), .Y(n_197) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_24), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_25), .B(n_199), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_26), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_27), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_28), .B(n_199), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_29), .B(n_161), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_30), .A2(n_94), .B1(n_859), .B2(n_860), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_30), .Y(n_859) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_31), .Y(n_137) );
OAI21xp33_ASAP7_75t_L g547 ( .A1(n_32), .A2(n_147), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_33), .B(n_136), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_34), .B(n_215), .Y(n_263) );
NAND2xp33_ASAP7_75t_SL g248 ( .A(n_35), .B(n_186), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_36), .B(n_136), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_37), .B(n_202), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_38), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_39), .B(n_139), .Y(n_217) );
INVx1_ASAP7_75t_L g112 ( .A(n_40), .Y(n_112) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_41), .A2(n_74), .B(n_130), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g872 ( .A(n_42), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_43), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_44), .B(n_136), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_45), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_46), .B(n_202), .Y(n_201) );
AND2x6_ASAP7_75t_L g148 ( .A(n_47), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_48), .B(n_172), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_49), .A2(n_87), .B1(n_529), .B2(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_50), .B(n_172), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_51), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_52), .B(n_127), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_53), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_54), .A2(n_843), .B1(n_846), .B2(n_847), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_54), .Y(n_847) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_55), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_56), .A2(n_101), .B1(n_844), .B2(n_845), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_56), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_57), .Y(n_530) );
INVx1_ASAP7_75t_L g149 ( .A(n_58), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_59), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_60), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_61), .B(n_550), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_62), .B(n_550), .Y(n_562) );
NAND2xp33_ASAP7_75t_L g246 ( .A(n_63), .B(n_186), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_64), .B(n_202), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_65), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_66), .B(n_127), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_67), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g879 ( .A(n_68), .Y(n_879) );
AND2x2_ASAP7_75t_L g110 ( .A(n_69), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g520 ( .A(n_70), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_71), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_72), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_73), .B(n_167), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_75), .B(n_136), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_76), .B(n_143), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_77), .B(n_161), .Y(n_195) );
INVx1_ASAP7_75t_L g514 ( .A(n_78), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_79), .B(n_202), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_80), .Y(n_614) );
BUFx10_ASAP7_75t_L g851 ( .A(n_81), .Y(n_851) );
INVx1_ASAP7_75t_L g608 ( .A(n_82), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_83), .B(n_143), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_84), .B(n_136), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_85), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_86), .B(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_88), .B(n_127), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_89), .B(n_143), .Y(n_194) );
INVx1_ASAP7_75t_L g523 ( .A(n_90), .Y(n_523) );
INVx2_ASAP7_75t_L g130 ( .A(n_92), .Y(n_130) );
INVx1_ASAP7_75t_L g113 ( .A(n_93), .Y(n_113) );
BUFx2_ASAP7_75t_L g483 ( .A(n_93), .Y(n_483) );
OR2x2_ASAP7_75t_L g867 ( .A(n_93), .B(n_868), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_93), .B(n_852), .Y(n_877) );
INVx1_ASAP7_75t_L g860 ( .A(n_94), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_95), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_96), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g111 ( .A(n_97), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_98), .B(n_180), .Y(n_187) );
NOR2xp67_ASAP7_75t_L g544 ( .A(n_99), .B(n_545), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_100), .Y(n_230) );
INVx1_ASAP7_75t_L g844 ( .A(n_101), .Y(n_844) );
NAND2xp33_ASAP7_75t_L g569 ( .A(n_102), .B(n_127), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_114), .B(n_878), .Y(n_103) );
INVx4_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx6_ASAP7_75t_L g880 ( .A(n_105), .Y(n_880) );
INVx6_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x4_ASAP7_75t_L g852 ( .A(n_107), .B(n_112), .Y(n_852) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .C(n_113), .Y(n_108) );
INVx4_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_848), .B(n_853), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
XNOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_842), .Y(n_117) );
OAI22x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_482), .B1(n_484), .B2(n_841), .Y(n_118) );
XNOR2xp5_ASAP7_75t_L g857 ( .A(n_119), .B(n_858), .Y(n_857) );
NAND3x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_357), .C(n_436), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_310), .Y(n_120) );
AOI211xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_204), .B(n_251), .C(n_301), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_153), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_124), .B(n_278), .Y(n_411) );
AND2x2_ASAP7_75t_L g442 ( .A(n_124), .B(n_174), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_124), .B(n_331), .Y(n_445) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2x1_ASAP7_75t_L g277 ( .A(n_125), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g329 ( .A(n_125), .B(n_290), .Y(n_329) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g254 ( .A(n_126), .B(n_176), .Y(n_254) );
INVx3_ASAP7_75t_L g289 ( .A(n_126), .Y(n_289) );
AND2x2_ASAP7_75t_L g309 ( .A(n_126), .B(n_155), .Y(n_309) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_131), .B(n_150), .Y(n_126) );
OAI21x1_ASAP7_75t_L g210 ( .A1(n_127), .A2(n_211), .B(n_220), .Y(n_210) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_127), .A2(n_224), .B(n_233), .Y(n_223) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_127), .A2(n_261), .B(n_269), .Y(n_260) );
INVx2_ASAP7_75t_L g542 ( .A(n_127), .Y(n_542) );
NOR2x1p5_ASAP7_75t_SL g578 ( .A(n_127), .B(n_579), .Y(n_578) );
BUFx5_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g173 ( .A(n_128), .Y(n_173) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_128), .Y(n_270) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g152 ( .A(n_129), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_135), .B(n_141), .C(n_148), .Y(n_131) );
AOI21x1_ASAP7_75t_L g163 ( .A1(n_132), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_132), .A2(n_248), .B(n_249), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_132), .A2(n_266), .B(n_268), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_132), .A2(n_500), .B(n_501), .Y(n_499) );
INVx2_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_133), .A2(n_160), .B(n_162), .Y(n_159) );
INVx2_ASAP7_75t_SL g200 ( .A(n_133), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_133), .A2(n_244), .B(n_245), .C(n_246), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_133), .A2(n_263), .B(n_264), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_133), .A2(n_497), .B(n_498), .Y(n_496) );
CKINVDCx6p67_ASAP7_75t_R g563 ( .A(n_133), .Y(n_563) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx12f_ASAP7_75t_L g147 ( .A(n_134), .Y(n_147) );
INVx5_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_138), .B1(n_139), .B2(n_140), .Y(n_135) );
INVx2_ASAP7_75t_L g512 ( .A(n_136), .Y(n_512) );
INVx2_ASAP7_75t_L g590 ( .A(n_136), .Y(n_590) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g139 ( .A(n_137), .Y(n_139) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_137), .Y(n_146) );
INVx1_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_137), .Y(n_186) );
INVx1_ASAP7_75t_L g245 ( .A(n_139), .Y(n_245) );
INVx2_ASAP7_75t_L g267 ( .A(n_139), .Y(n_267) );
INVx2_ASAP7_75t_L g529 ( .A(n_139), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_144), .B(n_147), .Y(n_141) );
INVx5_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
OR2x2_ASAP7_75t_L g610 ( .A(n_143), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g231 ( .A(n_145), .Y(n_231) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g199 ( .A(n_146), .Y(n_199) );
INVx2_ASAP7_75t_L g215 ( .A(n_146), .Y(n_215) );
INVx2_ASAP7_75t_L g227 ( .A(n_146), .Y(n_227) );
INVx2_ASAP7_75t_L g531 ( .A(n_146), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_147), .A2(n_184), .B(n_187), .Y(n_183) );
BUFx2_ASAP7_75t_L g515 ( .A(n_147), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_147), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_147), .B(n_536), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_147), .A2(n_544), .B1(n_547), .B2(n_549), .Y(n_543) );
INVx3_ASAP7_75t_L g591 ( .A(n_147), .Y(n_591) );
INVx8_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
OAI21x1_ASAP7_75t_SL g177 ( .A1(n_148), .A2(n_178), .B(n_183), .Y(n_177) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_148), .A2(n_193), .B(n_196), .Y(n_192) );
AOI21xp33_ASAP7_75t_L g524 ( .A1(n_148), .A2(n_203), .B(n_522), .Y(n_524) );
INVx1_ASAP7_75t_L g534 ( .A(n_148), .Y(n_534) );
INVx1_ASAP7_75t_L g579 ( .A(n_148), .Y(n_579) );
BUFx4f_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
OAI21x1_ASAP7_75t_L g176 ( .A1(n_151), .A2(n_177), .B(n_188), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_151), .B(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g558 ( .A(n_151), .Y(n_558) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
INVx2_ASAP7_75t_L g420 ( .A(n_153), .Y(n_420) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_174), .Y(n_153) );
AND2x2_ASAP7_75t_L g253 ( .A(n_154), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g345 ( .A(n_154), .Y(n_345) );
AND2x2_ASAP7_75t_L g441 ( .A(n_154), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g278 ( .A(n_155), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g288 ( .A(n_155), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVxp67_ASAP7_75t_R g339 ( .A(n_156), .Y(n_339) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_171), .Y(n_156) );
OAI21xp5_ASAP7_75t_L g323 ( .A1(n_157), .A2(n_158), .B(n_171), .Y(n_323) );
OAI21x1_ASAP7_75t_L g494 ( .A1(n_157), .A2(n_495), .B(n_502), .Y(n_494) );
OAI21x1_ASAP7_75t_SL g585 ( .A1(n_157), .A2(n_586), .B(n_596), .Y(n_585) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_163), .B(n_169), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_161), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_161), .A2(n_529), .B1(n_572), .B2(n_573), .Y(n_571) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g180 ( .A(n_168), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_169), .A2(n_225), .B(n_229), .Y(n_224) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_169), .A2(n_243), .B(n_247), .Y(n_242) );
OAI21x1_ASAP7_75t_L g495 ( .A1(n_169), .A2(n_496), .B(n_499), .Y(n_495) );
INVx2_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
INVx8_ASAP7_75t_L g219 ( .A(n_170), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g615 ( .A1(n_170), .A2(n_202), .B(n_616), .Y(n_615) );
OAI21x1_ASAP7_75t_L g191 ( .A1(n_172), .A2(n_192), .B(n_201), .Y(n_191) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_172), .A2(n_242), .B(n_250), .Y(n_241) );
INVx2_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g189 ( .A(n_173), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_173), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g338 ( .A(n_174), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_190), .Y(n_174) );
INVx2_ASAP7_75t_SL g291 ( .A(n_175), .Y(n_291) );
INVx1_ASAP7_75t_L g297 ( .A(n_175), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_175), .B(n_289), .Y(n_318) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_175), .Y(n_350) );
INVx1_ASAP7_75t_L g396 ( .A(n_175), .Y(n_396) );
AND2x2_ASAP7_75t_L g417 ( .A(n_175), .B(n_370), .Y(n_417) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_175), .Y(n_432) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .C(n_182), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_180), .A2(n_512), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_182), .A2(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_182), .A2(n_217), .B(n_218), .Y(n_216) );
O2A1O1Ixp5_ASAP7_75t_L g229 ( .A1(n_182), .A2(n_230), .B(n_231), .C(n_232), .Y(n_229) );
OAI21xp33_ASAP7_75t_L g527 ( .A1(n_182), .A2(n_528), .B(n_533), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_182), .A2(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g595 ( .A(n_182), .Y(n_595) );
INVx2_ASAP7_75t_L g518 ( .A(n_185), .Y(n_518) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g546 ( .A(n_186), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_186), .Y(n_548) );
INVx2_ASAP7_75t_L g550 ( .A(n_186), .Y(n_550) );
INVx1_ASAP7_75t_L g279 ( .A(n_190), .Y(n_279) );
AND2x2_ASAP7_75t_L g290 ( .A(n_190), .B(n_291), .Y(n_290) );
NOR2xp67_ASAP7_75t_L g296 ( .A(n_190), .B(n_297), .Y(n_296) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_190), .Y(n_308) );
AND2x2_ASAP7_75t_L g363 ( .A(n_190), .B(n_323), .Y(n_363) );
INVx1_ASAP7_75t_L g371 ( .A(n_190), .Y(n_371) );
INVx1_ASAP7_75t_L g433 ( .A(n_190), .Y(n_433) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g331 ( .A(n_191), .B(n_323), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_200), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_199), .B(n_514), .Y(n_513) );
INVxp67_ASAP7_75t_L g576 ( .A(n_199), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_199), .B(n_614), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_200), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_200), .A2(n_226), .B(n_228), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g574 ( .A1(n_200), .A2(n_575), .B(n_576), .C(n_577), .Y(n_574) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_203), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_203), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_234), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_206), .B(n_283), .Y(n_447) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g419 ( .A(n_207), .Y(n_419) );
OR2x2_ASAP7_75t_L g458 ( .A(n_207), .B(n_406), .Y(n_458) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g313 ( .A(n_208), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g390 ( .A(n_208), .B(n_342), .Y(n_390) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_221), .Y(n_208) );
INVx2_ASAP7_75t_L g276 ( .A(n_209), .Y(n_276) );
AND2x2_ASAP7_75t_L g282 ( .A(n_209), .B(n_222), .Y(n_282) );
INVx1_ASAP7_75t_L g294 ( .A(n_209), .Y(n_294) );
INVx1_ASAP7_75t_L g405 ( .A(n_209), .Y(n_405) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_216), .B(n_219), .Y(n_211) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_219), .A2(n_262), .B(n_265), .Y(n_261) );
AO31x2_ASAP7_75t_L g541 ( .A1(n_219), .A2(n_542), .A3(n_543), .B(n_551), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_219), .A2(n_560), .B(n_564), .Y(n_559) );
OAI21x1_ASAP7_75t_SL g586 ( .A1(n_219), .A2(n_587), .B(n_592), .Y(n_586) );
INVx1_ASAP7_75t_L g235 ( .A(n_221), .Y(n_235) );
AND2x2_ASAP7_75t_L g299 ( .A(n_221), .B(n_294), .Y(n_299) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_221), .Y(n_383) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g356 ( .A(n_222), .Y(n_356) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g271 ( .A(n_223), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
AND2x2_ASAP7_75t_L g460 ( .A(n_236), .B(n_392), .Y(n_460) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g304 ( .A(n_238), .Y(n_304) );
INVx1_ASAP7_75t_L g314 ( .A(n_238), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_238), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g300 ( .A(n_239), .B(n_259), .Y(n_300) );
AND2x2_ASAP7_75t_L g440 ( .A(n_239), .B(n_275), .Y(n_440) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g274 ( .A(n_240), .Y(n_274) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_240), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_240), .B(n_259), .Y(n_378) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g352 ( .A(n_241), .B(n_276), .Y(n_352) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_241), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_245), .A2(n_531), .B1(n_537), .B2(n_538), .Y(n_536) );
OAI221xp5_ASAP7_75t_SL g251 ( .A1(n_252), .A2(n_255), .B1(n_277), .B2(n_280), .C(n_286), .Y(n_251) );
OAI32xp33_ASAP7_75t_L g454 ( .A1(n_252), .A2(n_352), .A3(n_455), .B1(n_457), .B2(n_458), .Y(n_454) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g388 ( .A(n_254), .B(n_363), .Y(n_388) );
AND2x2_ASAP7_75t_L g392 ( .A(n_254), .B(n_284), .Y(n_392) );
INVx1_ASAP7_75t_L g479 ( .A(n_254), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_272), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_256), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g457 ( .A(n_256), .Y(n_457) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g360 ( .A(n_257), .B(n_326), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g257 ( .A(n_258), .B(n_271), .Y(n_257) );
BUFx2_ASAP7_75t_L g292 ( .A(n_258), .Y(n_292) );
INVx2_ASAP7_75t_L g335 ( .A(n_258), .Y(n_335) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g285 ( .A(n_260), .Y(n_285) );
INVx2_ASAP7_75t_L g401 ( .A(n_271), .Y(n_401) );
INVx1_ASAP7_75t_L g332 ( .A(n_272), .Y(n_332) );
AOI322xp5_ASAP7_75t_L g373 ( .A1(n_272), .A2(n_374), .A3(n_376), .B1(n_377), .B2(n_379), .C1(n_380), .C2(n_381), .Y(n_373) );
AND2x4_ASAP7_75t_SL g469 ( .A(n_272), .B(n_406), .Y(n_469) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g326 ( .A(n_274), .Y(n_326) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g456 ( .A(n_278), .Y(n_456) );
OAI221xp5_ASAP7_75t_L g336 ( .A1(n_280), .A2(n_337), .B1(n_340), .B2(n_343), .C(n_346), .Y(n_336) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g303 ( .A(n_282), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g372 ( .A(n_282), .B(n_326), .Y(n_372) );
INVx1_ASAP7_75t_L g475 ( .A(n_282), .Y(n_475) );
INVx1_ASAP7_75t_L g312 ( .A(n_283), .Y(n_312) );
AND2x2_ASAP7_75t_L g410 ( .A(n_283), .B(n_299), .Y(n_410) );
BUFx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_284), .B(n_356), .Y(n_375) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx3_ASAP7_75t_L g354 ( .A(n_285), .Y(n_354) );
AOI32xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_292), .A3(n_293), .B1(n_295), .B2(n_298), .Y(n_286) );
INVx1_ASAP7_75t_L g408 ( .A(n_287), .Y(n_408) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
AND2x4_ASAP7_75t_L g295 ( .A(n_288), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g434 ( .A(n_288), .Y(n_434) );
AND2x2_ASAP7_75t_L g365 ( .A(n_289), .B(n_291), .Y(n_365) );
INVx1_ASAP7_75t_L g370 ( .A(n_289), .Y(n_370) );
AND2x2_ASAP7_75t_L g481 ( .A(n_290), .B(n_309), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_292), .A2(n_302), .B(n_305), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_292), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_293), .B(n_335), .Y(n_334) );
NAND2x1_ASAP7_75t_L g435 ( .A(n_293), .B(n_353), .Y(n_435) );
BUFx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_295), .A2(n_319), .B(n_392), .Y(n_391) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_297), .Y(n_306) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
AND2x2_ASAP7_75t_L g341 ( .A(n_299), .B(n_342), .Y(n_341) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_299), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_299), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND3xp33_ASAP7_75t_SL g397 ( .A(n_305), .B(n_398), .C(n_402), .Y(n_397) );
INVx2_ASAP7_75t_L g422 ( .A(n_305), .Y(n_422) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
OR2x2_ASAP7_75t_L g455 ( .A(n_306), .B(n_456), .Y(n_455) );
BUFx3_ASAP7_75t_L g333 ( .A(n_307), .Y(n_333) );
NAND2x1_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AOI311xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_315), .A3(n_319), .B(n_324), .C(n_336), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_317), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g344 ( .A(n_317), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_318), .B(n_345), .Y(n_379) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g429 ( .A(n_321), .B(n_417), .Y(n_429) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g395 ( .A(n_322), .B(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_322), .Y(n_478) );
BUFx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI222xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_328), .B1(n_330), .B2(n_332), .C1(n_333), .C2(n_334), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OR2x2_ASAP7_75t_L g386 ( .A(n_326), .B(n_375), .Y(n_386) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_331), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g380 ( .A(n_331), .B(n_350), .Y(n_380) );
AND2x2_ASAP7_75t_L g416 ( .A(n_331), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g426 ( .A(n_331), .B(n_365), .Y(n_426) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_338), .A2(n_347), .B(n_351), .Y(n_346) );
AND2x2_ASAP7_75t_L g367 ( .A(n_339), .B(n_365), .Y(n_367) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_352), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g466 ( .A(n_352), .B(n_467), .Y(n_466) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_352), .Y(n_480) );
INVxp67_ASAP7_75t_SL g414 ( .A(n_353), .Y(n_414) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx3_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_354), .Y(n_467) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND3x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_393), .C(n_421), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_385), .Y(n_358) );
OAI211xp5_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_361), .B(n_366), .C(n_373), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_361), .B(n_477), .Y(n_476) );
OR2x6_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g376 ( .A(n_364), .Y(n_376) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI21xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B(n_372), .Y(n_366) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g394 ( .A(n_369), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_371), .Y(n_463) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_377), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g384 ( .A(n_378), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_380), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_389), .B2(n_391), .Y(n_385) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI211xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B(n_407), .C(n_412), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_398), .A2(n_408), .B1(n_409), .B2(n_411), .Y(n_407) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g451 ( .A(n_405), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_SL g425 ( .A(n_406), .Y(n_425) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_406), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_418), .B2(n_420), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_424), .B2(n_426), .C(n_427), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B(n_435), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OR2x6_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .Y(n_430) );
INVxp67_ASAP7_75t_SL g453 ( .A(n_431), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
AND4x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_443), .C(n_459), .D(n_471), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g470 ( .A(n_442), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_446), .B1(n_448), .B2(n_453), .C(n_454), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_464), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_468), .B(n_470), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_476), .B1(n_480), .B2(n_481), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_SL g841 ( .A(n_482), .Y(n_841) );
BUFx8_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND4xp75_ASAP7_75t_L g486 ( .A(n_487), .B(n_700), .C(n_755), .D(n_802), .Y(n_486) );
NOR2x1_ASAP7_75t_L g487 ( .A(n_488), .B(n_650), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_489), .B(n_629), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_553), .B1(n_597), .B2(n_617), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_503), .Y(n_491) );
AND2x2_ASAP7_75t_L g635 ( .A(n_492), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g675 ( .A(n_492), .B(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g689 ( .A(n_492), .B(n_622), .Y(n_689) );
INVx2_ASAP7_75t_L g706 ( .A(n_492), .Y(n_706) );
INVx2_ASAP7_75t_L g766 ( .A(n_492), .Y(n_766) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g620 ( .A(n_493), .B(n_621), .Y(n_620) );
AND2x4_ASAP7_75t_L g628 ( .A(n_493), .B(n_541), .Y(n_628) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g687 ( .A(n_494), .Y(n_687) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_525), .Y(n_503) );
INVx1_ASAP7_75t_L g637 ( .A(n_504), .Y(n_637) );
INVxp67_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g732 ( .A(n_505), .B(n_621), .Y(n_732) );
AND2x2_ASAP7_75t_L g746 ( .A(n_505), .B(n_526), .Y(n_746) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g623 ( .A(n_506), .B(n_526), .Y(n_623) );
AND2x2_ASAP7_75t_L g719 ( .A(n_506), .B(n_526), .Y(n_719) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g644 ( .A(n_507), .Y(n_644) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_516), .B(n_524), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_513), .B(n_515), .Y(n_508) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_521), .B(n_522), .Y(n_516) );
AO21x1_ASAP7_75t_L g603 ( .A1(n_521), .A2(n_604), .B(n_607), .Y(n_603) );
AOI21x1_ASAP7_75t_L g609 ( .A1(n_521), .A2(n_610), .B(n_612), .Y(n_609) );
AND2x2_ASAP7_75t_L g636 ( .A(n_525), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g676 ( .A(n_525), .Y(n_676) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_540), .Y(n_525) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_526), .Y(n_626) );
INVx2_ASAP7_75t_SL g661 ( .A(n_526), .Y(n_661) );
INVx1_ASAP7_75t_L g670 ( .A(n_526), .Y(n_670) );
AND2x2_ASAP7_75t_L g831 ( .A(n_526), .B(n_687), .Y(n_831) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_535), .B(n_539), .Y(n_526) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B1(n_531), .B2(n_532), .Y(n_528) );
INVx1_ASAP7_75t_L g704 ( .A(n_540), .Y(n_704) );
INVx2_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g621 ( .A(n_541), .Y(n_621) );
AND2x2_ASAP7_75t_L g669 ( .A(n_541), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g686 ( .A(n_541), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g759 ( .A(n_541), .Y(n_759) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_580), .Y(n_553) );
OR2x2_ASAP7_75t_L g837 ( .A(n_554), .B(n_798), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_568), .Y(n_554) );
INVx2_ASAP7_75t_L g598 ( .A(n_555), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_555), .B(n_584), .Y(n_667) );
AND2x2_ASAP7_75t_L g691 ( .A(n_555), .B(n_634), .Y(n_691) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g632 ( .A(n_556), .Y(n_632) );
OAI21x1_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_559), .B(n_567), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B(n_563), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_563), .A2(n_571), .B(n_574), .C(n_578), .Y(n_570) );
INVx1_ASAP7_75t_L g583 ( .A(n_568), .Y(n_583) );
INVx1_ASAP7_75t_L g600 ( .A(n_568), .Y(n_600) );
INVx2_ASAP7_75t_L g656 ( .A(n_568), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_568), .B(n_601), .Y(n_665) );
AND2x2_ASAP7_75t_L g697 ( .A(n_568), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g709 ( .A(n_568), .B(n_584), .Y(n_709) );
INVx1_ASAP7_75t_L g787 ( .A(n_568), .Y(n_787) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g639 ( .A(n_582), .Y(n_639) );
AND2x2_ASAP7_75t_L g733 ( .A(n_582), .B(n_647), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_582), .B(n_714), .Y(n_735) );
AND2x4_ASAP7_75t_L g794 ( .A(n_582), .B(n_749), .Y(n_794) );
AND2x4_ASAP7_75t_L g809 ( .A(n_582), .B(n_810), .Y(n_809) );
AND2x4_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g781 ( .A(n_584), .Y(n_781) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx3_ASAP7_75t_L g634 ( .A(n_585), .Y(n_634) );
AOI21x1_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_591), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B(n_595), .Y(n_592) );
AND2x4_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g726 ( .A(n_598), .B(n_664), .Y(n_726) );
INVx1_ASAP7_75t_L g761 ( .A(n_598), .Y(n_761) );
INVx2_ASAP7_75t_L g810 ( .A(n_598), .Y(n_810) );
AND2x2_ASAP7_75t_L g828 ( .A(n_598), .B(n_709), .Y(n_828) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_599), .Y(n_712) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g724 ( .A(n_601), .Y(n_724) );
AND2x2_ASAP7_75t_L g752 ( .A(n_601), .B(n_634), .Y(n_752) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx3_ASAP7_75t_L g649 ( .A(n_602), .Y(n_649) );
INVx1_ASAP7_75t_L g699 ( .A(n_602), .Y(n_699) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_609), .B(n_615), .Y(n_602) );
INVxp67_ASAP7_75t_L g616 ( .A(n_607), .Y(n_616) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_624), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
AND2x4_ASAP7_75t_SL g727 ( .A(n_620), .B(n_660), .Y(n_727) );
AND2x4_ASAP7_75t_L g777 ( .A(n_622), .B(n_628), .Y(n_777) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g763 ( .A(n_623), .B(n_647), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_623), .Y(n_767) );
OAI222xp33_ASAP7_75t_L g832 ( .A1(n_624), .A2(n_833), .B1(n_835), .B2(n_837), .C1(n_838), .C2(n_840), .Y(n_832) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g684 ( .A(n_626), .Y(n_684) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_628), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g658 ( .A(n_628), .Y(n_658) );
AND2x2_ASAP7_75t_L g694 ( .A(n_628), .B(n_684), .Y(n_694) );
AND2x2_ASAP7_75t_L g745 ( .A(n_628), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g783 ( .A(n_628), .B(n_718), .Y(n_783) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_635), .B(n_638), .C(n_645), .Y(n_629) );
AND2x4_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g673 ( .A(n_631), .Y(n_673) );
AND2x4_ASAP7_75t_L g682 ( .A(n_631), .B(n_634), .Y(n_682) );
BUFx2_ASAP7_75t_L g749 ( .A(n_631), .Y(n_749) );
AND2x2_ASAP7_75t_L g774 ( .A(n_631), .B(n_656), .Y(n_774) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x4_ASAP7_75t_L g714 ( .A(n_632), .B(n_649), .Y(n_714) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g655 ( .A(n_634), .B(n_656), .Y(n_655) );
BUFx2_ASAP7_75t_L g773 ( .A(n_634), .Y(n_773) );
INVx2_ASAP7_75t_SL g801 ( .A(n_636), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_642), .B(n_686), .Y(n_812) );
AND2x2_ASAP7_75t_L g821 ( .A(n_642), .B(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g703 ( .A(n_643), .B(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_643), .B(n_704), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_643), .B(n_687), .Y(n_818) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g660 ( .A(n_644), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g826 ( .A(n_644), .B(n_687), .Y(n_826) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g654 ( .A(n_647), .B(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g739 ( .A(n_647), .B(n_725), .Y(n_739) );
AND2x2_ASAP7_75t_L g793 ( .A(n_647), .B(n_794), .Y(n_793) );
AND2x2_ASAP7_75t_L g800 ( .A(n_647), .B(n_682), .Y(n_800) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_677), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_657), .B1(n_662), .B2(n_668), .C(n_671), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x4_ASAP7_75t_L g672 ( .A(n_655), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g814 ( .A(n_655), .Y(n_814) );
INVx1_ASAP7_75t_L g750 ( .A(n_656), .Y(n_750) );
OR2x6_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_659), .A2(n_711), .B1(n_713), .B2(n_715), .Y(n_710) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g705 ( .A(n_660), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g731 ( .A(n_661), .B(n_687), .Y(n_731) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_664), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g680 ( .A(n_665), .Y(n_680) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_L g825 ( .A(n_669), .B(n_826), .Y(n_825) );
AND2x2_ASAP7_75t_L g822 ( .A(n_670), .B(n_759), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_673), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_675), .A2(n_693), .B(n_695), .Y(n_692) );
OR2x2_ASAP7_75t_L g736 ( .A(n_676), .B(n_737), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_692), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_683), .B1(n_688), .B2(n_690), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx2_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g696 ( .A(n_682), .B(n_697), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_682), .A2(n_689), .B1(n_730), .B2(n_733), .C(n_734), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_682), .B(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g768 ( .A(n_686), .B(n_719), .Y(n_768) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_687), .Y(n_717) );
INVx1_ASAP7_75t_L g738 ( .A(n_687), .Y(n_738) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_691), .B(n_712), .Y(n_711) );
BUFx2_ASAP7_75t_L g784 ( .A(n_691), .Y(n_784) );
AND2x2_ASAP7_75t_L g797 ( .A(n_691), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g744 ( .A(n_697), .Y(n_744) );
INVx2_ASAP7_75t_L g798 ( .A(n_698), .Y(n_798) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_699), .Y(n_771) );
NOR2x1_ASAP7_75t_L g700 ( .A(n_701), .B(n_728), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_702), .B(n_720), .Y(n_701) );
O2A1O1Ixp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .B(n_707), .C(n_710), .Y(n_702) );
AND2x2_ASAP7_75t_L g789 ( .A(n_706), .B(n_746), .Y(n_789) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_706), .Y(n_806) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g725 ( .A(n_709), .Y(n_725) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g792 ( .A(n_718), .Y(n_792) );
BUFx3_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_719), .B(n_737), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_726), .B(n_727), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_721), .A2(n_765), .B1(n_768), .B2(n_769), .Y(n_764) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g829 ( .A(n_723), .Y(n_829) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_724), .B(n_781), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_741), .Y(n_728) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_731), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_SL g830 ( .A(n_732), .B(n_831), .Y(n_830) );
AND2x4_ASAP7_75t_L g834 ( .A(n_732), .B(n_737), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_732), .B(n_831), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_739), .B2(n_740), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OA22x2_ASAP7_75t_L g811 ( .A1(n_739), .A2(n_812), .B1(n_813), .B2(n_816), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_745), .B(n_747), .Y(n_741) );
INVxp67_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
AOI21xp33_ASAP7_75t_SL g747 ( .A1(n_748), .A2(n_751), .B(n_753), .Y(n_747) );
NAND2xp33_ASAP7_75t_SL g778 ( .A(n_748), .B(n_779), .Y(n_778) );
OR2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NOR2x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_775), .Y(n_755) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_760), .B(n_764), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g817 ( .A(n_758), .Y(n_817) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2x1_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
OA21x2_ASAP7_75t_L g804 ( .A1(n_763), .A2(n_805), .B(n_807), .Y(n_804) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
AND2x2_ASAP7_75t_L g791 ( .A(n_766), .B(n_792), .Y(n_791) );
INVx2_ASAP7_75t_SL g807 ( .A(n_768), .Y(n_807) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
INVx1_ASAP7_75t_L g782 ( .A(n_770), .Y(n_782) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g823 ( .A(n_772), .Y(n_823) );
AND2x4_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_790), .Y(n_775) );
AOI222xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B1(n_783), .B2(n_784), .C1(n_785), .C2(n_789), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_782), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_786), .A2(n_820), .B1(n_823), .B2(n_824), .C(n_827), .Y(n_819) );
OR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVxp67_ASAP7_75t_SL g836 ( .A(n_788), .Y(n_836) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_793), .B(n_795), .Y(n_790) );
AOI21xp5_ASAP7_75t_SL g795 ( .A1(n_796), .A2(n_799), .B(n_801), .Y(n_795) );
INVx2_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g815 ( .A(n_798), .Y(n_815) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NOR3x1_ASAP7_75t_L g802 ( .A(n_803), .B(n_819), .C(n_832), .Y(n_802) );
OAI21x1_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_808), .B(n_811), .Y(n_803) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
OR2x6_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVx1_ASAP7_75t_L g839 ( .A(n_814), .Y(n_839) );
OR2x2_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
OAI21xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_829), .B(n_830), .Y(n_827) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g846 ( .A(n_843), .Y(n_846) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
OR2x6_ASAP7_75t_L g849 ( .A(n_850), .B(n_852), .Y(n_849) );
OR2x2_ASAP7_75t_L g876 ( .A(n_850), .B(n_877), .Y(n_876) );
INVx2_ASAP7_75t_SL g850 ( .A(n_851), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g855 ( .A(n_851), .Y(n_855) );
INVx2_ASAP7_75t_L g868 ( .A(n_852), .Y(n_868) );
OAI21xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_856), .B(n_873), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g854 ( .A(n_855), .Y(n_854) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_861), .B1(n_869), .B2(n_870), .C(n_871), .Y(n_856) );
INVx1_ASAP7_75t_L g869 ( .A(n_857), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
INVx4_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_865), .B(n_872), .Y(n_871) );
BUFx12f_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
BUFx6f_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx5_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
BUFx12f_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
endmodule