module fake_netlist_5_464_n_1758 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1758);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1758;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_44),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_12),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_113),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_115),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_21),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_17),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_83),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_74),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_39),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_36),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_109),
.Y(n_177)
);

BUFx2_ASAP7_75t_SL g178 ( 
.A(n_85),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_94),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_75),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_140),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_95),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_91),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_25),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_50),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_55),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_126),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_122),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_116),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_78),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_39),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_35),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_43),
.Y(n_194)
);

BUFx2_ASAP7_75t_SL g195 ( 
.A(n_61),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_104),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_49),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_52),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_6),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_105),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_41),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_30),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_63),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_53),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_31),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_154),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_59),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_135),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_45),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_34),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_134),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_31),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_60),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_121),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_57),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_143),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_16),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_45),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_110),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_6),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_34),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_89),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_14),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_90),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_27),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_97),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_124),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_118),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_106),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_88),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_4),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_17),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_19),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_103),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_107),
.Y(n_238)
);

BUFx2_ASAP7_75t_SL g239 ( 
.A(n_80),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_10),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_36),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_84),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_19),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_13),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_21),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_26),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_15),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_150),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_133),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_28),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_1),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_117),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_13),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_18),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_30),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_93),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_5),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_51),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_62),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_54),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_123),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_66),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_20),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_138),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_142),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_3),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_37),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_7),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_67),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_1),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_10),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_25),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_44),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_77),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_100),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_111),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_11),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_38),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_146),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_56),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_43),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_70),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_76),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_40),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_64),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_29),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_38),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_79),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_2),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_16),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_11),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_108),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_96),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_72),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_3),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_48),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_35),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_12),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_46),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_87),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_15),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_155),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_65),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_14),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_68),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_92),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_24),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_4),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_32),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_192),
.B(n_0),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_212),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_254),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_234),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_185),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_234),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_268),
.B(n_2),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_5),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_199),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_193),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_161),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_193),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_201),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_198),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_193),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_208),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_169),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_193),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_193),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_207),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_202),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_220),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_220),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_222),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_248),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_275),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_301),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_164),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_206),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_220),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_221),
.Y(n_344)
);

INVxp33_ASAP7_75t_SL g345 ( 
.A(n_156),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_224),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_210),
.B(n_7),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_220),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_226),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_236),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_156),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_220),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_162),
.B(n_8),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_282),
.B(n_8),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_240),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_235),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_243),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_235),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_244),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_183),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_184),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_235),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_235),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_187),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_264),
.B(n_9),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_235),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_164),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_267),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_209),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_264),
.B(n_9),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_245),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_247),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_267),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_267),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_189),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_267),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_162),
.B(n_18),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_250),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_158),
.Y(n_381)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_331),
.A2(n_310),
.B(n_271),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_331),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_332),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_371),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_371),
.Y(n_386)
);

NAND2x1p5_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_230),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_371),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_371),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_322),
.B(n_186),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_325),
.B(n_267),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_328),
.B(n_230),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_335),
.B(n_157),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_336),
.B(n_157),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_371),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_313),
.B(n_186),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_312),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_378),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_378),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_343),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_352),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_356),
.B(n_359),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_364),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_280),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_368),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_370),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_375),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_315),
.B(n_280),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_317),
.A2(n_271),
.B(n_310),
.Y(n_413)
);

AND3x1_ASAP7_75t_L g414 ( 
.A(n_353),
.B(n_213),
.C(n_194),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_320),
.B(n_167),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_323),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_311),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_381),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_362),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_367),
.B(n_167),
.Y(n_420)
);

AND2x2_ASAP7_75t_SL g421 ( 
.A(n_379),
.B(n_173),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_363),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_311),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_312),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_372),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_327),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_319),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_329),
.Y(n_429)
);

BUFx8_ASAP7_75t_L g430 ( 
.A(n_360),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_314),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_354),
.A2(n_223),
.B(n_215),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_318),
.B(n_163),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_316),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_345),
.B(n_214),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_316),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_L g437 ( 
.A(n_314),
.B(n_209),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_321),
.Y(n_438)
);

AND3x2_ASAP7_75t_L g439 ( 
.A(n_358),
.B(n_216),
.C(n_173),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_321),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_351),
.A2(n_166),
.B1(n_305),
.B2(n_174),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_326),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_326),
.B(n_163),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_334),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_334),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_386),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_386),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_386),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_342),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_404),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

NOR3xp33_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_369),
.C(n_341),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_426),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_391),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_391),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_366),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_391),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_391),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_391),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_421),
.B(n_342),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_421),
.B(n_344),
.Y(n_467)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_386),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_410),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_392),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_410),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_392),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_407),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_410),
.Y(n_474)
);

NOR2x1p5_ASAP7_75t_L g475 ( 
.A(n_424),
.B(n_431),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_421),
.B(n_344),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_432),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_377),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_410),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_390),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_386),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_427),
.B(n_346),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_426),
.B(n_427),
.Y(n_483)
);

OAI22xp33_ASAP7_75t_SL g484 ( 
.A1(n_387),
.A2(n_380),
.B1(n_374),
.B2(n_373),
.Y(n_484)
);

OR2x6_ASAP7_75t_L g485 ( 
.A(n_426),
.B(n_427),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_407),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_427),
.B(n_346),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_417),
.B(n_216),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_429),
.B(n_349),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_417),
.B(n_349),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_417),
.B(n_350),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_429),
.B(n_350),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_387),
.B(n_306),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_417),
.B(n_355),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_432),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_394),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_417),
.B(n_159),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_419),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_390),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_386),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_426),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_400),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_426),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_423),
.A2(n_228),
.B1(n_241),
.B2(n_246),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_407),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_429),
.B(n_355),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_386),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_387),
.B(n_445),
.Y(n_511)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_435),
.B(n_361),
.C(n_357),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_423),
.B(n_306),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_423),
.B(n_357),
.Y(n_515)
);

AND2x6_ASAP7_75t_L g516 ( 
.A(n_423),
.B(n_209),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_419),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_387),
.B(n_209),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_429),
.B(n_361),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_432),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_400),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_440),
.B(n_373),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_388),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_401),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_407),
.Y(n_525)
);

BUFx10_ASAP7_75t_L g526 ( 
.A(n_445),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_401),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_402),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_445),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_423),
.B(n_374),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_398),
.B(n_324),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_388),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_402),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_415),
.B(n_397),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_387),
.B(n_209),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_401),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_413),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_418),
.B(n_269),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_413),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_399),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_426),
.Y(n_541)
);

INVx8_ASAP7_75t_L g542 ( 
.A(n_445),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_413),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_403),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_413),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_403),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_415),
.B(n_160),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_383),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_418),
.B(n_285),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_420),
.A2(n_432),
.B1(n_413),
.B2(n_382),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_433),
.B(n_170),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_445),
.B(n_307),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_433),
.B(n_190),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_388),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_388),
.Y(n_555)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_394),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_399),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_399),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_440),
.B(n_340),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_432),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_383),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_388),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_388),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_399),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_409),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_422),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_442),
.B(n_330),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_420),
.A2(n_195),
.B1(n_178),
.B2(n_239),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_428),
.B(n_191),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_413),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_426),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_388),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_388),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_445),
.B(n_307),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_406),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_426),
.B(n_176),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_384),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_389),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_422),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_445),
.B(n_307),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_389),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_430),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_409),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_389),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_445),
.B(n_307),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_428),
.B(n_307),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_389),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_389),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_384),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_430),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_405),
.Y(n_592)
);

OAI21xp33_ASAP7_75t_SL g593 ( 
.A1(n_428),
.A2(n_218),
.B(n_188),
.Y(n_593)
);

AO22x2_ASAP7_75t_L g594 ( 
.A1(n_414),
.A2(n_219),
.B1(n_297),
.B2(n_294),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_482),
.B(n_436),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_450),
.B(n_465),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_495),
.A2(n_499),
.B1(n_535),
.B2(n_518),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_467),
.B(n_446),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_476),
.B(n_446),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_498),
.B(n_434),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_556),
.B(n_434),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_522),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_487),
.B(n_434),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_491),
.B(n_436),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_494),
.B(n_434),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_534),
.B(n_456),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_508),
.B(n_436),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_511),
.B(n_526),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_542),
.B(n_442),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_480),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_519),
.B(n_434),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_457),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_592),
.B(n_444),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_511),
.B(n_526),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_480),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_489),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_526),
.B(n_444),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_470),
.B(n_444),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_492),
.A2(n_446),
.B1(n_444),
.B2(n_414),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_489),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_501),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_529),
.B(n_446),
.Y(n_622)
);

AND2x6_ASAP7_75t_L g623 ( 
.A(n_537),
.B(n_444),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_501),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_517),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_493),
.B(n_446),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_515),
.A2(n_424),
.B1(n_431),
.B2(n_338),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_529),
.B(n_484),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_461),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_462),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_496),
.B(n_438),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_472),
.B(n_551),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_504),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_492),
.B(n_395),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_534),
.B(n_499),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_529),
.B(n_438),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_463),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_534),
.B(n_395),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_504),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_509),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_499),
.B(n_420),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_458),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_530),
.B(n_420),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_553),
.B(n_420),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_473),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_568),
.B(n_420),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_456),
.B(n_438),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_503),
.B(n_424),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_460),
.A2(n_437),
.B1(n_333),
.B2(n_337),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_478),
.A2(n_437),
.B1(n_339),
.B2(n_431),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_537),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_509),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_542),
.B(n_197),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_458),
.Y(n_654)
);

INVx5_ASAP7_75t_L g655 ( 
.A(n_488),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_515),
.B(n_424),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_538),
.B(n_398),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_521),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_512),
.B(n_398),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_548),
.B(n_415),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_561),
.B(n_397),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_578),
.B(n_397),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_531),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_503),
.B(n_431),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_464),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_486),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_521),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_590),
.B(n_411),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_475),
.B(n_425),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_490),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_L g671 ( 
.A(n_542),
.B(n_200),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_507),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_569),
.B(n_430),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_505),
.B(n_430),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_538),
.Y(n_675)
);

OAI221xp5_ASAP7_75t_L g676 ( 
.A1(n_506),
.A2(n_441),
.B1(n_425),
.B2(n_416),
.C(n_393),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_539),
.A2(n_441),
.B(n_425),
.C(n_411),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_464),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_505),
.B(n_430),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_513),
.B(n_411),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_525),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_541),
.B(n_439),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_539),
.B(n_416),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_543),
.B(n_416),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_541),
.B(n_439),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_517),
.Y(n_686)
);

INVxp33_ASAP7_75t_L g687 ( 
.A(n_549),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_549),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_524),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_572),
.B(n_204),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_543),
.B(n_416),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_572),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_495),
.A2(n_382),
.B1(n_270),
.B2(n_231),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_545),
.B(n_382),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_545),
.B(n_382),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_483),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_528),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_524),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_571),
.B(n_382),
.Y(n_699)
);

NOR3xp33_ASAP7_75t_L g700 ( 
.A(n_559),
.B(n_253),
.C(n_257),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_567),
.B(n_393),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_527),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_483),
.B(n_168),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_527),
.Y(n_704)
);

AND2x6_ASAP7_75t_SL g705 ( 
.A(n_577),
.B(n_205),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_571),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_550),
.B(n_238),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_500),
.B(n_158),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_536),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_477),
.B(n_252),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_533),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_566),
.Y(n_712)
);

NOR3xp33_ASAP7_75t_L g713 ( 
.A(n_454),
.B(n_272),
.C(n_273),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_483),
.B(n_251),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_544),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_483),
.A2(n_217),
.B1(n_196),
.B2(n_203),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_547),
.B(n_546),
.C(n_485),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_547),
.B(n_382),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_565),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_536),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_485),
.B(n_255),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_485),
.B(n_258),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_565),
.Y(n_723)
);

AND2x2_ASAP7_75t_SL g724 ( 
.A(n_466),
.B(n_256),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_584),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_485),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_477),
.B(n_261),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_547),
.B(n_409),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_584),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_477),
.B(n_262),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_451),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_580),
.B(n_165),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_518),
.B(n_412),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_577),
.B(n_276),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_451),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_535),
.B(n_412),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_488),
.B(n_412),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_447),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_488),
.B(n_408),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_452),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_566),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_452),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_488),
.B(n_408),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_583),
.B(n_274),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_594),
.B(n_278),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_488),
.B(n_408),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_453),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_447),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_453),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_497),
.B(n_281),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_455),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_577),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_497),
.B(n_283),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_455),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_488),
.B(n_408),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_469),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_514),
.B(n_408),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_447),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_497),
.B(n_211),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_520),
.B(n_168),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_SL g761 ( 
.A(n_520),
.B(n_165),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_514),
.B(n_520),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_560),
.B(n_225),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_577),
.B(n_405),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_469),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_560),
.B(n_570),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_641),
.A2(n_542),
.B(n_570),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_766),
.A2(n_560),
.B(n_570),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_611),
.B(n_594),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_645),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_602),
.B(n_591),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_608),
.A2(n_552),
.B(n_575),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_608),
.A2(n_614),
.B(n_694),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_723),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_595),
.A2(n_593),
.B(n_575),
.C(n_552),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_634),
.B(n_594),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_604),
.B(n_591),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_596),
.B(n_594),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_675),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_607),
.B(n_581),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_614),
.A2(n_581),
.B(n_586),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_596),
.B(n_514),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_657),
.B(n_586),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_632),
.B(n_514),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_623),
.B(n_514),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_695),
.A2(n_523),
.B(n_502),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_699),
.A2(n_671),
.B(n_653),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_SL g788 ( 
.A1(n_712),
.A2(n_290),
.B1(n_171),
.B2(n_287),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_603),
.B(n_605),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_654),
.B(n_514),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_613),
.B(n_516),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_726),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_677),
.A2(n_471),
.B(n_474),
.C(n_479),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_666),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_723),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_683),
.A2(n_589),
.B(n_588),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_670),
.Y(n_797)
);

OAI321xp33_ASAP7_75t_L g798 ( 
.A1(n_619),
.A2(n_299),
.A3(n_287),
.B1(n_288),
.B2(n_290),
.C(n_291),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_626),
.B(n_516),
.Y(n_799)
);

O2A1O1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_677),
.A2(n_471),
.B(n_474),
.C(n_479),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_638),
.B(n_516),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_701),
.B(n_516),
.Y(n_802)
);

NOR2x1_ASAP7_75t_L g803 ( 
.A(n_636),
.B(n_656),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_600),
.B(n_601),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_684),
.A2(n_691),
.B(n_718),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_631),
.A2(n_589),
.B(n_588),
.C(n_585),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_610),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_708),
.Y(n_808)
);

CKINVDCx10_ASAP7_75t_R g809 ( 
.A(n_712),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_618),
.B(n_516),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_653),
.A2(n_448),
.B(n_502),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_651),
.B(n_516),
.Y(n_812)
);

O2A1O1Ixp5_ASAP7_75t_L g813 ( 
.A1(n_598),
.A2(n_589),
.B(n_588),
.C(n_459),
.Y(n_813)
);

NOR2xp67_ASAP7_75t_L g814 ( 
.A(n_650),
.B(n_227),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_671),
.A2(n_448),
.B(n_523),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_643),
.B(n_459),
.Y(n_816)
);

INVxp67_ASAP7_75t_SL g817 ( 
.A(n_706),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_644),
.A2(n_448),
.B(n_523),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_654),
.B(n_459),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_762),
.A2(n_502),
.B(n_523),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_597),
.A2(n_182),
.B1(n_304),
.B2(n_295),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_732),
.Y(n_822)
);

O2A1O1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_647),
.A2(n_557),
.B(n_540),
.C(n_558),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_706),
.B(n_481),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_635),
.A2(n_502),
.B(n_449),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_606),
.B(n_724),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_710),
.A2(n_555),
.B(n_585),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_707),
.A2(n_622),
.B(n_617),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_647),
.A2(n_557),
.B(n_540),
.C(n_558),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_687),
.B(n_171),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_606),
.A2(n_587),
.B1(n_585),
.B2(n_582),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_707),
.A2(n_449),
.B(n_448),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_617),
.A2(n_449),
.B(n_576),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_706),
.B(n_481),
.Y(n_834)
);

NOR3xp33_ASAP7_75t_L g835 ( 
.A(n_627),
.B(n_289),
.C(n_182),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_606),
.B(n_481),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_687),
.B(n_172),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_598),
.A2(n_564),
.B(n_582),
.C(n_579),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_672),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_659),
.B(n_172),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_681),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_680),
.B(n_510),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_726),
.A2(n_295),
.B1(n_304),
.B2(n_293),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_661),
.B(n_510),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_622),
.A2(n_609),
.B(n_710),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_760),
.A2(n_510),
.B(n_582),
.C(n_579),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_662),
.B(n_532),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_668),
.B(n_697),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_688),
.B(n_175),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_612),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_703),
.A2(n_599),
.B(n_673),
.C(n_717),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_609),
.A2(n_449),
.B(n_576),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_727),
.A2(n_576),
.B(n_562),
.Y(n_853)
);

INVx5_ASAP7_75t_L g854 ( 
.A(n_623),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_727),
.A2(n_579),
.B(n_573),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_610),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_642),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_663),
.B(n_174),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_665),
.Y(n_859)
);

AO21x1_ASAP7_75t_L g860 ( 
.A1(n_599),
.A2(n_564),
.B(n_396),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_642),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_761),
.A2(n_587),
.B1(n_555),
.B2(n_573),
.Y(n_862)
);

AOI21x1_ASAP7_75t_L g863 ( 
.A1(n_730),
.A2(n_385),
.B(n_396),
.Y(n_863)
);

BUFx12f_ASAP7_75t_L g864 ( 
.A(n_625),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_730),
.A2(n_562),
.B(n_574),
.Y(n_865)
);

NOR2x1_ASAP7_75t_L g866 ( 
.A(n_636),
.B(n_532),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_649),
.B(n_175),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_711),
.B(n_532),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_724),
.B(n_177),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_750),
.A2(n_562),
.B(n_574),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_615),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_623),
.B(n_555),
.Y(n_872)
);

INVx5_ASAP7_75t_L g873 ( 
.A(n_623),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_642),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_750),
.A2(n_574),
.B(n_563),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_623),
.B(n_573),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_753),
.A2(n_574),
.B(n_563),
.Y(n_877)
);

CKINVDCx16_ASAP7_75t_R g878 ( 
.A(n_745),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_744),
.B(n_288),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_753),
.A2(n_587),
.B(n_396),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_655),
.A2(n_574),
.B(n_563),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_615),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_655),
.A2(n_563),
.B(n_562),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_655),
.A2(n_563),
.B(n_562),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_655),
.A2(n_447),
.B(n_554),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_623),
.B(n_447),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_655),
.A2(n_692),
.B(n_759),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_665),
.B(n_177),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_678),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_686),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_669),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_616),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_676),
.A2(n_696),
.B(n_628),
.C(n_660),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_629),
.B(n_587),
.Y(n_894)
);

INVx6_ASAP7_75t_L g895 ( 
.A(n_705),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_646),
.A2(n_179),
.B1(n_181),
.B2(n_289),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_692),
.A2(n_554),
.B(n_468),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_759),
.A2(n_554),
.B(n_468),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_616),
.Y(n_899)
);

NAND2xp33_ASAP7_75t_L g900 ( 
.A(n_758),
.B(n_587),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_741),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_763),
.A2(n_554),
.B(n_468),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_715),
.B(n_179),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_630),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_763),
.A2(n_587),
.B(n_385),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_714),
.B(n_181),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_721),
.B(n_293),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_758),
.A2(n_554),
.B(n_468),
.Y(n_908)
);

NOR2x1_ASAP7_75t_L g909 ( 
.A(n_628),
.B(n_385),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_SL g910 ( 
.A1(n_739),
.A2(n_385),
.B(n_396),
.C(n_164),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_637),
.B(n_468),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_620),
.B(n_621),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_620),
.B(n_406),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_621),
.B(n_406),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_624),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_758),
.A2(n_389),
.B(n_406),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_624),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_633),
.Y(n_918)
);

AOI21x1_ASAP7_75t_L g919 ( 
.A1(n_743),
.A2(n_389),
.B(n_406),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_758),
.A2(n_389),
.B(n_406),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_648),
.A2(n_233),
.B(n_232),
.C(n_229),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_722),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_693),
.A2(n_284),
.B1(n_259),
.B2(n_237),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_728),
.A2(n_406),
.B(n_242),
.Y(n_924)
);

BUFx4f_ASAP7_75t_L g925 ( 
.A(n_734),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_737),
.A2(n_406),
.B(n_286),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_639),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_746),
.A2(n_249),
.B(n_260),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_734),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_761),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_639),
.B(n_640),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_678),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_755),
.A2(n_263),
.B(n_265),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_678),
.B(n_266),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_640),
.B(n_277),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_652),
.B(n_309),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_752),
.A2(n_679),
.B1(n_674),
.B2(n_664),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_757),
.A2(n_279),
.B(n_300),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_L g939 ( 
.A1(n_700),
.A2(n_309),
.B(n_296),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_652),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_658),
.B(n_291),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_658),
.B(n_292),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_682),
.A2(n_300),
.B(n_299),
.Y(n_943)
);

OAI321xp33_ASAP7_75t_L g944 ( 
.A1(n_685),
.A2(n_296),
.A3(n_292),
.B1(n_303),
.B2(n_180),
.C(n_26),
.Y(n_944)
);

O2A1O1Ixp5_ASAP7_75t_L g945 ( 
.A1(n_690),
.A2(n_303),
.B(n_180),
.C(n_73),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_667),
.B(n_71),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_764),
.B(n_303),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_648),
.A2(n_69),
.B(n_152),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_738),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_764),
.B(n_716),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_667),
.B(n_702),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_738),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_713),
.B(n_58),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_664),
.A2(n_736),
.B(n_733),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_792),
.B(n_674),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_774),
.Y(n_956)
);

BUFx2_ASAP7_75t_R g957 ( 
.A(n_890),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_770),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_780),
.A2(n_679),
.B1(n_764),
.B2(n_738),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_808),
.B(n_734),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_776),
.A2(n_690),
.B1(n_725),
.B2(n_729),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_840),
.A2(n_719),
.B(n_689),
.C(n_698),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_792),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_779),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_822),
.B(n_689),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_854),
.A2(n_748),
.B(n_702),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_859),
.B(n_698),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_L g968 ( 
.A(n_867),
.B(n_748),
.C(n_704),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_893),
.A2(n_704),
.B(n_709),
.C(n_720),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_854),
.A2(n_748),
.B(n_709),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_859),
.B(n_720),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_854),
.A2(n_765),
.B(n_756),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_863),
.A2(n_765),
.B(n_756),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_848),
.B(n_754),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_805),
.A2(n_754),
.B(n_751),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_944),
.A2(n_735),
.B(n_749),
.C(n_742),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_792),
.B(n_751),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_891),
.B(n_747),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_830),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_932),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_789),
.B(n_747),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_771),
.B(n_777),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_804),
.B(n_740),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_854),
.A2(n_740),
.B1(n_731),
.B2(n_180),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_873),
.A2(n_731),
.B(n_81),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_776),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_922),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_907),
.B(n_22),
.Y(n_988)
);

AO22x1_ASAP7_75t_L g989 ( 
.A1(n_835),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_989)
);

OR2x4_ASAP7_75t_L g990 ( 
.A(n_858),
.B(n_28),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_851),
.A2(n_29),
.B(n_32),
.C(n_33),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_773),
.A2(n_33),
.B(n_37),
.C(n_40),
.Y(n_992)
);

BUFx12f_ASAP7_75t_L g993 ( 
.A(n_864),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_SL g994 ( 
.A(n_878),
.B(n_41),
.C(n_42),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_879),
.B(n_42),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_873),
.A2(n_102),
.B1(n_141),
.B2(n_82),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_859),
.B(n_112),
.Y(n_997)
);

OR2x6_ASAP7_75t_L g998 ( 
.A(n_901),
.B(n_101),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_794),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_925),
.B(n_132),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_784),
.A2(n_46),
.B(n_47),
.C(n_86),
.Y(n_1001)
);

OAI21xp33_ASAP7_75t_SL g1002 ( 
.A1(n_826),
.A2(n_47),
.B(n_98),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_783),
.B(n_936),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_828),
.A2(n_99),
.B(n_136),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_795),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_797),
.B(n_137),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_807),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_873),
.A2(n_139),
.B1(n_148),
.B2(n_769),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_925),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_869),
.A2(n_769),
.B(n_798),
.C(n_778),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_788),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_839),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_888),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_841),
.B(n_850),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_932),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_904),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_778),
.A2(n_950),
.B1(n_803),
.B2(n_953),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_895),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_837),
.B(n_849),
.Y(n_1019)
);

CKINVDCx14_ASAP7_75t_R g1020 ( 
.A(n_895),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_784),
.A2(n_775),
.B(n_772),
.C(n_781),
.Y(n_1021)
);

BUFx10_ASAP7_75t_L g1022 ( 
.A(n_888),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_873),
.A2(n_785),
.B(n_845),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_816),
.A2(n_787),
.B(n_767),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_790),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_906),
.B(n_930),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_936),
.B(n_941),
.Y(n_1027)
);

NOR2xp67_ASAP7_75t_L g1028 ( 
.A(n_929),
.B(n_802),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_953),
.A2(n_896),
.B1(n_947),
.B2(n_790),
.Y(n_1029)
);

NAND2x1p5_ASAP7_75t_L g1030 ( 
.A(n_857),
.B(n_861),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_937),
.A2(n_782),
.B1(n_801),
.B2(n_844),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_817),
.A2(n_861),
.B1(n_857),
.B2(n_889),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_886),
.A2(n_818),
.B(n_887),
.Y(n_1033)
);

CKINVDCx16_ASAP7_75t_R g1034 ( 
.A(n_809),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_886),
.A2(n_786),
.B(n_768),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_941),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_895),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_927),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_856),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_874),
.B(n_889),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_820),
.A2(n_954),
.B(n_824),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_942),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_819),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_943),
.B(n_903),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_834),
.A2(n_796),
.B(n_876),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_942),
.Y(n_1046)
);

INVx8_ASAP7_75t_L g1047 ( 
.A(n_819),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_843),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_847),
.B(n_874),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_871),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_882),
.Y(n_1051)
);

NOR2x1_ASAP7_75t_L g1052 ( 
.A(n_814),
.B(n_934),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_892),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_909),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_939),
.B(n_821),
.C(n_938),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_872),
.A2(n_876),
.B(n_852),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_935),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_912),
.B(n_931),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_935),
.A2(n_806),
.B(n_782),
.C(n_846),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_899),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_949),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_872),
.A2(n_842),
.B(n_853),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_949),
.B(n_952),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_825),
.A2(n_833),
.B(n_812),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_SL g1065 ( 
.A1(n_921),
.A2(n_905),
.B(n_799),
.C(n_793),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_836),
.A2(n_831),
.B1(n_810),
.B2(n_791),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_915),
.B(n_918),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_865),
.A2(n_877),
.B(n_870),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_917),
.Y(n_1069)
);

NAND2xp33_ASAP7_75t_SL g1070 ( 
.A(n_952),
.B(n_946),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_940),
.B(n_868),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_946),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_912),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_931),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_923),
.B(n_951),
.Y(n_1075)
);

BUFx12f_ASAP7_75t_L g1076 ( 
.A(n_945),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_951),
.B(n_866),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_919),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_911),
.Y(n_1079)
);

OA21x2_ASAP7_75t_L g1080 ( 
.A1(n_813),
.A2(n_860),
.B(n_855),
.Y(n_1080)
);

INVx2_ASAP7_75t_SL g1081 ( 
.A(n_913),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_894),
.A2(n_911),
.B1(n_948),
.B2(n_914),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_875),
.A2(n_832),
.B(n_881),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_894),
.B(n_914),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_800),
.A2(n_838),
.B(n_823),
.C(n_829),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_928),
.B(n_933),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_883),
.A2(n_884),
.B(n_827),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_913),
.B(n_880),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_900),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_910),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_898),
.A2(n_902),
.B(n_815),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_811),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_862),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_924),
.A2(n_897),
.B1(n_926),
.B2(n_885),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_916),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_920),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_908),
.A2(n_840),
.B(n_604),
.C(n_607),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_808),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_779),
.Y(n_1099)
);

NOR2xp67_ASAP7_75t_L g1100 ( 
.A(n_891),
.B(n_717),
.Y(n_1100)
);

OAI22x1_ASAP7_75t_L g1101 ( 
.A1(n_988),
.A2(n_1019),
.B1(n_982),
.B2(n_1044),
.Y(n_1101)
);

AO21x2_ASAP7_75t_L g1102 ( 
.A1(n_1024),
.A2(n_1021),
.B(n_1035),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1023),
.A2(n_973),
.B(n_1056),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1027),
.B(n_1074),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_991),
.A2(n_992),
.B(n_1097),
.C(n_1036),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1091),
.A2(n_1033),
.B(n_1064),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1057),
.B(n_1003),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1057),
.B(n_960),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1041),
.A2(n_1058),
.B(n_1087),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1083),
.A2(n_1068),
.B(n_1062),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_975),
.A2(n_1045),
.B(n_1094),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_975),
.A2(n_1059),
.B(n_1078),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1070),
.A2(n_983),
.B(n_981),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1031),
.A2(n_1075),
.B(n_1085),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_SL g1115 ( 
.A(n_957),
.B(n_1093),
.Y(n_1115)
);

INVx8_ASAP7_75t_L g1116 ( 
.A(n_1047),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1073),
.B(n_1046),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1042),
.B(n_979),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1098),
.B(n_1026),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_1009),
.B(n_955),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1065),
.A2(n_1086),
.B(n_959),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1055),
.A2(n_1017),
.B(n_1010),
.C(n_1100),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_995),
.B(n_1098),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_SL g1124 ( 
.A1(n_1001),
.A2(n_1000),
.B(n_1006),
.C(n_997),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1029),
.A2(n_1017),
.B1(n_1100),
.B2(n_1013),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_978),
.B(n_974),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1014),
.B(n_999),
.Y(n_1127)
);

BUFx4f_ASAP7_75t_L g1128 ( 
.A(n_993),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1048),
.A2(n_1002),
.B(n_986),
.C(n_987),
.Y(n_1129)
);

AOI21xp33_ASAP7_75t_L g1130 ( 
.A1(n_1002),
.A2(n_1031),
.B(n_1066),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1012),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1016),
.Y(n_1132)
);

NOR2xp67_ASAP7_75t_L g1133 ( 
.A(n_964),
.B(n_1099),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1072),
.A2(n_962),
.B(n_1077),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_965),
.B(n_994),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1008),
.A2(n_1090),
.B(n_984),
.C(n_998),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_SL g1137 ( 
.A1(n_969),
.A2(n_1054),
.B(n_971),
.C(n_967),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1067),
.Y(n_1138)
);

OA21x2_ASAP7_75t_L g1139 ( 
.A1(n_1082),
.A2(n_961),
.B(n_1096),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1032),
.A2(n_1095),
.A3(n_1093),
.B(n_972),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1049),
.A2(n_1092),
.B(n_970),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1078),
.A2(n_966),
.B(n_1004),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1052),
.A2(n_1028),
.B(n_976),
.C(n_968),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_956),
.Y(n_1144)
);

OAI22x1_ASAP7_75t_L g1145 ( 
.A1(n_955),
.A2(n_961),
.B1(n_1037),
.B2(n_1038),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1082),
.A2(n_985),
.B(n_1040),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1084),
.B(n_1081),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1092),
.A2(n_1015),
.B(n_980),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1009),
.B(n_963),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1088),
.A2(n_1028),
.B(n_1080),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1030),
.A2(n_1040),
.B(n_980),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1030),
.A2(n_1015),
.B(n_1080),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1009),
.B(n_1025),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1043),
.B(n_1079),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1005),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1034),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1071),
.A2(n_1053),
.B(n_1060),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1079),
.B(n_1007),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1043),
.B(n_1079),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1039),
.A2(n_1050),
.B(n_1051),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1092),
.A2(n_1063),
.B(n_977),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1069),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1063),
.A2(n_977),
.B(n_1089),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1047),
.A2(n_996),
.B(n_1069),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1061),
.A2(n_1076),
.A3(n_989),
.B(n_1069),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1025),
.B(n_1047),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_998),
.A2(n_990),
.B1(n_1011),
.B2(n_1020),
.Y(n_1167)
);

AO21x1_ASAP7_75t_L g1168 ( 
.A1(n_998),
.A2(n_1022),
.B(n_1018),
.Y(n_1168)
);

BUFx12f_ASAP7_75t_L g1169 ( 
.A(n_1022),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1023),
.A2(n_542),
.B(n_854),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1034),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1023),
.A2(n_542),
.B(n_854),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1023),
.A2(n_973),
.B(n_1056),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1027),
.B(n_1074),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_958),
.Y(n_1175)
);

AOI221xp5_ASAP7_75t_SL g1176 ( 
.A1(n_988),
.A2(n_991),
.B1(n_1010),
.B2(n_776),
.C(n_677),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1021),
.A2(n_1085),
.A3(n_1090),
.B(n_851),
.Y(n_1177)
);

OA21x2_ASAP7_75t_L g1178 ( 
.A1(n_1021),
.A2(n_1085),
.B(n_1024),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1098),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1027),
.B(n_1074),
.Y(n_1180)
);

AOI221x1_ASAP7_75t_L g1181 ( 
.A1(n_988),
.A2(n_991),
.B1(n_1019),
.B2(n_1055),
.C(n_835),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_963),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_958),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1021),
.A2(n_1031),
.B(n_1059),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_964),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1023),
.A2(n_973),
.B(n_1056),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1018),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_988),
.A2(n_1019),
.B1(n_840),
.B2(n_1044),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_958),
.Y(n_1189)
);

INVx3_ASAP7_75t_SL g1190 ( 
.A(n_1034),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_958),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_963),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1034),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1023),
.A2(n_542),
.B(n_854),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1098),
.B(n_1003),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_L g1196 ( 
.A(n_1019),
.B(n_840),
.C(n_988),
.Y(n_1196)
);

AO32x2_ASAP7_75t_L g1197 ( 
.A1(n_959),
.A2(n_937),
.A3(n_1008),
.B1(n_1066),
.B2(n_1093),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1023),
.A2(n_973),
.B(n_1056),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1023),
.A2(n_542),
.B(n_854),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_958),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1027),
.B(n_1074),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1023),
.A2(n_973),
.B(n_1056),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1019),
.A2(n_1044),
.B(n_988),
.C(n_780),
.Y(n_1203)
);

CKINVDCx6p67_ASAP7_75t_R g1204 ( 
.A(n_1034),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_993),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1021),
.A2(n_1085),
.A3(n_1090),
.B(n_851),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1021),
.A2(n_1031),
.B(n_1059),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_SL g1208 ( 
.A(n_1009),
.B(n_591),
.Y(n_1208)
);

CKINVDCx11_ASAP7_75t_R g1209 ( 
.A(n_1034),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1035),
.A2(n_1091),
.B(n_1033),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1023),
.A2(n_542),
.B(n_854),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1098),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_SL g1213 ( 
.A1(n_1010),
.A2(n_893),
.B(n_778),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1018),
.Y(n_1214)
);

AO32x2_ASAP7_75t_L g1215 ( 
.A1(n_959),
.A2(n_937),
.A3(n_1008),
.B1(n_1066),
.B2(n_1093),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1023),
.A2(n_973),
.B(n_1056),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1019),
.A2(n_1044),
.B(n_988),
.C(n_780),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1027),
.B(n_1074),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1023),
.A2(n_973),
.B(n_1056),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1098),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1023),
.A2(n_542),
.B(n_854),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1023),
.A2(n_542),
.B(n_854),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1023),
.A2(n_542),
.B(n_854),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1063),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1023),
.A2(n_542),
.B(n_854),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_988),
.A2(n_1019),
.B1(n_840),
.B2(n_1044),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1023),
.A2(n_542),
.B(n_854),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1023),
.A2(n_973),
.B(n_1056),
.Y(n_1228)
);

O2A1O1Ixp5_ASAP7_75t_SL g1229 ( 
.A1(n_1090),
.A2(n_628),
.B(n_495),
.C(n_599),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1042),
.B(n_701),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1021),
.A2(n_1031),
.B(n_1059),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1021),
.A2(n_1031),
.B(n_1059),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1063),
.Y(n_1233)
);

AO22x2_ASAP7_75t_L g1234 ( 
.A1(n_1008),
.A2(n_835),
.B1(n_937),
.B2(n_959),
.Y(n_1234)
);

AOI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1035),
.A2(n_1091),
.B(n_1033),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1196),
.A2(n_1226),
.B1(n_1188),
.B2(n_1101),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1131),
.Y(n_1237)
);

INVx5_ASAP7_75t_L g1238 ( 
.A(n_1192),
.Y(n_1238)
);

INVx3_ASAP7_75t_SL g1239 ( 
.A(n_1204),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1230),
.B(n_1123),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1183),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1196),
.A2(n_1114),
.B1(n_1231),
.B2(n_1232),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1209),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1203),
.A2(n_1217),
.B1(n_1119),
.B2(n_1125),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1156),
.Y(n_1245)
);

INVx6_ASAP7_75t_L g1246 ( 
.A(n_1116),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1179),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1132),
.Y(n_1248)
);

CKINVDCx6p67_ASAP7_75t_R g1249 ( 
.A(n_1190),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1220),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1175),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1114),
.A2(n_1207),
.B1(n_1184),
.B2(n_1231),
.Y(n_1252)
);

INVxp67_ASAP7_75t_SL g1253 ( 
.A(n_1139),
.Y(n_1253)
);

CKINVDCx16_ASAP7_75t_R g1254 ( 
.A(n_1193),
.Y(n_1254)
);

CKINVDCx6p67_ASAP7_75t_R g1255 ( 
.A(n_1205),
.Y(n_1255)
);

INVx5_ASAP7_75t_L g1256 ( 
.A(n_1192),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1220),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1184),
.A2(n_1207),
.B1(n_1232),
.B2(n_1130),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1104),
.A2(n_1201),
.B1(n_1218),
.B2(n_1174),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_1169),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1130),
.A2(n_1234),
.B1(n_1213),
.B2(n_1107),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1115),
.A2(n_1167),
.B1(n_1234),
.B2(n_1107),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1104),
.A2(n_1180),
.B1(n_1201),
.B2(n_1218),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1189),
.Y(n_1264)
);

NAND2x1p5_ASAP7_75t_L g1265 ( 
.A(n_1151),
.B(n_1224),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1174),
.A2(n_1180),
.B1(n_1126),
.B2(n_1117),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1144),
.Y(n_1267)
);

BUFx2_ASAP7_75t_R g1268 ( 
.A(n_1171),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1177),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1155),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1117),
.A2(n_1108),
.B1(n_1127),
.B2(n_1195),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1191),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1115),
.A2(n_1167),
.B1(n_1178),
.B2(n_1139),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1177),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1212),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1116),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1118),
.Y(n_1277)
);

OAI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1181),
.A2(n_1147),
.B1(n_1138),
.B2(n_1200),
.Y(n_1278)
);

BUFx4f_ASAP7_75t_L g1279 ( 
.A(n_1116),
.Y(n_1279)
);

INVx6_ASAP7_75t_L g1280 ( 
.A(n_1149),
.Y(n_1280)
);

CKINVDCx11_ASAP7_75t_R g1281 ( 
.A(n_1187),
.Y(n_1281)
);

INVx5_ASAP7_75t_SL g1282 ( 
.A(n_1149),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1214),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1208),
.A2(n_1135),
.B1(n_1168),
.B2(n_1145),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1147),
.B(n_1157),
.Y(n_1285)
);

INVx6_ASAP7_75t_L g1286 ( 
.A(n_1182),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1158),
.Y(n_1287)
);

CKINVDCx11_ASAP7_75t_R g1288 ( 
.A(n_1192),
.Y(n_1288)
);

INVx6_ASAP7_75t_L g1289 ( 
.A(n_1182),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1185),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1178),
.A2(n_1157),
.B1(n_1128),
.B2(n_1121),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1153),
.A2(n_1133),
.B1(n_1122),
.B2(n_1176),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1224),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1158),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1160),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1233),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1160),
.Y(n_1297)
);

OAI21xp33_ASAP7_75t_L g1298 ( 
.A1(n_1105),
.A2(n_1143),
.B(n_1129),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1134),
.A2(n_1102),
.B1(n_1120),
.B2(n_1113),
.Y(n_1299)
);

CKINVDCx8_ASAP7_75t_R g1300 ( 
.A(n_1128),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1102),
.A2(n_1150),
.B1(n_1154),
.B2(n_1159),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1163),
.A2(n_1233),
.B1(n_1161),
.B2(n_1136),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1162),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1177),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1176),
.B(n_1166),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1124),
.A2(n_1141),
.B(n_1109),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1166),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1165),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1150),
.A2(n_1112),
.B1(n_1164),
.B2(n_1111),
.Y(n_1309)
);

CKINVDCx6p67_ASAP7_75t_R g1310 ( 
.A(n_1165),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1206),
.Y(n_1311)
);

BUFx2_ASAP7_75t_SL g1312 ( 
.A(n_1148),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1206),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1137),
.A2(n_1146),
.B1(n_1152),
.B2(n_1225),
.Y(n_1314)
);

INVx6_ASAP7_75t_L g1315 ( 
.A(n_1165),
.Y(n_1315)
);

BUFx8_ASAP7_75t_SL g1316 ( 
.A(n_1210),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1197),
.A2(n_1215),
.B1(n_1110),
.B2(n_1202),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1197),
.A2(n_1215),
.B1(n_1216),
.B2(n_1228),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1197),
.Y(n_1319)
);

OAI21xp33_ASAP7_75t_L g1320 ( 
.A1(n_1229),
.A2(n_1235),
.B(n_1215),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1140),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1140),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1142),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1103),
.A2(n_1219),
.B1(n_1198),
.B2(n_1173),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1186),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1170),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1106),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1172),
.A2(n_1194),
.B1(n_1199),
.B2(n_1211),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1221),
.A2(n_1222),
.B1(n_1223),
.B2(n_1227),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1188),
.A2(n_1226),
.B1(n_1217),
.B2(n_1203),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1209),
.Y(n_1331)
);

INVx6_ASAP7_75t_L g1332 ( 
.A(n_1116),
.Y(n_1332)
);

BUFx8_ASAP7_75t_SL g1333 ( 
.A(n_1193),
.Y(n_1333)
);

NAND2x1p5_ASAP7_75t_L g1334 ( 
.A(n_1151),
.B(n_1233),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1188),
.A2(n_1226),
.B1(n_1217),
.B2(n_1203),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1188),
.B(n_1226),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1116),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1179),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1209),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1179),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1196),
.A2(n_1226),
.B1(n_1188),
.B2(n_988),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1209),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1179),
.Y(n_1343)
);

BUFx4f_ASAP7_75t_SL g1344 ( 
.A(n_1205),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1188),
.A2(n_1226),
.B1(n_1217),
.B2(n_1203),
.Y(n_1345)
);

CKINVDCx6p67_ASAP7_75t_R g1346 ( 
.A(n_1190),
.Y(n_1346)
);

BUFx12f_ASAP7_75t_L g1347 ( 
.A(n_1209),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1196),
.A2(n_591),
.B1(n_430),
.B2(n_1114),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1326),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1322),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1252),
.B(n_1242),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1341),
.A2(n_1335),
.B(n_1330),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1247),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1306),
.A2(n_1324),
.B(n_1329),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1269),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1308),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1345),
.A2(n_1244),
.B1(n_1336),
.B2(n_1319),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1314),
.A2(n_1320),
.B(n_1323),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1338),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1274),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1266),
.B(n_1259),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1274),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1304),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1311),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1340),
.Y(n_1365)
);

BUFx2_ASAP7_75t_SL g1366 ( 
.A(n_1238),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1313),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1252),
.B(n_1242),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1324),
.A2(n_1329),
.B(n_1309),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1250),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1263),
.B(n_1271),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1316),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1265),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1321),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1325),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1253),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1261),
.B(n_1258),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1327),
.Y(n_1378)
);

AO21x1_ASAP7_75t_SL g1379 ( 
.A1(n_1258),
.A2(n_1298),
.B(n_1284),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1341),
.A2(n_1236),
.B1(n_1348),
.B2(n_1262),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1236),
.A2(n_1348),
.B1(n_1262),
.B2(n_1273),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1301),
.B(n_1295),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1287),
.B(n_1294),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1253),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1285),
.B(n_1305),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1309),
.A2(n_1299),
.B(n_1318),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1257),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1247),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1297),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1248),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1343),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1316),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1251),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1291),
.A2(n_1302),
.B(n_1299),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1291),
.A2(n_1292),
.B(n_1278),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1264),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1272),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1326),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1241),
.Y(n_1399)
);

INVx5_ASAP7_75t_L g1400 ( 
.A(n_1315),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1315),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1343),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1265),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1301),
.B(n_1240),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1334),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1273),
.B(n_1237),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1275),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1334),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1278),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1246),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1303),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1317),
.B(n_1318),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1276),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1310),
.Y(n_1414)
);

CKINVDCx14_ASAP7_75t_R g1415 ( 
.A(n_1243),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1246),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1277),
.B(n_1254),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1317),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1284),
.A2(n_1267),
.B(n_1270),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1293),
.A2(n_1328),
.B(n_1296),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1307),
.A2(n_1290),
.B(n_1293),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_1246),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1332),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1312),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1337),
.B(n_1276),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1332),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1280),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1238),
.A2(n_1256),
.B(n_1282),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1249),
.A2(n_1346),
.B1(n_1255),
.B2(n_1281),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1352),
.A2(n_1279),
.B(n_1283),
.C(n_1256),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1403),
.B(n_1256),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1403),
.B(n_1342),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1385),
.B(n_1280),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1405),
.B(n_1339),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1380),
.A2(n_1279),
.B(n_1245),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_SL g1436 ( 
.A1(n_1395),
.A2(n_1371),
.B(n_1361),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1394),
.A2(n_1331),
.B(n_1268),
.Y(n_1437)
);

AND2x6_ASAP7_75t_L g1438 ( 
.A(n_1401),
.B(n_1288),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1370),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1363),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1385),
.B(n_1239),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1376),
.B(n_1239),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1357),
.A2(n_1300),
.B(n_1333),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1411),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1356),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1386),
.B(n_1347),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1418),
.B(n_1288),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1418),
.B(n_1286),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1417),
.B(n_1333),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1387),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1356),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1419),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1404),
.B(n_1286),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1386),
.A2(n_1289),
.B(n_1281),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1376),
.B(n_1260),
.Y(n_1455)
);

AO21x1_ASAP7_75t_L g1456 ( 
.A1(n_1409),
.A2(n_1289),
.B(n_1260),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1404),
.B(n_1344),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1383),
.B(n_1344),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1419),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1381),
.A2(n_1372),
.B1(n_1392),
.B2(n_1368),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1351),
.A2(n_1368),
.B(n_1424),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1382),
.B(n_1412),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1382),
.B(n_1412),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1409),
.A2(n_1351),
.B1(n_1377),
.B2(n_1407),
.C(n_1382),
.Y(n_1464)
);

INVx4_ASAP7_75t_L g1465 ( 
.A(n_1428),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1383),
.B(n_1359),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1382),
.B(n_1406),
.Y(n_1467)
);

AO22x2_ASAP7_75t_L g1468 ( 
.A1(n_1374),
.A2(n_1360),
.B1(n_1355),
.B2(n_1362),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1390),
.B(n_1393),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1367),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1365),
.B(n_1399),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1415),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1367),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1354),
.A2(n_1369),
.B(n_1420),
.Y(n_1474)
);

AOI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1377),
.A2(n_1421),
.B1(n_1391),
.B2(n_1388),
.C(n_1402),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1396),
.B(n_1397),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1369),
.A2(n_1420),
.B(n_1364),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1353),
.Y(n_1478)
);

A2O1A1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1372),
.A2(n_1392),
.B(n_1379),
.C(n_1424),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1405),
.B(n_1408),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1349),
.A2(n_1398),
.B(n_1429),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1429),
.A2(n_1414),
.B1(n_1423),
.B2(n_1422),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1379),
.A2(n_1414),
.B(n_1349),
.C(n_1398),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1468),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1462),
.B(n_1384),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1468),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1440),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1436),
.A2(n_1349),
.B1(n_1398),
.B2(n_1427),
.Y(n_1488)
);

AND2x4_ASAP7_75t_SL g1489 ( 
.A(n_1431),
.B(n_1373),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1442),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1470),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1467),
.B(n_1378),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1480),
.B(n_1408),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1467),
.B(n_1378),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1462),
.B(n_1375),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1460),
.A2(n_1435),
.B1(n_1437),
.B2(n_1464),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1463),
.B(n_1469),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1452),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1440),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1473),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1444),
.B(n_1389),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1436),
.A2(n_1366),
.B1(n_1419),
.B2(n_1400),
.Y(n_1502)
);

INVxp67_ASAP7_75t_SL g1503 ( 
.A(n_1459),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1477),
.B(n_1358),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1477),
.B(n_1358),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1477),
.B(n_1358),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1477),
.B(n_1350),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1474),
.B(n_1350),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1457),
.A2(n_1349),
.B1(n_1398),
.B2(n_1427),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1468),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1441),
.B(n_1422),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1468),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1461),
.A2(n_1366),
.B1(n_1419),
.B2(n_1400),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1476),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1445),
.B(n_1360),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1496),
.B(n_1434),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1491),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1497),
.B(n_1490),
.Y(n_1518)
);

NAND3xp33_ASAP7_75t_L g1519 ( 
.A(n_1496),
.B(n_1475),
.C(n_1437),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1507),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1502),
.A2(n_1430),
.B(n_1483),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1490),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1497),
.B(n_1446),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1512),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1484),
.A2(n_1450),
.B1(n_1439),
.B2(n_1471),
.C(n_1466),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1484),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1507),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1495),
.B(n_1455),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1487),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1512),
.B(n_1486),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1486),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1508),
.Y(n_1532)
);

NOR2xp67_ASAP7_75t_L g1533 ( 
.A(n_1510),
.B(n_1465),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1510),
.Y(n_1534)
);

OAI31xp33_ASAP7_75t_L g1535 ( 
.A1(n_1488),
.A2(n_1479),
.A3(n_1482),
.B(n_1457),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1487),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1513),
.A2(n_1443),
.B1(n_1481),
.B2(n_1446),
.C(n_1455),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1499),
.Y(n_1538)
);

INVx4_ASAP7_75t_L g1539 ( 
.A(n_1489),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1492),
.B(n_1446),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1494),
.B(n_1446),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1489),
.Y(n_1542)
);

AOI211xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1511),
.A2(n_1449),
.B(n_1447),
.C(n_1448),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1485),
.B(n_1451),
.Y(n_1544)
);

INVx4_ASAP7_75t_L g1545 ( 
.A(n_1489),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1515),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1499),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1508),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1493),
.B(n_1465),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1500),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1500),
.Y(n_1551)
);

NAND4xp25_ASAP7_75t_L g1552 ( 
.A(n_1513),
.B(n_1458),
.C(n_1447),
.D(n_1442),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1530),
.B(n_1454),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1520),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1539),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1526),
.B(n_1498),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1550),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1530),
.B(n_1454),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1527),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_L g1560 ( 
.A(n_1519),
.B(n_1502),
.C(n_1472),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1530),
.B(n_1454),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1527),
.B(n_1504),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1527),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1530),
.B(n_1454),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1519),
.B(n_1516),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1529),
.Y(n_1566)
);

OAI211xp5_ASAP7_75t_L g1567 ( 
.A1(n_1535),
.A2(n_1498),
.B(n_1503),
.C(n_1433),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1532),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1550),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1531),
.B(n_1503),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1532),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1529),
.Y(n_1572)
);

INVxp67_ASAP7_75t_SL g1573 ( 
.A(n_1534),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1536),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1536),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1549),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1551),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1524),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1548),
.B(n_1505),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1546),
.B(n_1514),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1551),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1524),
.B(n_1515),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1548),
.B(n_1506),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1517),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1576),
.B(n_1523),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1565),
.B(n_1472),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1578),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1578),
.Y(n_1588)
);

OAI32xp33_ASAP7_75t_L g1589 ( 
.A1(n_1565),
.A2(n_1552),
.A3(n_1537),
.B1(n_1522),
.B2(n_1546),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1578),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1578),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1555),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1573),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1566),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1567),
.B(n_1525),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1566),
.Y(n_1596)
);

NAND2x1p5_ASAP7_75t_L g1597 ( 
.A(n_1555),
.B(n_1539),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1572),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1567),
.B(n_1543),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1559),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1572),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1573),
.B(n_1522),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1560),
.B(n_1543),
.Y(n_1603)
);

NOR2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1560),
.B(n_1552),
.Y(n_1604)
);

NOR4xp25_ASAP7_75t_SL g1605 ( 
.A(n_1555),
.B(n_1535),
.C(n_1538),
.D(n_1547),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1574),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1576),
.B(n_1523),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1555),
.B(n_1533),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1574),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1584),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1575),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1555),
.B(n_1521),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1553),
.A2(n_1456),
.B1(n_1438),
.B2(n_1453),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1575),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1576),
.B(n_1540),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1576),
.B(n_1540),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1582),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1576),
.B(n_1541),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1557),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1580),
.B(n_1518),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1557),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1559),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1559),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1556),
.B(n_1544),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1584),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1557),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1587),
.Y(n_1627)
);

NOR3xp33_ASAP7_75t_L g1628 ( 
.A(n_1589),
.B(n_1432),
.C(n_1478),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1585),
.B(n_1553),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1619),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1604),
.B(n_1553),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1604),
.B(n_1558),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1617),
.B(n_1556),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1599),
.B(n_1603),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1602),
.B(n_1556),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1595),
.B(n_1558),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1585),
.B(n_1558),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1587),
.B(n_1561),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1620),
.B(n_1528),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1619),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1621),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1602),
.B(n_1582),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_SL g1643 ( 
.A1(n_1612),
.A2(n_1564),
.B(n_1561),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1607),
.B(n_1561),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1621),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1593),
.B(n_1564),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1624),
.B(n_1582),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1588),
.B(n_1591),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1622),
.Y(n_1649)
);

OAI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1613),
.A2(n_1539),
.B1(n_1545),
.B2(n_1542),
.Y(n_1650)
);

AND2x4_ASAP7_75t_SL g1651 ( 
.A(n_1608),
.B(n_1539),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1626),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1588),
.B(n_1564),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1591),
.B(n_1518),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1586),
.A2(n_1456),
.B1(n_1474),
.B2(n_1506),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1624),
.B(n_1570),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1605),
.B(n_1509),
.C(n_1570),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1622),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1626),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1590),
.A2(n_1584),
.B(n_1568),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1597),
.Y(n_1661)
);

AOI211x1_ASAP7_75t_L g1662 ( 
.A1(n_1634),
.A2(n_1589),
.B(n_1607),
.C(n_1615),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1651),
.B(n_1615),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1631),
.A2(n_1592),
.B1(n_1590),
.B2(n_1597),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1627),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1634),
.B(n_1432),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1628),
.A2(n_1613),
.B(n_1592),
.C(n_1608),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1632),
.A2(n_1616),
.B1(n_1618),
.B2(n_1608),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1636),
.A2(n_1597),
.B(n_1590),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_L g1670 ( 
.A(n_1657),
.B(n_1596),
.C(n_1594),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1643),
.A2(n_1655),
.B(n_1650),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1639),
.B(n_1432),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1630),
.Y(n_1673)
);

OAI21xp33_ASAP7_75t_L g1674 ( 
.A1(n_1655),
.A2(n_1618),
.B(n_1616),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1648),
.B(n_1608),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1650),
.B(n_1542),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1661),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1651),
.A2(n_1542),
.B1(n_1545),
.B2(n_1533),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1635),
.B(n_1594),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1654),
.A2(n_1545),
.B1(n_1542),
.B2(n_1549),
.Y(n_1680)
);

AOI222xp33_ASAP7_75t_L g1681 ( 
.A1(n_1646),
.A2(n_1596),
.B1(n_1611),
.B2(n_1609),
.C1(n_1606),
.C2(n_1601),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1633),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1638),
.Y(n_1683)
);

OAI31xp33_ASAP7_75t_L g1684 ( 
.A1(n_1633),
.A2(n_1622),
.A3(n_1623),
.B(n_1570),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1635),
.B(n_1642),
.Y(n_1685)
);

OAI211xp5_ASAP7_75t_L g1686 ( 
.A1(n_1653),
.A2(n_1601),
.B(n_1606),
.C(n_1609),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1665),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1671),
.A2(n_1656),
.B1(n_1647),
.B2(n_1652),
.C(n_1659),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1682),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1677),
.B(n_1682),
.Y(n_1690)
);

XNOR2x1_ASAP7_75t_L g1691 ( 
.A(n_1670),
.B(n_1434),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1666),
.B(n_1638),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1673),
.Y(n_1693)
);

O2A1O1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1667),
.A2(n_1645),
.B(n_1640),
.C(n_1641),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_SL g1695 ( 
.A(n_1664),
.B(n_1658),
.C(n_1649),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_R g1696 ( 
.A(n_1685),
.B(n_1434),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1679),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1676),
.A2(n_1638),
.B1(n_1629),
.B2(n_1637),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1664),
.A2(n_1658),
.B(n_1649),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1662),
.B(n_1629),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1683),
.Y(n_1701)
);

AOI21xp33_ASAP7_75t_L g1702 ( 
.A1(n_1675),
.A2(n_1611),
.B(n_1598),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1672),
.B(n_1637),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1668),
.A2(n_1644),
.B1(n_1545),
.B2(n_1622),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1675),
.B(n_1644),
.Y(n_1705)
);

AOI211x1_ASAP7_75t_L g1706 ( 
.A1(n_1688),
.A2(n_1669),
.B(n_1674),
.C(n_1686),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1695),
.A2(n_1681),
.B(n_1663),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1696),
.B(n_1684),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1687),
.B(n_1680),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1698),
.A2(n_1678),
.B1(n_1623),
.B2(n_1600),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1690),
.B(n_1598),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1689),
.B(n_1614),
.Y(n_1712)
);

OAI21xp33_ASAP7_75t_SL g1713 ( 
.A1(n_1700),
.A2(n_1623),
.B(n_1600),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1692),
.B(n_1623),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1704),
.A2(n_1691),
.B1(n_1705),
.B2(n_1701),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_SL g1716 ( 
.A(n_1697),
.B(n_1600),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1703),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1717),
.B(n_1693),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1711),
.Y(n_1719)
);

AOI222xp33_ASAP7_75t_L g1720 ( 
.A1(n_1707),
.A2(n_1699),
.B1(n_1694),
.B2(n_1702),
.C1(n_1614),
.C2(n_1625),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1709),
.Y(n_1721)
);

AOI211xp5_ASAP7_75t_L g1722 ( 
.A1(n_1708),
.A2(n_1699),
.B(n_1625),
.C(n_1610),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1706),
.B(n_1569),
.Y(n_1723)
);

NAND4xp75_ASAP7_75t_L g1724 ( 
.A(n_1713),
.B(n_1715),
.C(n_1714),
.D(n_1712),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1716),
.Y(n_1725)
);

NOR3xp33_ASAP7_75t_SL g1726 ( 
.A(n_1710),
.B(n_1580),
.C(n_1501),
.Y(n_1726)
);

AOI211x1_ASAP7_75t_SL g1727 ( 
.A1(n_1723),
.A2(n_1610),
.B(n_1554),
.C(n_1571),
.Y(n_1727)
);

OAI21xp33_ASAP7_75t_SL g1728 ( 
.A1(n_1720),
.A2(n_1583),
.B(n_1579),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1718),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1725),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1721),
.B(n_1569),
.Y(n_1731)
);

AOI221x1_ASAP7_75t_SL g1732 ( 
.A1(n_1730),
.A2(n_1722),
.B1(n_1719),
.B2(n_1724),
.C(n_1726),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1729),
.Y(n_1733)
);

NOR2xp67_ASAP7_75t_L g1734 ( 
.A(n_1731),
.B(n_1722),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1727),
.B(n_1660),
.Y(n_1735)
);

XNOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1728),
.B(n_1425),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_L g1737 ( 
.A(n_1729),
.B(n_1423),
.C(n_1426),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1733),
.B(n_1559),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1734),
.Y(n_1739)
);

AO22x2_ASAP7_75t_L g1740 ( 
.A1(n_1732),
.A2(n_1584),
.B1(n_1571),
.B2(n_1568),
.Y(n_1740)
);

XNOR2xp5_ASAP7_75t_L g1741 ( 
.A(n_1736),
.B(n_1737),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1735),
.B(n_1660),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1740),
.A2(n_1581),
.B1(n_1577),
.B2(n_1569),
.C(n_1571),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_L g1744 ( 
.A(n_1739),
.B(n_1741),
.C(n_1742),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1740),
.B(n_1660),
.Y(n_1745)
);

AO22x2_ASAP7_75t_L g1746 ( 
.A1(n_1744),
.A2(n_1738),
.B1(n_1741),
.B2(n_1581),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1745),
.B1(n_1743),
.B2(n_1568),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1747),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1748),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1749),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1562),
.B1(n_1554),
.B2(n_1568),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1750),
.A2(n_1554),
.B1(n_1563),
.B2(n_1571),
.Y(n_1752)
);

OR2x6_ASAP7_75t_L g1753 ( 
.A(n_1752),
.B(n_1425),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1751),
.A2(n_1563),
.B1(n_1554),
.B2(n_1581),
.Y(n_1754)
);

OAI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1753),
.A2(n_1563),
.B1(n_1577),
.B2(n_1413),
.Y(n_1755)
);

XNOR2xp5_ASAP7_75t_L g1756 ( 
.A(n_1754),
.B(n_1425),
.Y(n_1756)
);

AOI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1755),
.A2(n_1577),
.B1(n_1563),
.B2(n_1562),
.C(n_1559),
.Y(n_1757)
);

OAI31xp33_ASAP7_75t_L g1758 ( 
.A1(n_1757),
.A2(n_1756),
.A3(n_1410),
.B(n_1416),
.Y(n_1758)
);


endmodule