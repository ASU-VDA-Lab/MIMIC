module fake_jpeg_2109_n_683 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_683);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_683;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_4),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_59),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_63),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g222 ( 
.A(n_64),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_65),
.B(n_95),
.Y(n_194)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_32),
.B(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_68),
.B(n_71),
.Y(n_137)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g212 ( 
.A(n_69),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_29),
.B(n_18),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_72),
.B(n_98),
.Y(n_149)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g192 ( 
.A(n_75),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_79),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_82),
.Y(n_214)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_85),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_87),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_89),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_32),
.B(n_16),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_100),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_48),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx11_ASAP7_75t_SL g110 ( 
.A(n_21),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_126),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_31),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_117),
.Y(n_225)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_118),
.Y(n_217)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_123),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_33),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_124),
.B(n_35),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_47),
.B(n_16),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_127),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_21),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_33),
.B(n_15),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_41),
.Y(n_131)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_43),
.B(n_53),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_134),
.B(n_170),
.C(n_193),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_113),
.A2(n_21),
.B1(n_37),
.B2(n_128),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_161),
.A2(n_26),
.B1(n_102),
.B2(n_96),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_104),
.B(n_43),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_166),
.B(n_181),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_168),
.Y(n_296)
);

OR2x2_ASAP7_75t_SL g170 ( 
.A(n_85),
.B(n_56),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_64),
.B(n_23),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_174),
.B(n_177),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_64),
.B(n_23),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_101),
.B(n_57),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_89),
.B(n_57),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_185),
.B(n_186),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_107),
.B(n_45),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_116),
.B(n_22),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_188),
.B(n_190),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_60),
.B(n_22),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_107),
.B(n_38),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_191),
.B(n_196),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_122),
.B(n_56),
.C(n_28),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_125),
.B(n_45),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_61),
.B(n_28),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_197),
.B(n_200),
.Y(n_312)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_67),
.A2(n_41),
.B1(n_37),
.B2(n_31),
.Y(n_198)
);

AO22x2_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_209),
.B1(n_173),
.B2(n_140),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_62),
.B(n_40),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_127),
.B(n_40),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_204),
.B(n_208),
.Y(n_315)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_85),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_206),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_75),
.B(n_39),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_207),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_99),
.B(n_39),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_63),
.A2(n_37),
.B1(n_38),
.B2(n_35),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_209),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_218),
.Y(n_233)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_92),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_213),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_70),
.B(n_34),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_216),
.B(n_223),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_121),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_79),
.B(n_26),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_220),
.B(n_14),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_82),
.B(n_34),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_84),
.Y(n_224)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_87),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_117),
.Y(n_235)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_90),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_231),
.Y(n_232)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_151),
.Y(n_234)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_234),
.Y(n_328)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_235),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_236),
.B(n_278),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_138),
.Y(n_237)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_237),
.Y(n_335)
);

OR2x2_ASAP7_75t_SL g238 ( 
.A(n_154),
.B(n_41),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_238),
.B(n_204),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_114),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_239),
.Y(n_358)
);

CKINVDCx12_ASAP7_75t_R g240 ( 
.A(n_228),
.Y(n_240)
);

INVx4_ASAP7_75t_SL g373 ( 
.A(n_240),
.Y(n_373)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_139),
.Y(n_242)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_242),
.Y(n_331)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_138),
.Y(n_244)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_244),
.Y(n_364)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_245),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_246),
.A2(n_285),
.B1(n_303),
.B2(n_305),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_155),
.Y(n_247)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_247),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_169),
.B(n_15),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_249),
.B(n_252),
.Y(n_322)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_151),
.Y(n_250)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_250),
.Y(n_338)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_152),
.Y(n_251)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_251),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_169),
.B(n_15),
.Y(n_252)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_144),
.Y(n_253)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_253),
.Y(n_366)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_136),
.Y(n_255)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_255),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_194),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_256),
.B(n_275),
.Y(n_356)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_257),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_161),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_258),
.B(n_277),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_149),
.B(n_106),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_259),
.B(n_270),
.Y(n_375)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_262),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_208),
.A2(n_91),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_263),
.A2(n_289),
.B1(n_298),
.B2(n_210),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_162),
.Y(n_264)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_264),
.Y(n_361)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_141),
.Y(n_265)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_265),
.Y(n_368)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

BUFx24_ASAP7_75t_L g365 ( 
.A(n_266),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_267),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_146),
.Y(n_269)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_269),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_149),
.B(n_0),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_163),
.Y(n_271)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_271),
.Y(n_354)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_272),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_146),
.Y(n_273)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_274),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_145),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_172),
.Y(n_276)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_276),
.Y(n_378)
);

INVx3_ASAP7_75t_SL g278 ( 
.A(n_212),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_179),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_279),
.B(n_286),
.Y(n_377)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_167),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_283),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_154),
.B(n_1),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_281),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_137),
.B(n_1),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_282),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_221),
.B(n_1),
.Y(n_283)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_179),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_171),
.Y(n_286)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_165),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_287),
.Y(n_330)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_199),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_288),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_220),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_289)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_165),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_290),
.Y(n_332)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_222),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_291),
.Y(n_380)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_148),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_293),
.Y(n_343)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_199),
.Y(n_293)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_222),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_294),
.Y(n_344)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_160),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_295),
.B(n_297),
.Y(n_346)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_201),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_137),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_299),
.A2(n_219),
.B1(n_175),
.B2(n_203),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_186),
.B(n_7),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_301),
.A2(n_306),
.B1(n_308),
.B2(n_317),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_145),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_302),
.Y(n_360)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_133),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_156),
.Y(n_304)
);

NOR2x1_ASAP7_75t_L g339 ( 
.A(n_304),
.B(n_314),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_219),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_191),
.B(n_8),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_164),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_310),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_198),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_185),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_196),
.B(n_10),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_316),
.Y(n_345)
);

CKINVDCx12_ASAP7_75t_R g314 ( 
.A(n_176),
.Y(n_314)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_184),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_174),
.B(n_10),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_198),
.A2(n_12),
.B1(n_13),
.B2(n_181),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_318),
.A2(n_177),
.B1(n_192),
.B2(n_135),
.Y(n_342)
);

AO21x1_ASAP7_75t_L g384 ( 
.A1(n_325),
.A2(n_281),
.B(n_282),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_143),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_340),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_261),
.B(n_132),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_342),
.A2(n_349),
.B1(n_350),
.B2(n_362),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_318),
.A2(n_153),
.B1(n_147),
.B2(n_192),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_243),
.A2(n_189),
.B1(n_214),
.B2(n_180),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_260),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_355),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_353),
.A2(n_371),
.B1(n_379),
.B2(n_278),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_284),
.B(n_230),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_248),
.B(n_217),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_266),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_308),
.A2(n_189),
.B1(n_202),
.B2(n_225),
.Y(n_362)
);

OAI32xp33_ASAP7_75t_L g363 ( 
.A1(n_239),
.A2(n_173),
.A3(n_212),
.B1(n_195),
.B2(n_142),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_266),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_258),
.A2(n_277),
.B(n_309),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_271),
.B(n_296),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_236),
.A2(n_195),
.B1(n_227),
.B2(n_150),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_L g381 ( 
.A1(n_337),
.A2(n_246),
.B1(n_236),
.B2(n_263),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_381),
.A2(n_386),
.B1(n_392),
.B2(n_403),
.Y(n_437)
);

AND2x2_ASAP7_75t_SL g382 ( 
.A(n_358),
.B(n_238),
.Y(n_382)
);

NAND2x1_ASAP7_75t_SL g458 ( 
.A(n_382),
.B(n_415),
.Y(n_458)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

AO21x1_ASAP7_75t_L g435 ( 
.A1(n_384),
.A2(n_389),
.B(n_395),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_385),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_299),
.B1(n_236),
.B2(n_268),
.Y(n_386)
);

BUFx16f_ASAP7_75t_L g387 ( 
.A(n_380),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_387),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_377),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_388),
.B(n_397),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_321),
.A2(n_337),
.B1(n_358),
.B2(n_342),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_371),
.A2(n_239),
.B1(n_233),
.B2(n_157),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_351),
.B(n_241),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_393),
.B(n_414),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_327),
.A2(n_303),
.B1(n_232),
.B2(n_273),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g450 ( 
.A1(n_394),
.A2(n_409),
.B1(n_424),
.B2(n_427),
.Y(n_450)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_396),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_373),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_335),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_398),
.Y(n_438)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_328),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_399),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_377),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_400),
.B(n_406),
.Y(n_464)
);

INVx13_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_401),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_402),
.B(n_412),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_355),
.A2(n_182),
.B1(n_210),
.B2(n_178),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_347),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_404),
.B(n_405),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_356),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_377),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g408 ( 
.A(n_325),
.B(n_294),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_408),
.B(n_411),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_373),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_327),
.B(n_290),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_413),
.A2(n_296),
.B(n_365),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_375),
.B(n_264),
.Y(n_414)
);

NAND2x1_ASAP7_75t_SL g415 ( 
.A(n_354),
.B(n_291),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_416),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_345),
.B(n_253),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_417),
.B(n_419),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_339),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_418),
.B(n_421),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_346),
.Y(n_419)
);

INVx6_ASAP7_75t_L g420 ( 
.A(n_330),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_420),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_326),
.B(n_300),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_329),
.B(n_311),
.Y(n_422)
);

MAJx2_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_378),
.C(n_352),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_328),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_423),
.B(n_426),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_357),
.A2(n_287),
.B1(n_244),
.B2(n_237),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_345),
.B(n_323),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_425),
.B(n_428),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_340),
.B(n_305),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_364),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_360),
.B(n_311),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_322),
.B(n_247),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_429),
.B(n_430),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_331),
.B(n_341),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_386),
.A2(n_319),
.B1(n_370),
.B2(n_374),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_433),
.A2(n_442),
.B1(n_456),
.B2(n_468),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_395),
.A2(n_362),
.B1(n_336),
.B2(n_319),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_436),
.A2(n_446),
.B(n_448),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_381),
.A2(n_349),
.B1(n_350),
.B2(n_334),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_367),
.C(n_372),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_443),
.B(n_385),
.C(n_419),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_413),
.A2(n_363),
.B(n_339),
.Y(n_446)
);

OAI22xp33_ASAP7_75t_L g447 ( 
.A1(n_407),
.A2(n_332),
.B1(n_344),
.B2(n_324),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_447),
.A2(n_390),
.B1(n_383),
.B2(n_396),
.Y(n_502)
);

A2O1A1Ixp33_ASAP7_75t_SL g449 ( 
.A1(n_395),
.A2(n_365),
.B(n_324),
.C(n_333),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_449),
.A2(n_453),
.B(n_461),
.Y(n_483)
);

XNOR2x1_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_422),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_389),
.A2(n_368),
.B(n_369),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_392),
.A2(n_333),
.B1(n_364),
.B2(n_376),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_387),
.Y(n_459)
);

INVx13_ASAP7_75t_L g480 ( 
.A(n_459),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_402),
.A2(n_368),
.B1(n_338),
.B2(n_320),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_460),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_406),
.A2(n_348),
.B(n_359),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_387),
.Y(n_462)
);

INVx13_ASAP7_75t_L g486 ( 
.A(n_462),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_415),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_382),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_407),
.A2(n_335),
.B1(n_369),
.B2(n_359),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_405),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_473),
.B(n_485),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_455),
.Y(n_474)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_474),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_471),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_475),
.B(n_459),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_451),
.B(n_410),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g550 ( 
.A(n_476),
.B(n_481),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_391),
.Y(n_477)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_477),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_437),
.A2(n_436),
.B1(n_442),
.B2(n_463),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_478),
.A2(n_494),
.B1(n_495),
.B2(n_446),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_479),
.B(n_503),
.Y(n_515)
);

OAI21xp33_ASAP7_75t_SL g540 ( 
.A1(n_482),
.A2(n_506),
.B(n_458),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_425),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_431),
.B(n_391),
.Y(n_488)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_431),
.B(n_417),
.Y(n_489)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_489),
.Y(n_520)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_467),
.Y(n_490)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_490),
.Y(n_521)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_445),
.Y(n_491)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_491),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_492),
.B(n_496),
.C(n_454),
.Y(n_527)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_467),
.Y(n_493)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_493),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_437),
.A2(n_412),
.B1(n_382),
.B2(n_408),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_465),
.A2(n_426),
.B1(n_400),
.B2(n_423),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_443),
.B(n_384),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_445),
.Y(n_497)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_441),
.B(n_404),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_498),
.B(n_507),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_466),
.A2(n_415),
.B(n_384),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_499),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_435),
.B(n_403),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_500),
.B(n_435),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_465),
.B(n_420),
.Y(n_501)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_501),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_502),
.A2(n_505),
.B1(n_450),
.B2(n_444),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_432),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_455),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_504),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_456),
.A2(n_399),
.B1(n_427),
.B2(n_398),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_458),
.B(n_416),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_439),
.B(n_361),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_444),
.B(n_398),
.Y(n_508)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_457),
.Y(n_509)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_509),
.Y(n_549)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_472),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_512),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_432),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_513),
.A2(n_528),
.B1(n_542),
.B2(n_511),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_439),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_514),
.B(n_532),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_464),
.Y(n_518)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_518),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_523),
.B(n_527),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_489),
.B(n_441),
.Y(n_524)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_524),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_477),
.B(n_449),
.Y(n_525)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_525),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_449),
.Y(n_526)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_526),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_484),
.A2(n_470),
.B1(n_433),
.B2(n_469),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_530),
.A2(n_511),
.B1(n_483),
.B2(n_506),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_479),
.A2(n_435),
.B(n_453),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_531),
.A2(n_536),
.B(n_499),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_474),
.B(n_434),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_495),
.Y(n_533)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_533),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_494),
.B(n_469),
.Y(n_535)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_535),
.Y(n_552)
);

A2O1A1O1Ixp25_ASAP7_75t_L g536 ( 
.A1(n_482),
.A2(n_458),
.B(n_461),
.C(n_449),
.D(n_462),
.Y(n_536)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_537),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_540),
.B(n_440),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_503),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_496),
.B(n_460),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_478),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_512),
.B(n_432),
.Y(n_548)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_548),
.Y(n_555)
);

AOI21x1_ASAP7_75t_L g588 ( 
.A1(n_551),
.A2(n_577),
.B(n_515),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_554),
.B(n_580),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_544),
.A2(n_487),
.B(n_482),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_556),
.A2(n_579),
.B(n_536),
.Y(n_596)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_518),
.Y(n_557)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_557),
.Y(n_586)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_549),
.Y(n_558)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_558),
.Y(n_603)
);

AOI21xp33_ASAP7_75t_L g561 ( 
.A1(n_538),
.A2(n_487),
.B(n_506),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_561),
.B(n_574),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_527),
.B(n_476),
.C(n_481),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_562),
.B(n_573),
.C(n_575),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_564),
.A2(n_544),
.B1(n_546),
.B2(n_525),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_566),
.A2(n_559),
.B1(n_577),
.B2(n_576),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_533),
.A2(n_500),
.B1(n_483),
.B2(n_502),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_567),
.A2(n_570),
.B1(n_546),
.B2(n_526),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_531),
.A2(n_449),
.B(n_486),
.Y(n_568)
);

CKINVDCx14_ASAP7_75t_R g593 ( 
.A(n_568),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_542),
.B(n_510),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_569),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_543),
.A2(n_468),
.B1(n_504),
.B2(n_490),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_516),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_571),
.B(n_578),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_545),
.B(n_457),
.C(n_338),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_538),
.B(n_440),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_550),
.B(n_472),
.C(n_486),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_547),
.B(n_361),
.Y(n_578)
);

NAND2x1p5_ASAP7_75t_L g579 ( 
.A(n_523),
.B(n_480),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_550),
.B(n_480),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_567),
.A2(n_530),
.B1(n_543),
.B2(n_517),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_582),
.A2(n_590),
.B1(n_594),
.B2(n_572),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_581),
.B(n_515),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_585),
.B(n_589),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_587),
.A2(n_600),
.B1(n_493),
.B2(n_522),
.Y(n_620)
);

O2A1O1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_588),
.A2(n_596),
.B(n_565),
.C(n_577),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_581),
.B(n_524),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_575),
.B(n_519),
.C(n_520),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_597),
.B(n_598),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_573),
.B(n_519),
.C(n_520),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_562),
.B(n_517),
.C(n_516),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_599),
.B(n_605),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_576),
.A2(n_547),
.B1(n_541),
.B2(n_549),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_580),
.B(n_539),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_601),
.B(n_602),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_554),
.B(n_539),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g604 ( 
.A1(n_556),
.A2(n_541),
.B(n_534),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_604),
.B(n_568),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_579),
.B(n_551),
.C(n_564),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_559),
.B(n_529),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_606),
.B(n_563),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_606),
.B(n_555),
.Y(n_608)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_608),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_587),
.A2(n_579),
.B(n_572),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_610),
.A2(n_623),
.B(n_601),
.Y(n_635)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_611),
.Y(n_633)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_612),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_582),
.A2(n_565),
.B1(n_552),
.B2(n_563),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_613),
.A2(n_622),
.B1(n_624),
.B2(n_625),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_614),
.B(n_619),
.Y(n_628)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_595),
.Y(n_615)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_615),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_616),
.B(n_618),
.Y(n_639)
);

AOI322xp5_ASAP7_75t_L g617 ( 
.A1(n_586),
.A2(n_553),
.A3(n_569),
.B1(n_560),
.B2(n_529),
.C1(n_521),
.C2(n_534),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_617),
.B(n_603),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_592),
.B(n_521),
.C(n_570),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_SL g619 ( 
.A(n_584),
.B(n_522),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_620),
.B(n_598),
.Y(n_636)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_600),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_621),
.B(n_597),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_591),
.A2(n_605),
.B1(n_593),
.B2(n_596),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_SL g623 ( 
.A1(n_591),
.A2(n_401),
.B(n_250),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_602),
.A2(n_438),
.B1(n_269),
.B2(n_267),
.Y(n_624)
);

AOI221xp5_ASAP7_75t_L g625 ( 
.A1(n_583),
.A2(n_438),
.B1(n_320),
.B2(n_176),
.C(n_285),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_618),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_629),
.B(n_631),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_607),
.B(n_589),
.Y(n_631)
);

INVx11_ASAP7_75t_L g634 ( 
.A(n_620),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_634),
.A2(n_623),
.B1(n_438),
.B2(n_254),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_635),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_SL g652 ( 
.A1(n_636),
.A2(n_641),
.B1(n_613),
.B2(n_619),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_609),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_637),
.B(n_638),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_607),
.B(n_585),
.Y(n_638)
);

CKINVDCx14_ASAP7_75t_R g650 ( 
.A(n_640),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_627),
.B(n_599),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_643),
.B(n_644),
.Y(n_647)
);

CKINVDCx16_ASAP7_75t_R g644 ( 
.A(n_608),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_643),
.B(n_626),
.C(n_592),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_649),
.B(n_654),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_642),
.A2(n_622),
.B(n_614),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_651),
.A2(n_636),
.B(n_632),
.Y(n_665)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_652),
.Y(n_660)
);

XOR2xp5_ASAP7_75t_L g653 ( 
.A(n_631),
.B(n_627),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_653),
.B(n_638),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_639),
.B(n_611),
.C(n_610),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_636),
.B(n_584),
.C(n_624),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_655),
.B(n_656),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_SL g657 ( 
.A(n_645),
.B(n_288),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_657),
.B(n_234),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_661),
.B(n_662),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_649),
.B(n_646),
.C(n_654),
.Y(n_662)
);

XOR2xp5_ASAP7_75t_L g673 ( 
.A(n_663),
.B(n_628),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_665),
.A2(n_667),
.B1(n_658),
.B2(n_650),
.Y(n_668)
);

NAND2xp67_ASAP7_75t_SL g666 ( 
.A(n_658),
.B(n_633),
.Y(n_666)
);

XNOR2xp5_ASAP7_75t_SL g670 ( 
.A(n_666),
.B(n_628),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_648),
.B(n_630),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_668),
.A2(n_669),
.B(n_664),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_662),
.B(n_647),
.C(n_653),
.Y(n_669)
);

AO21x1_ASAP7_75t_SL g676 ( 
.A1(n_670),
.A2(n_666),
.B(n_634),
.Y(n_676)
);

XOR2xp5_ASAP7_75t_L g671 ( 
.A(n_659),
.B(n_655),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_671),
.B(n_673),
.C(n_660),
.Y(n_675)
);

XOR2xp5_ASAP7_75t_L g677 ( 
.A(n_674),
.B(n_675),
.Y(n_677)
);

AOI322xp5_ASAP7_75t_L g678 ( 
.A1(n_676),
.A2(n_670),
.A3(n_672),
.B1(n_671),
.B2(n_176),
.C1(n_254),
.C2(n_279),
.Y(n_678)
);

OAI311xp33_ASAP7_75t_L g679 ( 
.A1(n_678),
.A2(n_293),
.A3(n_158),
.B1(n_159),
.C1(n_205),
.Y(n_679)
);

OAI21xp33_ASAP7_75t_L g680 ( 
.A1(n_679),
.A2(n_677),
.B(n_227),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g681 ( 
.A(n_680),
.B(n_178),
.C(n_12),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_681),
.A2(n_12),
.B1(n_13),
.B2(n_440),
.Y(n_682)
);

XNOR2xp5_ASAP7_75t_L g683 ( 
.A(n_682),
.B(n_13),
.Y(n_683)
);


endmodule