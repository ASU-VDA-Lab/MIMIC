module fake_ariane_1247_n_834 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_834);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_834;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_259;
wire n_808;
wire n_553;
wire n_446;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_569;
wire n_247;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_604;
wire n_439;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_571;
wire n_414;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_804;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_626;
wire n_430;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_517;
wire n_246;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_650;
wire n_258;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx2_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_22),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_93),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_135),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_102),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_55),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_22),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_51),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_20),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_89),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_85),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_118),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_142),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_108),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_119),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_14),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_54),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_57),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_3),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_109),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_13),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_7),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_33),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_8),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_132),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_11),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_67),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_129),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_3),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_151),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_1),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_120),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_92),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_16),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_80),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_1),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_117),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_158),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_148),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_144),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_79),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_84),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_116),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_160),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_136),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_103),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_88),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_0),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_172),
.B(n_173),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_176),
.B(n_0),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_181),
.B(n_185),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_186),
.B(n_187),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_2),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_193),
.B(n_4),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_175),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_4),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_5),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_207),
.B(n_5),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_171),
.B(n_30),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_171),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_184),
.B(n_6),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_220),
.B(n_6),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_205),
.B(n_7),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_184),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g269 ( 
.A(n_177),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_208),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_221),
.B(n_222),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_204),
.B(n_8),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_227),
.B(n_9),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_9),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_174),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_10),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_204),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_182),
.B(n_10),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_180),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_178),
.B(n_11),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_188),
.B(n_12),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g285 ( 
.A(n_210),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_240),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_211),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_240),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_201),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_179),
.Y(n_291)
);

OR2x6_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_269),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

AO22x2_ASAP7_75t_L g294 ( 
.A1(n_264),
.A2(n_219),
.B1(n_229),
.B2(n_224),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_251),
.A2(n_216),
.B1(n_218),
.B2(n_225),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_179),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_183),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

AO22x2_ASAP7_75t_L g299 ( 
.A1(n_264),
.A2(n_237),
.B1(n_194),
.B2(n_189),
.Y(n_299)
);

AO22x2_ASAP7_75t_L g300 ( 
.A1(n_264),
.A2(n_237),
.B1(n_194),
.B2(n_189),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_269),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_272),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_241),
.B(n_190),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_248),
.A2(n_235),
.B1(n_234),
.B2(n_233),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_241),
.B(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

OA22x2_ASAP7_75t_L g309 ( 
.A1(n_252),
.A2(n_232),
.B1(n_230),
.B2(n_228),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_191),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_277),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

OA22x2_ASAP7_75t_L g313 ( 
.A1(n_252),
.A2(n_226),
.B1(n_217),
.B2(n_215),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_192),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_254),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_L g316 ( 
.A1(n_285),
.A2(n_206),
.B1(n_203),
.B2(n_200),
.Y(n_316)
);

OA22x2_ASAP7_75t_L g317 ( 
.A1(n_270),
.A2(n_198),
.B1(n_195),
.B2(n_14),
.Y(n_317)
);

OR2x6_ASAP7_75t_L g318 ( 
.A(n_272),
.B(n_12),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_L g319 ( 
.A1(n_271),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_L g320 ( 
.A1(n_243),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_L g321 ( 
.A1(n_253),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_270),
.B(n_19),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_284),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_257),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_273),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_273),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_256),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_L g328 ( 
.A1(n_266),
.A2(n_275),
.B1(n_250),
.B2(n_239),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_264),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_249),
.Y(n_330)
);

AO22x2_ASAP7_75t_L g331 ( 
.A1(n_239),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_260),
.B(n_265),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_260),
.B(n_36),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_L g334 ( 
.A1(n_239),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_265),
.B(n_40),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_L g336 ( 
.A1(n_239),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_250),
.B(n_274),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_332),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_286),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_267),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_296),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_263),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_330),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_289),
.B(n_267),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

XOR2x2_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_281),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_307),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_290),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_263),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_314),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_293),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_302),
.B(n_250),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_303),
.B(n_250),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_263),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_287),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_335),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

NAND2xp33_ASAP7_75t_SL g374 ( 
.A(n_331),
.B(n_276),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_317),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_293),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_309),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_313),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_292),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_328),
.Y(n_380)
);

BUFx5_ASAP7_75t_L g381 ( 
.A(n_331),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_329),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_327),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_294),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_292),
.B(n_279),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_325),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_334),
.B(n_263),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_294),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_299),
.B(n_44),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_300),
.B(n_318),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_305),
.B(n_295),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_300),
.B(n_45),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_316),
.B(n_46),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_318),
.Y(n_396)
);

NAND2x1p5_ASAP7_75t_L g397 ( 
.A(n_336),
.B(n_268),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_324),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_319),
.B(n_47),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_320),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_321),
.B(n_263),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_306),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_289),
.B(n_259),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_298),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_364),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_342),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_349),
.B(n_263),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_268),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_370),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_350),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_387),
.A2(n_259),
.B(n_278),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_367),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_368),
.A2(n_259),
.B(n_282),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_355),
.B(n_268),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_368),
.A2(n_259),
.B(n_282),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_259),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_354),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_344),
.B(n_268),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_361),
.B(n_268),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_362),
.B(n_268),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_340),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_346),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_354),
.B(n_278),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_404),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_404),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_380),
.B(n_259),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_371),
.B(n_259),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_278),
.Y(n_432)
);

INVx8_ASAP7_75t_L g433 ( 
.A(n_370),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_351),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_356),
.B(n_278),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_372),
.B(n_278),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_48),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_370),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_357),
.Y(n_441)
);

INVx3_ASAP7_75t_SL g442 ( 
.A(n_379),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_358),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_363),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_397),
.Y(n_445)
);

NAND2x1p5_ASAP7_75t_L g446 ( 
.A(n_387),
.B(n_244),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_359),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_356),
.B(n_278),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

AND2x2_ASAP7_75t_SL g450 ( 
.A(n_381),
.B(n_238),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_365),
.B(n_238),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_338),
.B(n_238),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_341),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_343),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_386),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_381),
.B(n_401),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_345),
.B(n_282),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_402),
.Y(n_461)
);

BUFx4f_ASAP7_75t_L g462 ( 
.A(n_397),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_339),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_373),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_382),
.B(n_49),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_381),
.B(n_282),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_381),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_375),
.B(n_238),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_401),
.B(n_282),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_400),
.B(n_245),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_381),
.B(n_282),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_403),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_377),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_378),
.B(n_245),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_383),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_394),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_413),
.B(n_352),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_391),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_392),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_406),
.B(n_415),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_420),
.B(n_352),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_392),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_407),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_458),
.B(n_384),
.Y(n_485)
);

OR2x6_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_390),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_457),
.B(n_388),
.Y(n_487)
);

CKINVDCx11_ASAP7_75t_R g488 ( 
.A(n_442),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_420),
.B(n_366),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_433),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_433),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_433),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_442),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_433),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_457),
.B(n_379),
.Y(n_495)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_374),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_456),
.B(n_396),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_433),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_407),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_458),
.B(n_374),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_445),
.B(n_396),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_459),
.B(n_347),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_458),
.B(n_348),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_437),
.B(n_348),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_475),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_421),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_465),
.B(n_366),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_437),
.B(n_399),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_425),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_437),
.B(n_395),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_451),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_425),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_412),
.Y(n_518)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_405),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_442),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_462),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_434),
.Y(n_522)
);

NOR2x1_ASAP7_75t_L g523 ( 
.A(n_449),
.B(n_389),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_424),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_441),
.B(n_393),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_408),
.B(n_347),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_450),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_441),
.B(n_245),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_462),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_464),
.B(n_245),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_464),
.B(n_245),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_450),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_514),
.Y(n_533)
);

BUFx4f_ASAP7_75t_SL g534 ( 
.A(n_493),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_494),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_490),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_490),
.Y(n_537)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_490),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_502),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_488),
.Y(n_540)
);

NAND2x1p5_ASAP7_75t_L g541 ( 
.A(n_505),
.B(n_468),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_526),
.Y(n_542)
);

BUFx2_ASAP7_75t_R g543 ( 
.A(n_478),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_517),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_493),
.Y(n_545)
);

INVx5_ASAP7_75t_SL g546 ( 
.A(n_495),
.Y(n_546)
);

BUFx12f_ASAP7_75t_L g547 ( 
.A(n_488),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_505),
.Y(n_548)
);

NAND2x1p5_ASAP7_75t_L g549 ( 
.A(n_505),
.B(n_468),
.Y(n_549)
);

INVx6_ASAP7_75t_L g550 ( 
.A(n_490),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_495),
.B(n_466),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_524),
.Y(n_552)
);

INVx3_ASAP7_75t_SL g553 ( 
.A(n_520),
.Y(n_553)
);

CKINVDCx8_ASAP7_75t_R g554 ( 
.A(n_526),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_522),
.Y(n_555)
);

NAND2x1p5_ASAP7_75t_L g556 ( 
.A(n_505),
.B(n_449),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_518),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_501),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_518),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_491),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_494),
.Y(n_561)
);

BUFx4f_ASAP7_75t_L g562 ( 
.A(n_496),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_476),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g564 ( 
.A(n_501),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_492),
.Y(n_565)
);

BUFx8_ASAP7_75t_L g566 ( 
.A(n_516),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g567 ( 
.A1(n_515),
.A2(n_466),
.B1(n_450),
.B2(n_461),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_482),
.B(n_461),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_502),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_501),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_491),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_508),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_513),
.B(n_434),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_509),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_525),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_524),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_497),
.Y(n_577)
);

BUFx4_ASAP7_75t_SL g578 ( 
.A(n_492),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_491),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_513),
.B(n_440),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_497),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_551),
.A2(n_515),
.B1(n_481),
.B2(n_476),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_572),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_551),
.A2(n_481),
.B1(n_476),
.B2(n_506),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_574),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_547),
.Y(n_586)
);

INVxp67_ASAP7_75t_SL g587 ( 
.A(n_557),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_567),
.A2(n_476),
.B1(n_523),
.B2(n_525),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_573),
.A2(n_510),
.B1(n_580),
.B2(n_449),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_568),
.A2(n_476),
.B1(n_506),
.B2(n_466),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_575),
.A2(n_506),
.B1(n_466),
.B2(n_480),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_566),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_575),
.A2(n_506),
.B1(n_480),
.B2(n_483),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_L g594 ( 
.A1(n_554),
.A2(n_500),
.B1(n_510),
.B2(n_504),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_533),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_553),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_544),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_SL g598 ( 
.A1(n_539),
.A2(n_506),
.B1(n_500),
.B2(n_483),
.Y(n_598)
);

INVx6_ASAP7_75t_L g599 ( 
.A(n_566),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_548),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_566),
.Y(n_601)
);

OAI21xp33_ASAP7_75t_L g602 ( 
.A1(n_555),
.A2(n_443),
.B(n_440),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_552),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_552),
.Y(n_604)
);

INVx6_ASAP7_75t_L g605 ( 
.A(n_547),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_551),
.A2(n_443),
.B1(n_447),
.B2(n_504),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_557),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_576),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_546),
.A2(n_447),
.B1(n_532),
.B2(n_527),
.Y(n_609)
);

CKINVDCx14_ASAP7_75t_R g610 ( 
.A(n_540),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_SL g611 ( 
.A1(n_563),
.A2(n_479),
.B1(n_477),
.B2(n_487),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_577),
.A2(n_512),
.B1(n_477),
.B2(n_479),
.Y(n_612)
);

OAI22xp33_ASAP7_75t_L g613 ( 
.A1(n_553),
.A2(n_496),
.B1(n_532),
.B2(n_527),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_569),
.A2(n_487),
.B1(n_529),
.B2(n_521),
.Y(n_614)
);

INVx11_ASAP7_75t_L g615 ( 
.A(n_564),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_L g616 ( 
.A1(n_542),
.A2(n_485),
.B1(n_486),
.B2(n_454),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_581),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_576),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_558),
.A2(n_534),
.B1(n_545),
.B2(n_562),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_545),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_534),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_546),
.A2(n_562),
.B1(n_563),
.B2(n_556),
.Y(n_622)
);

OAI22xp33_ASAP7_75t_L g623 ( 
.A1(n_558),
.A2(n_485),
.B1(n_486),
.B2(n_454),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_564),
.A2(n_489),
.B1(n_486),
.B2(n_421),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_559),
.Y(n_625)
);

BUFx4_ASAP7_75t_R g626 ( 
.A(n_559),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_570),
.A2(n_426),
.B1(n_509),
.B2(n_503),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_590),
.A2(n_570),
.B1(n_435),
.B2(n_448),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_606),
.A2(n_563),
.B1(n_543),
.B2(n_546),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_591),
.A2(n_563),
.B1(n_428),
.B2(n_429),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_588),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_596),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_594),
.A2(n_427),
.B1(n_424),
.B2(n_499),
.Y(n_633)
);

OAI22xp33_ASAP7_75t_L g634 ( 
.A1(n_582),
.A2(n_548),
.B1(n_556),
.B2(n_540),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_589),
.A2(n_484),
.B1(n_455),
.B2(n_507),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_623),
.A2(n_455),
.B1(n_473),
.B2(n_423),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_584),
.A2(n_561),
.B1(n_535),
.B2(n_565),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_583),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_587),
.Y(n_639)
);

BUFx8_ASAP7_75t_SL g640 ( 
.A(n_621),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_606),
.A2(n_549),
.B(n_541),
.Y(n_641)
);

OAI21xp33_ASAP7_75t_SL g642 ( 
.A1(n_627),
.A2(n_548),
.B(n_535),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_616),
.A2(n_455),
.B1(n_422),
.B2(n_531),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_612),
.A2(n_455),
.B1(n_530),
.B2(n_452),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_607),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_596),
.B(n_620),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_619),
.A2(n_578),
.B(n_561),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_595),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_597),
.B(n_585),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_626),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_603),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_613),
.B(n_536),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_598),
.A2(n_455),
.B1(n_452),
.B2(n_453),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_593),
.A2(n_453),
.B1(n_471),
.B2(n_419),
.Y(n_654)
);

AND2x4_ASAP7_75t_SL g655 ( 
.A(n_607),
.B(n_537),
.Y(n_655)
);

AOI211xp5_ASAP7_75t_L g656 ( 
.A1(n_592),
.A2(n_602),
.B(n_625),
.C(n_601),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_599),
.A2(n_565),
.B1(n_446),
.B2(n_538),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_599),
.A2(n_446),
.B1(n_538),
.B2(n_550),
.Y(n_658)
);

INVx6_ASAP7_75t_L g659 ( 
.A(n_607),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_605),
.A2(n_549),
.B1(n_541),
.B2(n_446),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_604),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_624),
.A2(n_471),
.B1(n_419),
.B2(n_474),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_608),
.Y(n_663)
);

INVx5_ASAP7_75t_SL g664 ( 
.A(n_615),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_614),
.A2(n_550),
.B1(n_538),
.B2(n_503),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_605),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_586),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_617),
.A2(n_550),
.B1(n_519),
.B2(n_571),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_610),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_609),
.A2(n_419),
.B1(n_474),
.B2(n_431),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_611),
.A2(n_519),
.B1(n_571),
.B2(n_560),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_618),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_609),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_600),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_622),
.A2(n_414),
.B1(n_470),
.B2(n_430),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_622),
.A2(n_414),
.B1(n_430),
.B2(n_416),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_SL g677 ( 
.A1(n_600),
.A2(n_418),
.B1(n_419),
.B2(n_431),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_629),
.A2(n_460),
.B1(n_432),
.B2(n_436),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_672),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_SL g680 ( 
.A1(n_647),
.A2(n_578),
.B(n_410),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_639),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_648),
.Y(n_682)
);

AOI222xp33_ASAP7_75t_L g683 ( 
.A1(n_673),
.A2(n_469),
.B1(n_528),
.B2(n_444),
.C1(n_439),
.C2(n_463),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_649),
.Y(n_684)
);

AOI221xp5_ASAP7_75t_L g685 ( 
.A1(n_632),
.A2(n_469),
.B1(n_528),
.B2(n_463),
.C(n_439),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_631),
.A2(n_662),
.B1(n_638),
.B2(n_670),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_650),
.A2(n_579),
.B1(n_560),
.B2(n_536),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_631),
.A2(n_460),
.B1(n_463),
.B2(n_444),
.Y(n_688)
);

OA21x2_ASAP7_75t_L g689 ( 
.A1(n_635),
.A2(n_411),
.B(n_417),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_646),
.B(n_579),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_628),
.A2(n_444),
.B1(n_439),
.B2(n_467),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_651),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_657),
.A2(n_536),
.B1(n_560),
.B2(n_519),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_636),
.A2(n_643),
.B1(n_654),
.B2(n_644),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_SL g695 ( 
.A1(n_634),
.A2(n_536),
.B(n_498),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_656),
.A2(n_511),
.B1(n_498),
.B2(n_491),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_661),
.Y(n_697)
);

AO22x1_ASAP7_75t_L g698 ( 
.A1(n_637),
.A2(n_658),
.B1(n_645),
.B2(n_666),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_663),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_635),
.A2(n_630),
.B1(n_653),
.B2(n_634),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_645),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_652),
.A2(n_472),
.B1(n_438),
.B2(n_412),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_630),
.A2(n_633),
.B1(n_675),
.B2(n_677),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_660),
.A2(n_438),
.B1(n_511),
.B2(n_537),
.Y(n_704)
);

INVxp67_ASAP7_75t_SL g705 ( 
.A(n_674),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_633),
.A2(n_438),
.B1(n_511),
.B2(n_405),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_675),
.A2(n_511),
.B1(n_405),
.B2(n_537),
.Y(n_707)
);

AOI222xp33_ASAP7_75t_L g708 ( 
.A1(n_642),
.A2(n_676),
.B1(n_660),
.B2(n_665),
.C1(n_668),
.C2(n_671),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_676),
.A2(n_405),
.B1(n_247),
.B2(n_246),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_641),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_659),
.A2(n_247),
.B1(n_246),
.B2(n_258),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_659),
.A2(n_247),
.B1(n_246),
.B2(n_258),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_645),
.B(n_246),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_SL g714 ( 
.A1(n_659),
.A2(n_247),
.B1(n_246),
.B2(n_255),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_645),
.A2(n_247),
.B1(n_255),
.B2(n_258),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_667),
.A2(n_258),
.B1(n_255),
.B2(n_244),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_655),
.B(n_50),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_667),
.A2(n_258),
.B1(n_255),
.B2(n_244),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g719 ( 
.A(n_681),
.B(n_710),
.C(n_708),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_682),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_705),
.B(n_669),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_703),
.A2(n_664),
.B1(n_640),
.B2(n_258),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_682),
.B(n_664),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_684),
.B(n_664),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_679),
.B(n_52),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_679),
.B(n_53),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_690),
.B(n_56),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_701),
.B(n_58),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_692),
.B(n_59),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_710),
.B(n_255),
.C(n_244),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_L g731 ( 
.A(n_700),
.B(n_255),
.C(n_244),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_692),
.B(n_60),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_680),
.B(n_695),
.C(n_696),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_698),
.B(n_61),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_697),
.B(n_62),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_697),
.B(n_63),
.Y(n_736)
);

OAI221xp5_ASAP7_75t_L g737 ( 
.A1(n_694),
.A2(n_244),
.B1(n_65),
.B2(n_66),
.C(n_68),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_689),
.B(n_64),
.C(n_70),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_699),
.B(n_689),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_SL g740 ( 
.A1(n_707),
.A2(n_72),
.B(n_73),
.Y(n_740)
);

OA21x2_ASAP7_75t_L g741 ( 
.A1(n_713),
.A2(n_74),
.B(n_75),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_699),
.B(n_169),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_689),
.B(n_76),
.Y(n_743)
);

NAND3xp33_ASAP7_75t_L g744 ( 
.A(n_683),
.B(n_77),
.C(n_78),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_698),
.B(n_168),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_687),
.B(n_686),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_704),
.B(n_81),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_693),
.B(n_167),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_720),
.Y(n_749)
);

NOR2x1_ASAP7_75t_L g750 ( 
.A(n_719),
.B(n_717),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_740),
.B(n_685),
.C(n_714),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_L g752 ( 
.A(n_744),
.B(n_737),
.C(n_722),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_739),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_733),
.B(n_709),
.C(n_691),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_723),
.Y(n_755)
);

NOR2x1_ASAP7_75t_L g756 ( 
.A(n_724),
.B(n_721),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_733),
.A2(n_678),
.B1(n_702),
.B2(n_706),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_L g758 ( 
.A(n_738),
.B(n_688),
.C(n_716),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_739),
.B(n_718),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_743),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_746),
.B(n_712),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_731),
.B(n_711),
.C(n_715),
.Y(n_762)
);

NAND4xp75_ASAP7_75t_L g763 ( 
.A(n_734),
.B(n_82),
.C(n_83),
.D(n_86),
.Y(n_763)
);

XOR2x2_ASAP7_75t_L g764 ( 
.A(n_734),
.B(n_87),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_725),
.Y(n_765)
);

NAND4xp75_ASAP7_75t_L g766 ( 
.A(n_745),
.B(n_90),
.C(n_91),
.D(n_94),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_755),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_755),
.B(n_743),
.Y(n_768)
);

NAND4xp75_ASAP7_75t_L g769 ( 
.A(n_750),
.B(n_727),
.C(n_748),
.D(n_741),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_765),
.B(n_726),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_749),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_753),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_752),
.B(n_747),
.C(n_735),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_756),
.B(n_728),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_764),
.Y(n_775)
);

NAND4xp75_ASAP7_75t_SL g776 ( 
.A(n_759),
.B(n_741),
.C(n_730),
.D(n_736),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_760),
.B(n_732),
.Y(n_777)
);

NAND4xp75_ASAP7_75t_L g778 ( 
.A(n_757),
.B(n_741),
.C(n_729),
.D(n_742),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_774),
.Y(n_779)
);

OA22x2_ASAP7_75t_L g780 ( 
.A1(n_775),
.A2(n_754),
.B1(n_751),
.B2(n_763),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_771),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_772),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_770),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_777),
.Y(n_784)
);

XOR2x2_ASAP7_75t_L g785 ( 
.A(n_780),
.B(n_769),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_779),
.A2(n_778),
.B1(n_767),
.B2(n_773),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_783),
.B(n_784),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_782),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_788),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_787),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_785),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_786),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_789),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_790),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_791),
.A2(n_780),
.B1(n_773),
.B2(n_754),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_793),
.A2(n_792),
.B(n_761),
.C(n_758),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_794),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_795),
.A2(n_792),
.B1(n_767),
.B2(n_768),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_795),
.A2(n_758),
.B(n_781),
.C(n_776),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_799),
.A2(n_766),
.B1(n_776),
.B2(n_762),
.Y(n_800)
);

NOR4xp25_ASAP7_75t_L g801 ( 
.A(n_796),
.B(n_762),
.C(n_96),
.D(n_97),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_797),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_798),
.A2(n_95),
.B1(n_99),
.B2(n_101),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_797),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_802),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_804),
.B(n_104),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_800),
.A2(n_105),
.B1(n_107),
.B2(n_110),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_803),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_801),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_800),
.A2(n_115),
.B1(n_121),
.B2(n_123),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_805),
.Y(n_811)
);

AND4x1_ASAP7_75t_L g812 ( 
.A(n_806),
.B(n_125),
.C(n_126),
.D(n_127),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_808),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_810),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_811),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_813),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_814),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_812),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_811),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_816),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_817),
.Y(n_821)
);

OAI22x1_ASAP7_75t_L g822 ( 
.A1(n_816),
.A2(n_807),
.B1(n_809),
.B2(n_133),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_815),
.A2(n_128),
.B1(n_130),
.B2(n_137),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_820),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_821),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_822),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_826),
.A2(n_818),
.B1(n_819),
.B2(n_823),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_825),
.A2(n_166),
.B1(n_146),
.B2(n_149),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_824),
.A2(n_145),
.B1(n_150),
.B2(n_153),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_827),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_830),
.A2(n_824),
.B1(n_828),
.B2(n_829),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_831),
.B(n_154),
.Y(n_832)
);

AOI221xp5_ASAP7_75t_L g833 ( 
.A1(n_832),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.C(n_159),
.Y(n_833)
);

AOI211xp5_ASAP7_75t_L g834 ( 
.A1(n_833),
.A2(n_161),
.B(n_162),
.C(n_164),
.Y(n_834)
);


endmodule