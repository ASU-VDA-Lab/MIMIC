module real_jpeg_6976_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_L g233 ( 
.A(n_0),
.B(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_0),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_0),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_0),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_0),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_0),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_0),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_0),
.B(n_373),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_1),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_1),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_1),
.B(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_1),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_1),
.B(n_216),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_1),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_1),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_2),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_2),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_2),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_2),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_2),
.B(n_34),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_2),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_3),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_3),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_3),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_3),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_190),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_3),
.B(n_288),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_3),
.B(n_421),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_4),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_4),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_4),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_4),
.B(n_437),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_5),
.Y(n_98)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_5),
.Y(n_192)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_5),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_5),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_5),
.Y(n_318)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_6),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_6),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_6),
.Y(n_169)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_6),
.Y(n_209)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_6),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_7),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_8),
.B(n_161),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_8),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_8),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_8),
.B(n_190),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_8),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_8),
.B(n_282),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_8),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_8),
.B(n_169),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_9),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_9),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_9),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_9),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_9),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g377 ( 
.A(n_9),
.B(n_286),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_9),
.B(n_446),
.Y(n_445)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_11),
.Y(n_518)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_12),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_12),
.Y(n_282)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_14),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_14),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_14),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_14),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_14),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_14),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_14),
.B(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_15),
.Y(n_448)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_17),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_17),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_17),
.B(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_17),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_17),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_17),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_17),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_17),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_18),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_18),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_18),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_18),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_18),
.B(n_305),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_18),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_18),
.B(n_373),
.Y(n_372)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_517),
.B(n_519),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_171),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_170),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_149),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_24),
.B(n_149),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_111),
.C(n_122),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_25),
.B(n_502),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_79),
.C(n_93),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_26),
.B(n_505),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_47),
.C(n_60),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_27),
.B(n_47),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_28),
.B(n_38),
.C(n_46),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_29),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_29),
.B(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_31),
.Y(n_266)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_31),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_38),
.B1(n_39),
.B2(n_46),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_36),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_36),
.Y(n_439)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_37),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_37),
.Y(n_249)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_37),
.Y(n_338)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_43),
.Y(n_390)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_44),
.Y(n_310)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_45),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_45),
.Y(n_237)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_45),
.Y(n_245)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_45),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.C(n_57),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_48),
.B(n_57),
.Y(n_466)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_52),
.B(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_55),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_56),
.Y(n_217)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_60),
.B(n_494),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_61),
.B(n_69),
.C(n_78),
.Y(n_120)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_67),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_78),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_70),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_114),
.C(n_117),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_96),
.C(n_99),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_73),
.A2(n_78),
.B1(n_96),
.B2(n_97),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_76),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_77),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_77),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_79),
.A2(n_93),
.B1(n_94),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_79),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_84),
.C(n_88),
.Y(n_138)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_86),
.Y(n_262)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.C(n_106),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_95),
.B(n_492),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_96),
.A2(n_97),
.B1(n_445),
.B2(n_449),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_96),
.B(n_445),
.C(n_450),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_99),
.B(n_462),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_102),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_492)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_106),
.A2(n_107),
.B1(n_475),
.B2(n_476),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_107),
.B(n_476),
.C(n_490),
.Y(n_489)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_111),
.B(n_122),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_120),
.C(n_121),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_112),
.B(n_508),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_115),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_132),
.C(n_134),
.Y(n_167)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_120),
.B(n_121),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_137),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_135),
.B2(n_136),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_136),
.C(n_137),
.Y(n_150)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_130),
.B1(n_131),
.B2(n_134),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_132),
.A2(n_133),
.B1(n_160),
.B2(n_164),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_143),
.C(n_148),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_143),
.B1(n_144),
.B2(n_148),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_165),
.B2(n_166),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_160),
.Y(n_164)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g242 ( 
.A(n_163),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_163),
.Y(n_404)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

AO21x1_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_497),
.B(n_514),
.Y(n_171)
);

OAI21x1_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_481),
.B(n_496),
.Y(n_172)
);

AOI21x1_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_455),
.B(n_480),
.Y(n_173)
);

OAI21x1_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_408),
.B(n_454),
.Y(n_174)
);

AOI21x1_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_365),
.B(n_407),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_291),
.B(n_364),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_275),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_178),
.B(n_275),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_220),
.B2(n_274),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_179),
.B(n_221),
.C(n_258),
.Y(n_406)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_199),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_181),
.B(n_200),
.C(n_219),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_193),
.C(n_197),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_182),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_188),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_183),
.A2(n_184),
.B1(n_188),
.B2(n_189),
.Y(n_280)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_185),
.Y(n_299)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_187),
.Y(n_288)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_192),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_193),
.B(n_197),
.Y(n_290)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_204),
.B1(n_218),
.B2(n_219),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B(n_203),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_203),
.B(n_381),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_203),
.B(n_370),
.C(n_381),
.Y(n_415)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_205),
.B(n_211),
.C(n_215),
.Y(n_405)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx8_ASAP7_75t_L g401 ( 
.A(n_217),
.Y(n_401)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_258),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_238),
.C(n_250),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_233),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_224),
.B(n_228),
.C(n_233),
.Y(n_273)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_238),
.A2(n_239),
.B1(n_250),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.C(n_246),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_240),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_357)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_243),
.B(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_255),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_255),
.Y(n_272)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2x1_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_271),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_259),
.B(n_272),
.C(n_273),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g381 ( 
.A(n_260),
.B(n_267),
.C(n_269),
.Y(n_381)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_267),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.C(n_289),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_276),
.B(n_362),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_279),
.B(n_289),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.C(n_283),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_280),
.B(n_281),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_283),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_287),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_359),
.B(n_363),
.Y(n_291)
);

OA21x2_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_344),
.B(n_358),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_328),
.B(n_343),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_319),
.B(n_327),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_301),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_301),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_300),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_311),
.B2(n_312),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_307),
.C(n_311),
.Y(n_342)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_335),
.Y(n_334)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_317),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_317),
.Y(n_332)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_323),
.B(n_326),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_322),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_342),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_342),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_332),
.C(n_346),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_336),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_339),
.C(n_341),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_336)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_337),
.Y(n_341)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_347),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_351),
.B2(n_352),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_348),
.B(n_354),
.C(n_355),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_360),
.B(n_361),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_406),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_366),
.B(n_406),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_383),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_368),
.B(n_369),
.C(n_383),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_371),
.B1(n_380),
.B2(n_382),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_375),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_372),
.B(n_377),
.C(n_378),
.Y(n_425)
);

INVx8_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_380),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_386),
.C(n_398),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_398),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_391),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_387),
.B(n_392),
.C(n_395),
.Y(n_441)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx6_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_405),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_402),
.C(n_405),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_409),
.B(n_410),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_411),
.B(n_427),
.C(n_452),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_413),
.A2(n_427),
.B1(n_452),
.B2(n_453),
.Y(n_412)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_413),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_416),
.B2(n_426),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_417),
.C(n_418),
.Y(n_457)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_416),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_425),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_422),
.C(n_425),
.Y(n_472)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_427),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_440),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_428),
.B(n_441),
.C(n_442),
.Y(n_470)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_428),
.Y(n_523)
);

FAx1_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_433),
.CI(n_436),
.CON(n_428),
.SN(n_428)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_429),
.B(n_433),
.C(n_436),
.Y(n_477)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_443),
.A2(n_444),
.B1(n_450),
.B2(n_451),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_445),
.Y(n_449)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_479),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_479),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_457),
.B(n_459),
.C(n_468),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_468),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_461),
.B1(n_463),
.B2(n_467),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_464),
.C(n_465),
.Y(n_486)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_463),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_470),
.B1(n_471),
.B2(n_478),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_472),
.C(n_473),
.Y(n_483)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_471),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_477),
.Y(n_473)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_475),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_477),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_495),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_495),
.Y(n_496)
);

BUFx24_ASAP7_75t_SL g524 ( 
.A(n_482),
.Y(n_524)
);

FAx1_ASAP7_75t_SL g482 ( 
.A(n_483),
.B(n_484),
.CI(n_493),
.CON(n_482),
.SN(n_482)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_483),
.B(n_484),
.C(n_493),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_489),
.C(n_491),
.Y(n_509)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_491),
.Y(n_488)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_510),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_500),
.A2(n_515),
.B(n_516),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_503),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_501),
.B(n_503),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_507),
.C(n_509),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_507),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_509),
.B(n_512),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_513),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_513),
.Y(n_515)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx13_ASAP7_75t_L g521 ( 
.A(n_518),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_522),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);


endmodule