module fake_netlist_5_585_n_2920 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_551, n_17, n_382, n_554, n_254, n_33, n_23, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2920);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_551;
input n_17;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2920;

wire n_924;
wire n_1263;
wire n_1378;
wire n_977;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_2899;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_1695;
wire n_688;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_854;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_2244;
wire n_933;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_2031;
wire n_2076;
wire n_1728;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_2127;
wire n_1818;
wire n_1576;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2249;
wire n_926;
wire n_2180;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_1547;
wire n_777;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_1473;
wire n_1587;
wire n_680;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_2118;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_1447;
wire n_907;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1463;
wire n_1581;
wire n_1002;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_2919;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2674;
wire n_2606;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_1276;
wire n_702;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_728;
wire n_1538;
wire n_1162;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_931;
wire n_1711;
wire n_599;
wire n_1891;
wire n_1662;
wire n_870;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_1876;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_1537;
wire n_913;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_2022;
wire n_1798;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2913;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_1539;
wire n_946;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1994;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2339;
wire n_2320;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_750;
wire n_2029;
wire n_742;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_602;
wire n_574;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_1684;
wire n_921;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_1437;
wire n_701;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_1897;
wire n_890;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_2916;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_1954;
wire n_802;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_1644;
wire n_762;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_1983;
wire n_883;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_2169;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2751;
wire n_2707;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_669;
wire n_2471;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_1848;
wire n_1928;
wire n_783;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_1401;
wire n_969;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_876;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_703;
wire n_1115;
wire n_698;
wire n_980;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_2884;
wire n_1268;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_737;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_733;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2774;
wire n_2726;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2778;
wire n_1756;
wire n_771;
wire n_2678;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_1567;
wire n_682;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2742;
wire n_2673;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_598;
wire n_685;
wire n_1367;
wire n_608;
wire n_928;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_2208;
wire n_1404;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_722;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_2918;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2505;
wire n_2438;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_1089;
wire n_2013;
wire n_927;
wire n_1990;
wire n_2689;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_185),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_554),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_536),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_565),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_316),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_521),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_491),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_511),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_375),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_404),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_287),
.Y(n_584)
);

CKINVDCx14_ASAP7_75t_R g585 ( 
.A(n_504),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_450),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_445),
.Y(n_587)
);

INVxp67_ASAP7_75t_SL g588 ( 
.A(n_215),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_43),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_528),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_541),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_533),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_485),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_29),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_36),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_49),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_18),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_415),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_463),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_342),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_255),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_191),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_530),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_327),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_266),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_510),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_232),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_547),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_434),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_83),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_100),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_22),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_61),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_503),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_140),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_307),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_522),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_90),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_567),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_500),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_497),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_501),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_523),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_212),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_418),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_213),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_5),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_275),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_268),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_175),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_516),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_75),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_142),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_570),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_185),
.Y(n_635)
);

CKINVDCx16_ASAP7_75t_R g636 ( 
.A(n_548),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_516),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_482),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_440),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_408),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_358),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_93),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_419),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_354),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_32),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_128),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_327),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_283),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_363),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_330),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_134),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_498),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_351),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_12),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_543),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_172),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_435),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_453),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_157),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_293),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_27),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_90),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_527),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_346),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_96),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_9),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_204),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_507),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_505),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_217),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_58),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_180),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_310),
.Y(n_673)
);

INVxp33_ASAP7_75t_SL g674 ( 
.A(n_429),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_1),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_482),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_495),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_449),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_107),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_513),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_345),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_473),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_434),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_18),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_266),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_509),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_82),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_397),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_469),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_341),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_459),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_487),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_116),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_471),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_526),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_549),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_221),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_497),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_564),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_517),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_335),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_355),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_47),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_474),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_77),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_226),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_92),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_143),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_518),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_219),
.Y(n_710)
);

BUFx5_ASAP7_75t_L g711 ( 
.A(n_249),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_305),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_125),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_194),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_236),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_108),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_417),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_488),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_495),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_131),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_315),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_103),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_433),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_525),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_344),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_572),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_34),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_180),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_496),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_262),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_203),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_21),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_351),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_519),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_563),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_34),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_172),
.Y(n_737)
);

BUFx5_ASAP7_75t_L g738 ( 
.A(n_390),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_11),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_399),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_350),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_215),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_358),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_57),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_12),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_177),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_242),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_535),
.Y(n_748)
);

CKINVDCx16_ASAP7_75t_R g749 ( 
.A(n_458),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_556),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_300),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_519),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_506),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_546),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_357),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_183),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_325),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_258),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_504),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_8),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_349),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_499),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_245),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_139),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_129),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_310),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_242),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_195),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_226),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_365),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_485),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_521),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_385),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_366),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_348),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_560),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_103),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_488),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_0),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_359),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_205),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_539),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_496),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_489),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_193),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_133),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_261),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_494),
.Y(n_788)
);

BUFx2_ASAP7_75t_SL g789 ( 
.A(n_544),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_178),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_538),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_303),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_346),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_44),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_386),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_220),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_57),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_196),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_69),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_380),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_532),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_512),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_552),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_335),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_87),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_159),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_198),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_367),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_26),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_28),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_289),
.Y(n_811)
);

BUFx10_ASAP7_75t_L g812 ( 
.A(n_158),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_503),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_334),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_422),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_555),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_81),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_394),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_269),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_441),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_250),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_553),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_56),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_118),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_45),
.Y(n_825)
);

BUFx2_ASAP7_75t_SL g826 ( 
.A(n_534),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_33),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_566),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_347),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_502),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_433),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_515),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_233),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_522),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_133),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_489),
.Y(n_836)
);

BUFx2_ASAP7_75t_R g837 ( 
.A(n_511),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_558),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_22),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_139),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_573),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_182),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_427),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_98),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_481),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_272),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_275),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_141),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_440),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_203),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_525),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_537),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_40),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_292),
.Y(n_854)
);

CKINVDCx14_ASAP7_75t_R g855 ( 
.A(n_99),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_404),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_540),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_415),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_58),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_461),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_321),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_267),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_437),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_480),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_399),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_234),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_229),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_285),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_45),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_514),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_365),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_542),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_268),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_557),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_403),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_28),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_493),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_499),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_95),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_451),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_420),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_119),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_280),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_237),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_431),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_453),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_462),
.Y(n_887)
);

BUFx10_ASAP7_75t_L g888 ( 
.A(n_508),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_512),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_448),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_390),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_314),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_464),
.Y(n_893)
);

CKINVDCx16_ASAP7_75t_R g894 ( 
.A(n_230),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_213),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_144),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_473),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_265),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_14),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_160),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_380),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_461),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_221),
.Y(n_903)
);

BUFx10_ASAP7_75t_L g904 ( 
.A(n_160),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_450),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_111),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_517),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_510),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_91),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_314),
.Y(n_910)
);

CKINVDCx16_ASAP7_75t_R g911 ( 
.A(n_158),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_164),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_144),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_321),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_531),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_245),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_65),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_437),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_97),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_318),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_269),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_138),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_490),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_181),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_291),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_145),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_325),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_59),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_38),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_311),
.Y(n_930)
);

CKINVDCx16_ASAP7_75t_R g931 ( 
.A(n_568),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_0),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_467),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_344),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_397),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_561),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_123),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_562),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_498),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_373),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_148),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_520),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_289),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_214),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_569),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_227),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_432),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_193),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_13),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_235),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_338),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_25),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_74),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_239),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_395),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_524),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_551),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_356),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_227),
.Y(n_959)
);

BUFx10_ASAP7_75t_L g960 ( 
.A(n_306),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_559),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_571),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_292),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_105),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_457),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_486),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_13),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_270),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_68),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_408),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_439),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_214),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_387),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_65),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_130),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_545),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_444),
.Y(n_977)
);

BUFx10_ASAP7_75t_L g978 ( 
.A(n_419),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_427),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_220),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_106),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_5),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_373),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_173),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_301),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_135),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_118),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_48),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_274),
.Y(n_989)
);

BUFx10_ASAP7_75t_L g990 ( 
.A(n_140),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_297),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_479),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_64),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_550),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_135),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_223),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_109),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_295),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_246),
.Y(n_999)
);

BUFx8_ASAP7_75t_SL g1000 ( 
.A(n_484),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_353),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_455),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_212),
.Y(n_1003)
);

BUFx10_ASAP7_75t_L g1004 ( 
.A(n_432),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_182),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_146),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_7),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_192),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_106),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_264),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_452),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_492),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_150),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_265),
.Y(n_1014)
);

INVxp67_ASAP7_75t_SL g1015 ( 
.A(n_645),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_866),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_1000),
.Y(n_1017)
);

INVxp67_ASAP7_75t_SL g1018 ( 
.A(n_645),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_711),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_711),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_711),
.Y(n_1021)
);

INVxp33_ASAP7_75t_L g1022 ( 
.A(n_769),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_711),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_575),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_577),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_711),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_735),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_711),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_711),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_711),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_636),
.Y(n_1031)
);

CKINVDCx16_ASAP7_75t_R g1032 ( 
.A(n_585),
.Y(n_1032)
);

INVxp67_ASAP7_75t_SL g1033 ( 
.A(n_645),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_711),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_590),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_591),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_636),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_738),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_592),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_738),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_866),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_738),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_931),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_619),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_634),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_931),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_738),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_880),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_663),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_575),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_738),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_738),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_880),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_738),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_596),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_696),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_738),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_738),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_855),
.Y(n_1059)
);

INVxp33_ASAP7_75t_L g1060 ( 
.A(n_877),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_581),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_581),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_581),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_645),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_579),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_581),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_581),
.Y(n_1067)
);

INVxp67_ASAP7_75t_SL g1068 ( 
.A(n_945),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_581),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_699),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_610),
.Y(n_1071)
);

INVxp67_ASAP7_75t_SL g1072 ( 
.A(n_945),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_726),
.Y(n_1073)
);

INVxp67_ASAP7_75t_L g1074 ( 
.A(n_579),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_748),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_610),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_610),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_610),
.Y(n_1078)
);

INVxp67_ASAP7_75t_SL g1079 ( 
.A(n_610),
.Y(n_1079)
);

INVxp33_ASAP7_75t_SL g1080 ( 
.A(n_574),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_583),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_791),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_610),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_639),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_874),
.Y(n_1085)
);

CKINVDCx16_ASAP7_75t_R g1086 ( 
.A(n_749),
.Y(n_1086)
);

INVxp67_ASAP7_75t_SL g1087 ( 
.A(n_639),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_639),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_803),
.Y(n_1089)
);

OA21x2_ASAP7_75t_L g1090 ( 
.A1(n_1061),
.A2(n_1063),
.B(n_1062),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1079),
.B(n_639),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1026),
.A2(n_957),
.B(n_754),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1026),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_1085),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_1025),
.Y(n_1095)
);

CKINVDCx6p67_ASAP7_75t_R g1096 ( 
.A(n_1032),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_1085),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1061),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1062),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_1087),
.B(n_603),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1088),
.B(n_603),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1029),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1029),
.Y(n_1103)
);

INVx5_ASAP7_75t_L g1104 ( 
.A(n_1085),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_1085),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1064),
.B(n_915),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1030),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1063),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_1085),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1030),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1015),
.B(n_639),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1066),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1066),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1067),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1085),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_1080),
.B(n_915),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1018),
.B(n_1033),
.Y(n_1117)
);

INVx5_ASAP7_75t_L g1118 ( 
.A(n_1064),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1068),
.B(n_639),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1067),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1069),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1069),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1072),
.B(n_657),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1071),
.B(n_657),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1071),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1055),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_SL g1127 ( 
.A1(n_1031),
.A2(n_578),
.B1(n_595),
.B2(n_582),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1076),
.B(n_1077),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_L g1129 ( 
.A(n_1076),
.B(n_789),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1019),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1019),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1077),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1032),
.B(n_749),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1078),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1078),
.B(n_657),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1020),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1083),
.B(n_657),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1083),
.B(n_657),
.Y(n_1138)
);

INVx5_ASAP7_75t_L g1139 ( 
.A(n_1024),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1084),
.B(n_657),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1084),
.B(n_957),
.Y(n_1141)
);

CKINVDCx11_ASAP7_75t_R g1142 ( 
.A(n_1059),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1020),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1021),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1021),
.B(n_750),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1023),
.B(n_750),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1024),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_1023),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1028),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1028),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1024),
.B(n_660),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1124),
.A2(n_1038),
.B(n_1034),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1116),
.B(n_1035),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1149),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1126),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1149),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1096),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_R g1158 ( 
.A(n_1095),
.B(n_1036),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1096),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1096),
.Y(n_1160)
);

BUFx10_ASAP7_75t_L g1161 ( 
.A(n_1117),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1139),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1130),
.Y(n_1163)
);

CKINVDCx16_ASAP7_75t_R g1164 ( 
.A(n_1126),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1142),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_1133),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1130),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1093),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1130),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1093),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1130),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1127),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1127),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1136),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1147),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1147),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1147),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1117),
.B(n_1039),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1136),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1117),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_1119),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1093),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1136),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1094),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_1111),
.B(n_1044),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1102),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1136),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1119),
.Y(n_1188)
);

NOR2xp67_ASAP7_75t_L g1189 ( 
.A(n_1139),
.B(n_1056),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_1123),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1145),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1148),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1117),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1145),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1145),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1148),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_1123),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1092),
.A2(n_1038),
.B(n_1034),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1145),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1111),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1145),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1151),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1148),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_1151),
.Y(n_1204)
);

CKINVDCx16_ASAP7_75t_R g1205 ( 
.A(n_1100),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1148),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1091),
.Y(n_1207)
);

INVxp67_ASAP7_75t_SL g1208 ( 
.A(n_1091),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1094),
.Y(n_1209)
);

AND2x2_ASAP7_75t_SL g1210 ( 
.A(n_1205),
.B(n_894),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1180),
.B(n_1146),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1180),
.Y(n_1212)
);

AND2x2_ASAP7_75t_SL g1213 ( 
.A(n_1153),
.B(n_894),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1193),
.Y(n_1214)
);

INVxp67_ASAP7_75t_SL g1215 ( 
.A(n_1193),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1178),
.B(n_1070),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1198),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1161),
.B(n_1045),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1191),
.B(n_1194),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1161),
.B(n_1049),
.Y(n_1220)
);

INVx4_ASAP7_75t_L g1221 ( 
.A(n_1161),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1191),
.A2(n_1075),
.B1(n_1100),
.B2(n_1027),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1198),
.Y(n_1223)
);

NOR2x1p5_ASAP7_75t_L g1224 ( 
.A(n_1157),
.B(n_1017),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1168),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1154),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1168),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_1164),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1170),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1170),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1188),
.B(n_1208),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1207),
.B(n_1073),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1156),
.B(n_1100),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1200),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1181),
.B(n_1053),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1190),
.B(n_1146),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1182),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1197),
.B(n_1082),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1163),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1152),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1167),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1155),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1202),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1169),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1194),
.B(n_1146),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1185),
.B(n_1089),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1162),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1195),
.B(n_1146),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1204),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1195),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1165),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1182),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1199),
.B(n_1146),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1199),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1201),
.B(n_1175),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1175),
.B(n_1086),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1165),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1201),
.A2(n_1101),
.B1(n_1100),
.B2(n_1106),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1176),
.B(n_1086),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1171),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1174),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1176),
.B(n_1106),
.Y(n_1262)
);

INVx5_ASAP7_75t_L g1263 ( 
.A(n_1162),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1177),
.B(n_1037),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1177),
.B(n_1101),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1179),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1183),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1158),
.Y(n_1268)
);

INVx4_ASAP7_75t_L g1269 ( 
.A(n_1184),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1157),
.B(n_1101),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1186),
.Y(n_1271)
);

BUFx4_ASAP7_75t_L g1272 ( 
.A(n_1159),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1159),
.B(n_1101),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1152),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1184),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1172),
.B(n_1016),
.Y(n_1276)
);

AND2x4_ASAP7_75t_SL g1277 ( 
.A(n_1166),
.B(n_1043),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1187),
.B(n_1101),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1184),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1192),
.B(n_1046),
.Y(n_1280)
);

INVx4_ASAP7_75t_L g1281 ( 
.A(n_1184),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1196),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_SL g1283 ( 
.A(n_1160),
.B(n_837),
.Y(n_1283)
);

AND2x6_ASAP7_75t_L g1284 ( 
.A(n_1203),
.B(n_754),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1206),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1184),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1186),
.B(n_1050),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1235),
.Y(n_1288)
);

OR2x6_ASAP7_75t_L g1289 ( 
.A(n_1249),
.B(n_1016),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1231),
.B(n_1189),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1214),
.B(n_1160),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1235),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1232),
.B(n_1173),
.C(n_1172),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1231),
.B(n_1209),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1255),
.B(n_1173),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1221),
.B(n_1092),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1226),
.B(n_1209),
.Y(n_1297)
);

OR2x6_ASAP7_75t_L g1298 ( 
.A(n_1249),
.B(n_1219),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1212),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_L g1300 ( 
.A(n_1238),
.B(n_1048),
.C(n_1041),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1225),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1226),
.B(n_1209),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1233),
.B(n_1209),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1242),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1214),
.B(n_1209),
.Y(n_1305)
);

AND3x1_ASAP7_75t_L g1306 ( 
.A(n_1283),
.B(n_844),
.C(n_774),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1258),
.B(n_1143),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1234),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1255),
.B(n_1139),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1255),
.B(n_1139),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1225),
.Y(n_1311)
);

AND2x6_ASAP7_75t_SL g1312 ( 
.A(n_1264),
.B(n_583),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1255),
.B(n_1139),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1213),
.B(n_674),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1213),
.A2(n_587),
.B1(n_599),
.B2(n_598),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1213),
.A2(n_1248),
.B(n_1253),
.C(n_1212),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1248),
.A2(n_776),
.B(n_822),
.C(n_801),
.Y(n_1317)
);

AND2x2_ASAP7_75t_SL g1318 ( 
.A(n_1210),
.B(n_776),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1215),
.A2(n_655),
.B1(n_782),
.B2(n_576),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1268),
.B(n_911),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1216),
.B(n_911),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1239),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1262),
.B(n_1139),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1227),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1287),
.B(n_1143),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1236),
.B(n_633),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1253),
.A2(n_1129),
.B1(n_841),
.B2(n_1141),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1262),
.B(n_1139),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1227),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1287),
.B(n_1143),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1214),
.B(n_1144),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1236),
.B(n_665),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1214),
.B(n_1106),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1284),
.A2(n_1211),
.B1(n_1274),
.B2(n_1240),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1214),
.B(n_1106),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1265),
.A2(n_801),
.B1(n_872),
.B2(n_822),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1229),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1284),
.A2(n_587),
.B1(n_599),
.B2(n_598),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1229),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1211),
.B(n_1106),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1211),
.B(n_1129),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1228),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1210),
.B(n_1022),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1239),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1211),
.B(n_1131),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1241),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1245),
.A2(n_1141),
.B1(n_816),
.B2(n_838),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1245),
.B(n_1131),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1222),
.B(n_704),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1245),
.B(n_1131),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1245),
.A2(n_1141),
.B1(n_852),
.B2(n_857),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1241),
.B(n_1131),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1219),
.A2(n_1141),
.B1(n_936),
.B2(n_938),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1244),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1219),
.B(n_1144),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1284),
.A2(n_602),
.B1(n_615),
.B2(n_605),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1219),
.B(n_1144),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1262),
.B(n_828),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1250),
.B(n_709),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1230),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1234),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1262),
.B(n_1144),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1210),
.B(n_1060),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1244),
.B(n_1131),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1260),
.Y(n_1365)
);

OAI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1250),
.A2(n_872),
.B1(n_757),
.B2(n_779),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1260),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1270),
.A2(n_1273),
.B(n_1278),
.C(n_1266),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1254),
.B(n_1055),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1230),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1254),
.B(n_1050),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1256),
.B(n_720),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1261),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1261),
.B(n_1131),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1266),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1221),
.B(n_961),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1275),
.B(n_1131),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1267),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1259),
.B(n_784),
.Y(n_1379)
);

NOR3xp33_ASAP7_75t_L g1380 ( 
.A(n_1243),
.B(n_588),
.C(n_586),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1267),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_1276),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1221),
.B(n_1280),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1282),
.B(n_1144),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1246),
.B(n_962),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1275),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1237),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1218),
.B(n_976),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1282),
.B(n_1144),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1285),
.A2(n_1141),
.B1(n_994),
.B2(n_826),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1318),
.B(n_1220),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1301),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1342),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1318),
.B(n_1315),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1315),
.B(n_1277),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1322),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1321),
.A2(n_1285),
.B(n_1276),
.C(n_1237),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1298),
.B(n_1224),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1344),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1303),
.A2(n_1269),
.B(n_1281),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1311),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1321),
.B(n_1240),
.Y(n_1402)
);

OAI321xp33_ASAP7_75t_L g1403 ( 
.A1(n_1314),
.A2(n_805),
.A3(n_909),
.B1(n_912),
.B2(n_844),
.C(n_774),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1314),
.A2(n_1277),
.B1(n_1224),
.B2(n_1284),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1333),
.A2(n_1269),
.B(n_1281),
.Y(n_1405)
);

AOI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1305),
.A2(n_1223),
.B(n_1217),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1346),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_L g1408 ( 
.A(n_1383),
.B(n_1269),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1334),
.A2(n_1223),
.B1(n_1269),
.B2(n_1217),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1386),
.Y(n_1410)
);

NOR2xp67_ASAP7_75t_L g1411 ( 
.A(n_1293),
.B(n_1251),
.Y(n_1411)
);

AOI21xp33_ASAP7_75t_L g1412 ( 
.A1(n_1349),
.A2(n_1257),
.B(n_1251),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1294),
.B(n_1354),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1365),
.B(n_1240),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1335),
.A2(n_1281),
.B(n_1263),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1320),
.B(n_1257),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1367),
.B(n_1274),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1348),
.A2(n_1263),
.B(n_1247),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1373),
.B(n_1274),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1350),
.A2(n_1263),
.B(n_1247),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1316),
.A2(n_912),
.B(n_947),
.C(n_909),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1317),
.A2(n_979),
.B(n_1001),
.C(n_947),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1375),
.B(n_1252),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1290),
.A2(n_1263),
.B(n_1247),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1325),
.A2(n_1263),
.B(n_1247),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1307),
.A2(n_1271),
.B(n_1252),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1330),
.A2(n_1263),
.B(n_1247),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1378),
.B(n_1271),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1341),
.A2(n_1345),
.B(n_1368),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1355),
.A2(n_1247),
.B(n_1275),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1381),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1371),
.B(n_1286),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1304),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1334),
.A2(n_1355),
.B1(n_1357),
.B2(n_1340),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1288),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1299),
.B(n_1284),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1357),
.A2(n_1284),
.B(n_1092),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1362),
.A2(n_1279),
.B(n_1275),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1320),
.B(n_792),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1297),
.A2(n_1279),
.B(n_1275),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1298),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1295),
.A2(n_1284),
.B1(n_1286),
.B2(n_1279),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1369),
.B(n_1279),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1382),
.B(n_1065),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1362),
.A2(n_1286),
.B(n_1279),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1371),
.B(n_1286),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1326),
.B(n_1286),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1326),
.B(n_1098),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1332),
.B(n_1098),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1386),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1324),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1292),
.B(n_797),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1329),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1298),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1349),
.B(n_823),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1337),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1302),
.A2(n_1353),
.B1(n_1327),
.B2(n_1351),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1339),
.Y(n_1458)
);

A2O1A1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1372),
.A2(n_1001),
.B(n_1008),
.C(n_979),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1305),
.A2(n_1162),
.B(n_1094),
.Y(n_1460)
);

OR2x6_ASAP7_75t_L g1461 ( 
.A(n_1361),
.B(n_1272),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1360),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1332),
.B(n_1108),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1336),
.A2(n_1379),
.B1(n_1372),
.B2(n_1363),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1331),
.A2(n_1094),
.B(n_1102),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1331),
.A2(n_1094),
.B(n_1102),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1370),
.B(n_1108),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1366),
.B(n_608),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1289),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1379),
.B(n_834),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1309),
.A2(n_1094),
.B(n_1103),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1308),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1387),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1319),
.A2(n_1291),
.B(n_1388),
.C(n_1380),
.Y(n_1474)
);

OAI21xp33_ASAP7_75t_L g1475 ( 
.A1(n_1359),
.A2(n_1300),
.B(n_1343),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1352),
.A2(n_1107),
.B(n_1103),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1364),
.A2(n_1107),
.B(n_1103),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1291),
.B(n_1099),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1359),
.B(n_1099),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1338),
.B(n_1112),
.Y(n_1480)
);

AND2x2_ASAP7_75t_SL g1481 ( 
.A(n_1306),
.B(n_1272),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1374),
.A2(n_1110),
.B(n_1107),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1338),
.B(n_1356),
.Y(n_1483)
);

AOI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1384),
.A2(n_1135),
.B(n_1124),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1289),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1389),
.A2(n_1110),
.B(n_1144),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1385),
.A2(n_1008),
.B(n_602),
.C(n_615),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1377),
.A2(n_1110),
.B(n_1150),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1429),
.A2(n_1296),
.B(n_1310),
.Y(n_1489)
);

NAND2x1p5_ASAP7_75t_L g1490 ( 
.A(n_1441),
.B(n_1313),
.Y(n_1490)
);

A2O1A1Ixp33_ASAP7_75t_SL g1491 ( 
.A1(n_1416),
.A2(n_1390),
.B(n_1347),
.C(n_1356),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1429),
.A2(n_1296),
.B(n_1323),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1394),
.A2(n_1289),
.B1(n_875),
.B2(n_878),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1475),
.B(n_1358),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1410),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1396),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1399),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1413),
.B(n_1377),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1400),
.A2(n_1328),
.B(n_1376),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1398),
.B(n_1074),
.Y(n_1500)
);

AO32x1_ASAP7_75t_L g1501 ( 
.A1(n_1457),
.A2(n_1409),
.A3(n_1434),
.B1(n_1431),
.B2(n_1407),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_SL g1502 ( 
.A(n_1470),
.B(n_916),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1405),
.A2(n_1094),
.B(n_1150),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1402),
.A2(n_1150),
.B(n_1104),
.Y(n_1504)
);

A2O1A1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1474),
.A2(n_596),
.B(n_716),
.C(n_658),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1393),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1406),
.A2(n_1137),
.B(n_1135),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1464),
.B(n_1312),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1433),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1415),
.A2(n_1150),
.B(n_1104),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1451),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1448),
.B(n_597),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1461),
.Y(n_1513)
);

NOR2xp67_ASAP7_75t_SL g1514 ( 
.A(n_1485),
.B(n_789),
.Y(n_1514)
);

OR2x6_ASAP7_75t_L g1515 ( 
.A(n_1461),
.B(n_826),
.Y(n_1515)
);

AO22x1_ASAP7_75t_L g1516 ( 
.A1(n_1455),
.A2(n_635),
.B1(n_661),
.B2(n_611),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1472),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1453),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1427),
.A2(n_1150),
.B(n_1104),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1392),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1461),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1456),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1452),
.B(n_1081),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1449),
.B(n_670),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1469),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1463),
.B(n_679),
.Y(n_1526)
);

BUFx8_ASAP7_75t_SL g1527 ( 
.A(n_1398),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1462),
.Y(n_1528)
);

INVx2_ASAP7_75t_SL g1529 ( 
.A(n_1435),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1425),
.A2(n_1150),
.B(n_1104),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1425),
.A2(n_1150),
.B(n_1104),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1441),
.Y(n_1532)
);

AOI33xp33_ASAP7_75t_L g1533 ( 
.A1(n_1487),
.A2(n_843),
.A3(n_719),
.B1(n_850),
.B2(n_756),
.B3(n_686),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1412),
.B(n_835),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1401),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1439),
.A2(n_1391),
.B1(n_1395),
.B2(n_1404),
.Y(n_1536)
);

NOR2xp67_ASAP7_75t_SL g1537 ( 
.A(n_1441),
.B(n_658),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1479),
.B(n_966),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1458),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1483),
.A2(n_943),
.B1(n_950),
.B2(n_921),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1473),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1454),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1468),
.A2(n_981),
.B(n_605),
.C(n_618),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1443),
.B(n_580),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1424),
.A2(n_1104),
.B(n_1097),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1444),
.B(n_621),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1423),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1454),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1428),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1424),
.A2(n_1104),
.B(n_1097),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1454),
.B(n_1112),
.Y(n_1551)
);

A2O1A1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1397),
.A2(n_743),
.B(n_811),
.C(n_716),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1410),
.Y(n_1553)
);

AOI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1484),
.A2(n_1138),
.B(n_1137),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1450),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1447),
.B(n_584),
.Y(n_1556)
);

OAI21xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1436),
.A2(n_618),
.B(n_617),
.Y(n_1557)
);

AO31x2_ASAP7_75t_L g1558 ( 
.A1(n_1440),
.A2(n_1140),
.A3(n_1138),
.B(n_1114),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1418),
.A2(n_1105),
.B(n_1097),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1467),
.Y(n_1560)
);

AND2x6_ASAP7_75t_SL g1561 ( 
.A(n_1411),
.B(n_617),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1459),
.B(n_589),
.Y(n_1562)
);

BUFx12f_ASAP7_75t_L g1563 ( 
.A(n_1481),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1414),
.B(n_1090),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1417),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1419),
.B(n_1090),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1420),
.A2(n_1105),
.B(n_1097),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1432),
.B(n_594),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1450),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1478),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1442),
.A2(n_1480),
.B1(n_1446),
.B2(n_1421),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1408),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1403),
.Y(n_1573)
);

BUFx12f_ASAP7_75t_L g1574 ( 
.A(n_1422),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1438),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1440),
.A2(n_1109),
.B(n_1105),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1426),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1445),
.B(n_953),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_SL g1579 ( 
.A1(n_1437),
.A2(n_1114),
.B(n_1125),
.C(n_1113),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1430),
.A2(n_1486),
.B(n_1477),
.Y(n_1580)
);

NOR2xp67_ASAP7_75t_L g1581 ( 
.A(n_1471),
.B(n_529),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1488),
.Y(n_1582)
);

A2O1A1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1486),
.A2(n_811),
.B(n_818),
.C(n_743),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1476),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1488),
.B(n_969),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1460),
.A2(n_971),
.B1(n_988),
.B2(n_993),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1476),
.A2(n_637),
.B1(n_650),
.B2(n_593),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1477),
.B(n_1482),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1482),
.A2(n_600),
.B1(n_604),
.B2(n_601),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1465),
.A2(n_1109),
.B(n_1105),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1489),
.A2(n_1466),
.B(n_874),
.Y(n_1591)
);

O2A1O1Ixp33_ASAP7_75t_SL g1592 ( 
.A1(n_1491),
.A2(n_622),
.B(n_624),
.C(n_623),
.Y(n_1592)
);

AOI221x1_ASAP7_75t_L g1593 ( 
.A1(n_1578),
.A2(n_622),
.B1(n_627),
.B2(n_624),
.C(n_623),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1570),
.B(n_1113),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1506),
.Y(n_1595)
);

AO31x2_ASAP7_75t_L g1596 ( 
.A1(n_1580),
.A2(n_637),
.A3(n_650),
.B(n_593),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1527),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1502),
.B(n_606),
.Y(n_1598)
);

AOI21x1_ASAP7_75t_L g1599 ( 
.A1(n_1554),
.A2(n_1140),
.B(n_1132),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1496),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1523),
.B(n_608),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1520),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1547),
.B(n_1125),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1565),
.B(n_1132),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1588),
.A2(n_1134),
.B(n_1128),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1517),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1525),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1571),
.A2(n_1134),
.B(n_1128),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1509),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1512),
.B(n_607),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1542),
.B(n_627),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1549),
.B(n_631),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1502),
.B(n_609),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1534),
.A2(n_1508),
.B1(n_1536),
.B2(n_1516),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1492),
.A2(n_1121),
.B(n_1120),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1497),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1499),
.A2(n_874),
.B(n_1115),
.Y(n_1617)
);

AO32x2_ASAP7_75t_L g1618 ( 
.A1(n_1540),
.A2(n_812),
.A3(n_888),
.B1(n_685),
.B2(n_621),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1501),
.A2(n_874),
.B(n_1115),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1584),
.A2(n_1042),
.B(n_1040),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1503),
.A2(n_1121),
.B(n_1120),
.Y(n_1621)
);

NAND3xp33_ASAP7_75t_L g1622 ( 
.A(n_1586),
.B(n_613),
.C(n_612),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1576),
.A2(n_1121),
.B(n_1120),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1501),
.A2(n_874),
.B(n_1115),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1529),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1555),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1511),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1501),
.A2(n_874),
.B(n_1118),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1573),
.B(n_1546),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1571),
.A2(n_1118),
.B(n_1122),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1518),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1555),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1498),
.B(n_631),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1522),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1528),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1532),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1548),
.Y(n_1637)
);

AO32x2_ASAP7_75t_L g1638 ( 
.A1(n_1540),
.A2(n_812),
.A3(n_888),
.B1(n_685),
.B2(n_621),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1530),
.A2(n_1122),
.B(n_1042),
.Y(n_1639)
);

AO31x2_ASAP7_75t_L g1640 ( 
.A1(n_1577),
.A2(n_697),
.A3(n_729),
.B(n_664),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1500),
.B(n_632),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_SL g1642 ( 
.A(n_1543),
.B(n_616),
.C(n_614),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1535),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1539),
.Y(n_1644)
);

INVx4_ASAP7_75t_L g1645 ( 
.A(n_1555),
.Y(n_1645)
);

AO21x1_ASAP7_75t_L g1646 ( 
.A1(n_1494),
.A2(n_638),
.B(n_632),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1531),
.A2(n_1122),
.B(n_1047),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1579),
.A2(n_1118),
.B(n_1109),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1507),
.A2(n_1047),
.B(n_1040),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1585),
.A2(n_648),
.B(n_638),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1500),
.B(n_608),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1498),
.A2(n_1118),
.B(n_1109),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1560),
.B(n_648),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1541),
.B(n_652),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_SL g1655 ( 
.A1(n_1587),
.A2(n_697),
.B(n_664),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1505),
.B(n_652),
.Y(n_1656)
);

A2O1A1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1552),
.A2(n_1557),
.B(n_1533),
.C(n_1562),
.Y(n_1657)
);

OA21x2_ASAP7_75t_L g1658 ( 
.A1(n_1583),
.A2(n_1052),
.B(n_1051),
.Y(n_1658)
);

AO21x1_ASAP7_75t_L g1659 ( 
.A1(n_1556),
.A2(n_659),
.B(n_654),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1553),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1524),
.B(n_654),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1575),
.A2(n_1118),
.B(n_1052),
.Y(n_1662)
);

AOI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1545),
.A2(n_1054),
.B(n_1051),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1544),
.B(n_659),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1569),
.B(n_668),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_SL g1666 ( 
.A1(n_1587),
.A2(n_765),
.B(n_729),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1526),
.B(n_668),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1575),
.A2(n_1118),
.B(n_1057),
.Y(n_1668)
);

O2A1O1Ixp5_ASAP7_75t_L g1669 ( 
.A1(n_1537),
.A2(n_669),
.B(n_678),
.C(n_673),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1568),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1493),
.A2(n_917),
.B1(n_924),
.B2(n_818),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_SL g1672 ( 
.A1(n_1493),
.A2(n_1538),
.B(n_1589),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1551),
.B(n_1574),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1616),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1627),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1614),
.A2(n_1515),
.B1(n_1563),
.B2(n_1521),
.Y(n_1676)
);

OAI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1672),
.A2(n_1593),
.B1(n_1622),
.B2(n_1671),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1615),
.A2(n_1591),
.B(n_1617),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1673),
.B(n_1515),
.Y(n_1679)
);

OA21x2_ASAP7_75t_L g1680 ( 
.A1(n_1619),
.A2(n_1567),
.B(n_1559),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1597),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1598),
.A2(n_1581),
.B(n_1490),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1596),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1608),
.A2(n_1510),
.B(n_1572),
.Y(n_1684)
);

A2O1A1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1672),
.A2(n_924),
.B(n_917),
.C(n_770),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1649),
.A2(n_1519),
.B(n_1550),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1613),
.A2(n_1490),
.B(n_1551),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1631),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1599),
.A2(n_1504),
.B(n_1590),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1670),
.B(n_1513),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1634),
.B(n_1572),
.Y(n_1691)
);

AO21x1_ASAP7_75t_L g1692 ( 
.A1(n_1650),
.A2(n_673),
.B(n_669),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1595),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1606),
.B(n_1633),
.Y(n_1694)
);

INVx2_ASAP7_75t_SL g1695 ( 
.A(n_1607),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_SL g1696 ( 
.A1(n_1608),
.A2(n_1514),
.B(n_1495),
.C(n_770),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1663),
.A2(n_1566),
.B(n_1564),
.Y(n_1697)
);

AOI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1671),
.A2(n_681),
.B(n_684),
.C(n_678),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1622),
.A2(n_1515),
.B1(n_1495),
.B2(n_620),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1629),
.B(n_608),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1635),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1645),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1659),
.B(n_1582),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1633),
.B(n_1561),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1624),
.A2(n_1566),
.B(n_1564),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1645),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1621),
.A2(n_1558),
.B(n_1582),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1600),
.B(n_1558),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_1637),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1650),
.A2(n_781),
.B(n_824),
.C(n_765),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1642),
.A2(n_685),
.B1(n_812),
.B2(n_621),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1646),
.B(n_1582),
.Y(n_1712)
);

OAI21x1_ASAP7_75t_L g1713 ( 
.A1(n_1652),
.A2(n_1558),
.B(n_1057),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1625),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1643),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1665),
.B(n_1007),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_SL g1717 ( 
.A1(n_1601),
.A2(n_812),
.B1(n_888),
.B2(n_685),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1644),
.Y(n_1718)
);

AOI22x1_ASAP7_75t_L g1719 ( 
.A1(n_1664),
.A2(n_626),
.B1(n_628),
.B2(n_625),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1636),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1628),
.A2(n_684),
.B(n_681),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1640),
.Y(n_1722)
);

OAI21x1_ASAP7_75t_L g1723 ( 
.A1(n_1623),
.A2(n_1058),
.B(n_1054),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1658),
.B(n_689),
.Y(n_1724)
);

INVx2_ASAP7_75t_R g1725 ( 
.A(n_1660),
.Y(n_1725)
);

AOI21x1_ASAP7_75t_L g1726 ( 
.A1(n_1656),
.A2(n_690),
.B(n_689),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1596),
.Y(n_1727)
);

NAND2x1p5_ASAP7_75t_L g1728 ( 
.A(n_1658),
.B(n_690),
.Y(n_1728)
);

CKINVDCx11_ASAP7_75t_R g1729 ( 
.A(n_1609),
.Y(n_1729)
);

OA21x2_ASAP7_75t_L g1730 ( 
.A1(n_1630),
.A2(n_698),
.B(n_692),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1640),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1640),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1596),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1694),
.B(n_1602),
.Y(n_1734)
);

CKINVDCx11_ASAP7_75t_R g1735 ( 
.A(n_1709),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1689),
.A2(n_1656),
.B(n_1657),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1691),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1674),
.B(n_1605),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1722),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1684),
.A2(n_1592),
.B(n_1605),
.Y(n_1740)
);

AOI21xp33_ASAP7_75t_SL g1741 ( 
.A1(n_1676),
.A2(n_1651),
.B(n_1610),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1675),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1691),
.B(n_1626),
.Y(n_1743)
);

A2O1A1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1698),
.A2(n_1669),
.B(n_1667),
.C(n_1661),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1682),
.A2(n_1668),
.B(n_1662),
.Y(n_1745)
);

BUFx12f_ASAP7_75t_L g1746 ( 
.A(n_1681),
.Y(n_1746)
);

AO21x2_ASAP7_75t_L g1747 ( 
.A1(n_1731),
.A2(n_1666),
.B(n_1655),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1715),
.B(n_1718),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1688),
.B(n_1665),
.Y(n_1749)
);

OAI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1677),
.A2(n_1667),
.B(n_1661),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1677),
.A2(n_1641),
.B1(n_1611),
.B2(n_1654),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1683),
.B(n_1612),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1676),
.A2(n_1711),
.B1(n_1704),
.B2(n_1717),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1691),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1711),
.A2(n_1641),
.B1(n_1611),
.B2(n_1654),
.Y(n_1755)
);

OA21x2_ASAP7_75t_L g1756 ( 
.A1(n_1689),
.A2(n_1648),
.B(n_1647),
.Y(n_1756)
);

INVx5_ASAP7_75t_L g1757 ( 
.A(n_1724),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1732),
.Y(n_1758)
);

INVx4_ASAP7_75t_L g1759 ( 
.A(n_1679),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1687),
.B(n_1653),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1708),
.Y(n_1761)
);

OAI21x1_ASAP7_75t_L g1762 ( 
.A1(n_1678),
.A2(n_1639),
.B(n_1620),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1703),
.A2(n_1620),
.B(n_1604),
.Y(n_1763)
);

OA21x2_ASAP7_75t_L g1764 ( 
.A1(n_1727),
.A2(n_1594),
.B(n_1604),
.Y(n_1764)
);

OAI21x1_ASAP7_75t_L g1765 ( 
.A1(n_1678),
.A2(n_1594),
.B(n_1603),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1701),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1714),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1683),
.B(n_1618),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1679),
.A2(n_1653),
.B1(n_1612),
.B2(n_630),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1714),
.B(n_1626),
.Y(n_1770)
);

A2O1A1Ixp33_ASAP7_75t_L g1771 ( 
.A1(n_1685),
.A2(n_1638),
.B(n_1618),
.C(n_698),
.Y(n_1771)
);

OR2x2_ASAP7_75t_SL g1772 ( 
.A(n_1727),
.B(n_1618),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1679),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1733),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_1702),
.Y(n_1775)
);

OAI21x1_ASAP7_75t_L g1776 ( 
.A1(n_1686),
.A2(n_1603),
.B(n_1632),
.Y(n_1776)
);

AO31x2_ASAP7_75t_L g1777 ( 
.A1(n_1733),
.A2(n_824),
.A3(n_871),
.B(n_781),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1705),
.Y(n_1778)
);

OAI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1685),
.A2(n_701),
.B(n_692),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1695),
.B(n_1632),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1690),
.B(n_629),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1703),
.A2(n_1638),
.B(n_922),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1777),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1761),
.B(n_1705),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1777),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1773),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1738),
.B(n_1705),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1739),
.Y(n_1788)
);

OAI21x1_ASAP7_75t_L g1789 ( 
.A1(n_1778),
.A2(n_1707),
.B(n_1713),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1739),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1758),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1758),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_1737),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1761),
.B(n_1725),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1777),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1777),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1750),
.A2(n_1710),
.B(n_1726),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1777),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1778),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1774),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1742),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1776),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1773),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1774),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1738),
.B(n_1725),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1768),
.B(n_1680),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1742),
.Y(n_1807)
);

AO21x2_ASAP7_75t_L g1808 ( 
.A1(n_1740),
.A2(n_1696),
.B(n_1710),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1766),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1766),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1764),
.Y(n_1811)
);

OAI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1744),
.A2(n_1696),
.B(n_1699),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1748),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1764),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1776),
.Y(n_1815)
);

AO21x2_ASAP7_75t_L g1816 ( 
.A1(n_1762),
.A2(n_1692),
.B(n_1697),
.Y(n_1816)
);

AOI21x1_ASAP7_75t_L g1817 ( 
.A1(n_1782),
.A2(n_1724),
.B(n_1730),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1764),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1764),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1736),
.Y(n_1820)
);

BUFx5_ASAP7_75t_L g1821 ( 
.A(n_1768),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1772),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1772),
.Y(n_1823)
);

INVx4_ASAP7_75t_L g1824 ( 
.A(n_1757),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1752),
.Y(n_1825)
);

OAI21x1_ASAP7_75t_L g1826 ( 
.A1(n_1762),
.A2(n_1765),
.B(n_1745),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1754),
.B(n_1680),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1736),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1736),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1752),
.Y(n_1830)
);

AO21x2_ASAP7_75t_L g1831 ( 
.A1(n_1763),
.A2(n_1697),
.B(n_1723),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1734),
.B(n_1721),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1754),
.Y(n_1833)
);

AO21x2_ASAP7_75t_L g1834 ( 
.A1(n_1771),
.A2(n_703),
.B(n_701),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1736),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1754),
.Y(n_1836)
);

CKINVDCx16_ASAP7_75t_R g1837 ( 
.A(n_1803),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1788),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1812),
.A2(n_1753),
.B1(n_1759),
.B2(n_1773),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1821),
.B(n_1822),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1788),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1822),
.B(n_1767),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1821),
.B(n_1754),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1799),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1812),
.A2(n_1759),
.B1(n_1773),
.B2(n_1760),
.Y(n_1845)
);

NAND3xp33_ASAP7_75t_L g1846 ( 
.A(n_1797),
.B(n_1741),
.C(n_1779),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1797),
.A2(n_1757),
.B1(n_1759),
.B2(n_1773),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1788),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1799),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1799),
.Y(n_1850)
);

OAI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1822),
.A2(n_1769),
.B1(n_1751),
.B2(n_1781),
.C(n_1755),
.Y(n_1851)
);

OAI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1823),
.A2(n_1719),
.B1(n_1749),
.B2(n_1700),
.C(n_708),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1824),
.B(n_1754),
.Y(n_1853)
);

AO221x2_ASAP7_75t_L g1854 ( 
.A1(n_1823),
.A2(n_1638),
.B1(n_845),
.B2(n_856),
.C(n_766),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1823),
.A2(n_708),
.B1(n_710),
.B2(n_705),
.C(n_703),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1821),
.B(n_1767),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1803),
.A2(n_1757),
.B1(n_1709),
.B2(n_1743),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1799),
.Y(n_1858)
);

AOI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1813),
.A2(n_712),
.B1(n_724),
.B2(n_710),
.C(n_705),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1821),
.B(n_1743),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_SL g1861 ( 
.A1(n_1834),
.A2(n_1757),
.B1(n_1746),
.B2(n_1743),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1813),
.B(n_1770),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1834),
.A2(n_1757),
.B1(n_1729),
.B2(n_1735),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1821),
.B(n_1775),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1790),
.Y(n_1865)
);

OAI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1826),
.A2(n_1765),
.B(n_1756),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1834),
.A2(n_1746),
.B1(n_1730),
.B2(n_1716),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1808),
.A2(n_1712),
.B(n_1730),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1840),
.B(n_1821),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1838),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1840),
.B(n_1824),
.Y(n_1871)
);

INVxp67_ASAP7_75t_SL g1872 ( 
.A(n_1858),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1838),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1858),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1843),
.B(n_1824),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1843),
.B(n_1821),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1858),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1841),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1841),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1858),
.B(n_1821),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1860),
.B(n_1821),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1860),
.B(n_1821),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1848),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1853),
.B(n_1824),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1864),
.B(n_1821),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1864),
.B(n_1821),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1844),
.B(n_1821),
.Y(n_1887)
);

AND2x4_ASAP7_75t_L g1888 ( 
.A(n_1853),
.B(n_1824),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1848),
.Y(n_1889)
);

BUFx4f_ASAP7_75t_L g1890 ( 
.A(n_1853),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1865),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1844),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1865),
.Y(n_1893)
);

BUFx3_ASAP7_75t_L g1894 ( 
.A(n_1853),
.Y(n_1894)
);

BUFx2_ASAP7_75t_L g1895 ( 
.A(n_1856),
.Y(n_1895)
);

INVxp67_ASAP7_75t_SL g1896 ( 
.A(n_1844),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1850),
.B(n_1821),
.Y(n_1897)
);

INVx6_ASAP7_75t_L g1898 ( 
.A(n_1837),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1850),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1884),
.B(n_1862),
.Y(n_1900)
);

INVx4_ASAP7_75t_L g1901 ( 
.A(n_1898),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1870),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1890),
.B(n_1837),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1870),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1884),
.B(n_1813),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1873),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1898),
.B(n_1735),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1873),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1892),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1894),
.B(n_1850),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1898),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1878),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1878),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1879),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1890),
.B(n_1856),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1884),
.B(n_1854),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1890),
.B(n_1842),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1879),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1890),
.B(n_1842),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1883),
.B(n_1825),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1883),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1889),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1894),
.B(n_1803),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1890),
.B(n_1803),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1889),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1891),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1891),
.Y(n_1927)
);

AOI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1899),
.A2(n_1849),
.B(n_1814),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1898),
.B(n_1786),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1894),
.B(n_1819),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1893),
.Y(n_1931)
);

BUFx2_ASAP7_75t_SL g1932 ( 
.A(n_1894),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1904),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1900),
.B(n_1895),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1916),
.B(n_1895),
.Y(n_1935)
);

AOI33xp33_ASAP7_75t_L g1936 ( 
.A1(n_1903),
.A2(n_731),
.A3(n_724),
.B1(n_734),
.B2(n_727),
.B3(n_712),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1921),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1931),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1902),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1902),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1906),
.Y(n_1941)
);

AOI221xp5_ASAP7_75t_L g1942 ( 
.A1(n_1901),
.A2(n_1846),
.B1(n_1855),
.B2(n_1851),
.C(n_1852),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1906),
.Y(n_1943)
);

OAI211xp5_ASAP7_75t_L g1944 ( 
.A1(n_1901),
.A2(n_1846),
.B(n_1839),
.C(n_1845),
.Y(n_1944)
);

AOI33xp33_ASAP7_75t_L g1945 ( 
.A1(n_1903),
.A2(n_736),
.A3(n_731),
.B1(n_740),
.B2(n_734),
.B3(n_727),
.Y(n_1945)
);

AND3x1_ASAP7_75t_L g1946 ( 
.A(n_1907),
.B(n_1911),
.C(n_1924),
.Y(n_1946)
);

OAI211xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1911),
.A2(n_1859),
.B(n_1863),
.C(n_1729),
.Y(n_1947)
);

OAI31xp33_ASAP7_75t_L g1948 ( 
.A1(n_1911),
.A2(n_1847),
.A3(n_1888),
.B(n_1884),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1910),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1908),
.Y(n_1950)
);

AND2x4_ASAP7_75t_SL g1951 ( 
.A(n_1901),
.B(n_1888),
.Y(n_1951)
);

OAI31xp33_ASAP7_75t_SL g1952 ( 
.A1(n_1917),
.A2(n_1861),
.A3(n_1888),
.B(n_1884),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1901),
.B(n_1888),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1908),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1912),
.Y(n_1955)
);

AO221x2_ASAP7_75t_L g1956 ( 
.A1(n_1932),
.A2(n_1857),
.B1(n_1854),
.B2(n_1898),
.C(n_747),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1924),
.B(n_1898),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1917),
.B(n_1888),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1910),
.Y(n_1959)
);

NAND3xp33_ASAP7_75t_L g1960 ( 
.A(n_1905),
.B(n_1854),
.C(n_1867),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1912),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1919),
.B(n_1895),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1910),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1935),
.B(n_1919),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1957),
.B(n_1915),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1951),
.Y(n_1966)
);

INVxp67_ASAP7_75t_L g1967 ( 
.A(n_1938),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1962),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1944),
.B(n_1681),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1942),
.B(n_1929),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1960),
.A2(n_1929),
.B(n_1923),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1936),
.B(n_1923),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1951),
.B(n_1932),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1938),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1955),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1934),
.B(n_1920),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1955),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1939),
.Y(n_1978)
);

NAND2xp67_ASAP7_75t_L g1979 ( 
.A(n_1949),
.B(n_1915),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1933),
.B(n_1923),
.Y(n_1980)
);

NAND3xp33_ASAP7_75t_L g1981 ( 
.A(n_1952),
.B(n_1854),
.C(n_1930),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1958),
.B(n_1953),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1958),
.B(n_1923),
.Y(n_1983)
);

NOR2xp67_ASAP7_75t_SL g1984 ( 
.A(n_1937),
.B(n_1693),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1940),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1949),
.Y(n_1986)
);

INVx1_ASAP7_75t_SL g1987 ( 
.A(n_1953),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1959),
.Y(n_1988)
);

AND2x4_ASAP7_75t_L g1989 ( 
.A(n_1958),
.B(n_1913),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1953),
.B(n_1871),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1941),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1943),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1950),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1956),
.B(n_1920),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1946),
.B(n_1871),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1954),
.Y(n_1996)
);

AND2x4_ASAP7_75t_L g1997 ( 
.A(n_1959),
.B(n_1913),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1961),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1963),
.B(n_1948),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1936),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1945),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1945),
.Y(n_2002)
);

OR2x6_ASAP7_75t_L g2003 ( 
.A(n_1963),
.B(n_1720),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1956),
.B(n_1871),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1956),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1947),
.B(n_1914),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1957),
.B(n_1875),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1967),
.Y(n_2008)
);

INVx1_ASAP7_75t_SL g2009 ( 
.A(n_1973),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_2000),
.B(n_1910),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1968),
.B(n_1914),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_2001),
.B(n_1875),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1965),
.B(n_1930),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1968),
.B(n_1918),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1982),
.B(n_1930),
.Y(n_2015)
);

BUFx2_ASAP7_75t_SL g2016 ( 
.A(n_1973),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1995),
.B(n_1983),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1995),
.B(n_1930),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1967),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1966),
.B(n_1871),
.Y(n_2020)
);

INVxp67_ASAP7_75t_L g2021 ( 
.A(n_1969),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1989),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1989),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1989),
.B(n_1918),
.Y(n_2024)
);

INVxp67_ASAP7_75t_SL g2025 ( 
.A(n_2005),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1990),
.B(n_1871),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1979),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1994),
.Y(n_2028)
);

INVxp67_ASAP7_75t_L g2029 ( 
.A(n_1969),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1975),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1990),
.B(n_2004),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_2002),
.B(n_1922),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2004),
.B(n_1875),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_2003),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2005),
.B(n_1922),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1977),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1974),
.B(n_1925),
.Y(n_2037)
);

INVxp33_ASAP7_75t_SL g2038 ( 
.A(n_1984),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_2003),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1999),
.B(n_1875),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1999),
.B(n_1875),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1986),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1987),
.B(n_1869),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_1970),
.A2(n_1926),
.B(n_1925),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_2007),
.B(n_1869),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2007),
.B(n_1869),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1986),
.B(n_1926),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1980),
.B(n_1927),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1980),
.B(n_1927),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1972),
.B(n_1887),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1964),
.B(n_1887),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1988),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_2003),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1997),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1971),
.B(n_2006),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1988),
.B(n_1887),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_1976),
.B(n_1909),
.Y(n_2057)
);

BUFx6f_ASAP7_75t_L g2058 ( 
.A(n_1997),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_2006),
.B(n_1881),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1978),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1985),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1991),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1992),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1993),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1996),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1998),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_1997),
.Y(n_2067)
);

INVx1_ASAP7_75t_SL g2068 ( 
.A(n_2006),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_1981),
.B(n_1909),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1967),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2000),
.B(n_1897),
.Y(n_2071)
);

OAI21xp5_ASAP7_75t_SL g2072 ( 
.A1(n_2055),
.A2(n_740),
.B(n_736),
.Y(n_2072)
);

CKINVDCx16_ASAP7_75t_R g2073 ( 
.A(n_2028),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_2010),
.B(n_1897),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2009),
.B(n_2069),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2058),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2067),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_2038),
.B(n_1882),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2023),
.Y(n_2079)
);

OAI21xp33_ASAP7_75t_L g2080 ( 
.A1(n_2055),
.A2(n_1897),
.B(n_1882),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2008),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_2022),
.B(n_1881),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2021),
.B(n_1876),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2029),
.B(n_1876),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2058),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2058),
.Y(n_2086)
);

AOI322xp5_ASAP7_75t_L g2087 ( 
.A1(n_2068),
.A2(n_1872),
.A3(n_764),
.B1(n_766),
.B2(n_759),
.C1(n_771),
.C2(n_762),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2058),
.Y(n_2088)
);

AOI221xp5_ASAP7_75t_L g2089 ( 
.A1(n_2044),
.A2(n_762),
.B1(n_764),
.B2(n_759),
.C(n_747),
.Y(n_2089)
);

NAND3xp33_ASAP7_75t_SL g2090 ( 
.A(n_2069),
.B(n_641),
.C(n_640),
.Y(n_2090)
);

OAI21xp33_ASAP7_75t_L g2091 ( 
.A1(n_2012),
.A2(n_2070),
.B(n_2019),
.Y(n_2091)
);

AOI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_2038),
.A2(n_1824),
.B1(n_1834),
.B2(n_1868),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2017),
.B(n_1881),
.Y(n_2093)
);

AOI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_2016),
.A2(n_1834),
.B1(n_773),
.B2(n_785),
.Y(n_2094)
);

INVxp67_ASAP7_75t_L g2095 ( 
.A(n_2016),
.Y(n_2095)
);

A2O1A1Ixp33_ASAP7_75t_L g2096 ( 
.A1(n_2059),
.A2(n_832),
.B(n_859),
.C(n_795),
.Y(n_2096)
);

OAI21xp33_ASAP7_75t_SL g2097 ( 
.A1(n_2025),
.A2(n_1882),
.B(n_1872),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2032),
.A2(n_773),
.B1(n_785),
.B2(n_771),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_2017),
.A2(n_1876),
.B1(n_1886),
.B2(n_1885),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2058),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2031),
.B(n_1885),
.Y(n_2101)
);

OAI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2040),
.A2(n_1885),
.B1(n_1886),
.B2(n_1880),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2054),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2027),
.B(n_1886),
.Y(n_2104)
);

OAI211xp5_ASAP7_75t_L g2105 ( 
.A1(n_2027),
.A2(n_2071),
.B(n_2030),
.C(n_2036),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_SL g2106 ( 
.A(n_2040),
.B(n_1786),
.Y(n_2106)
);

CKINVDCx16_ASAP7_75t_R g2107 ( 
.A(n_2041),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2050),
.B(n_1892),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2031),
.B(n_2041),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2015),
.B(n_1880),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2054),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2022),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2035),
.B(n_1892),
.Y(n_2113)
);

AOI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2060),
.A2(n_795),
.B1(n_798),
.B2(n_787),
.Y(n_2114)
);

AOI32xp33_ASAP7_75t_L g2115 ( 
.A1(n_2020),
.A2(n_2018),
.A3(n_2015),
.B1(n_2013),
.B2(n_2043),
.Y(n_2115)
);

OAI21xp33_ASAP7_75t_L g2116 ( 
.A1(n_2020),
.A2(n_1880),
.B(n_1896),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2042),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2018),
.Y(n_2118)
);

BUFx2_ASAP7_75t_L g2119 ( 
.A(n_2024),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2033),
.B(n_2013),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2052),
.Y(n_2121)
);

INVx2_ASAP7_75t_SL g2122 ( 
.A(n_2033),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2026),
.B(n_1893),
.Y(n_2123)
);

OAI32xp33_ASAP7_75t_L g2124 ( 
.A1(n_2034),
.A2(n_1877),
.A3(n_1874),
.B1(n_1829),
.B2(n_1835),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2026),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2048),
.B(n_1896),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2011),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2048),
.B(n_1899),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2049),
.B(n_1899),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2024),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2049),
.B(n_787),
.Y(n_2131)
);

OR3x1_ASAP7_75t_L g2132 ( 
.A(n_2061),
.B(n_799),
.C(n_798),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_2024),
.Y(n_2133)
);

AOI322xp5_ASAP7_75t_L g2134 ( 
.A1(n_2062),
.A2(n_2065),
.A3(n_2064),
.B1(n_2066),
.B2(n_2063),
.C1(n_2043),
.C2(n_2046),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2034),
.B(n_799),
.Y(n_2135)
);

INVx2_ASAP7_75t_SL g2136 ( 
.A(n_2039),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2011),
.Y(n_2137)
);

INVx1_ASAP7_75t_SL g2138 ( 
.A(n_2014),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2014),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_2039),
.A2(n_1786),
.B1(n_1830),
.B2(n_1825),
.Y(n_2140)
);

HB1xp67_ASAP7_75t_L g2141 ( 
.A(n_2053),
.Y(n_2141)
);

INVx1_ASAP7_75t_SL g2142 ( 
.A(n_2053),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2047),
.Y(n_2143)
);

AOI32xp33_ASAP7_75t_L g2144 ( 
.A1(n_2045),
.A2(n_829),
.A3(n_831),
.B1(n_821),
.B2(n_813),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2045),
.B(n_2046),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2037),
.B(n_813),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2037),
.B(n_821),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2047),
.Y(n_2148)
);

AOI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_2051),
.A2(n_831),
.B1(n_832),
.B2(n_829),
.Y(n_2149)
);

NAND3xp33_ASAP7_75t_L g2150 ( 
.A(n_2057),
.B(n_840),
.C(n_836),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2057),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2056),
.B(n_836),
.Y(n_2152)
);

HB1xp67_ASAP7_75t_L g2153 ( 
.A(n_2058),
.Y(n_2153)
);

AND2x4_ASAP7_75t_L g2154 ( 
.A(n_2023),
.B(n_1928),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2058),
.Y(n_2155)
);

NAND2xp33_ASAP7_75t_SL g2156 ( 
.A(n_2017),
.B(n_1780),
.Y(n_2156)
);

INVx1_ASAP7_75t_SL g2157 ( 
.A(n_2016),
.Y(n_2157)
);

OAI311xp33_ASAP7_75t_L g2158 ( 
.A1(n_2021),
.A2(n_848),
.A3(n_849),
.B1(n_845),
.C1(n_840),
.Y(n_2158)
);

INVxp67_ASAP7_75t_L g2159 ( 
.A(n_2153),
.Y(n_2159)
);

HB1xp67_ASAP7_75t_L g2160 ( 
.A(n_2133),
.Y(n_2160)
);

OAI211xp5_ASAP7_75t_L g2161 ( 
.A1(n_2091),
.A2(n_2095),
.B(n_2157),
.C(n_2105),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2073),
.B(n_848),
.Y(n_2162)
);

AOI221xp5_ASAP7_75t_L g2163 ( 
.A1(n_2091),
.A2(n_2081),
.B1(n_2090),
.B2(n_2142),
.C(n_2089),
.Y(n_2163)
);

INVxp33_ASAP7_75t_L g2164 ( 
.A(n_2078),
.Y(n_2164)
);

OAI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_2107),
.A2(n_1928),
.B1(n_1877),
.B2(n_1874),
.Y(n_2165)
);

AOI21xp33_ASAP7_75t_L g2166 ( 
.A1(n_2075),
.A2(n_853),
.B(n_849),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2122),
.A2(n_1877),
.B1(n_1874),
.B2(n_1825),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_2136),
.B(n_2141),
.Y(n_2168)
);

OAI21xp33_ASAP7_75t_L g2169 ( 
.A1(n_2115),
.A2(n_1892),
.B(n_1836),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2109),
.B(n_853),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2120),
.B(n_2118),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2119),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2125),
.B(n_1874),
.Y(n_2173)
);

NOR2x1_ASAP7_75t_L g2174 ( 
.A(n_2132),
.B(n_856),
.Y(n_2174)
);

OAI221xp5_ASAP7_75t_L g2175 ( 
.A1(n_2092),
.A2(n_865),
.B1(n_867),
.B2(n_864),
.C(n_859),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2079),
.B(n_1877),
.Y(n_2176)
);

OAI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_2145),
.A2(n_1830),
.B1(n_1793),
.B2(n_1833),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2112),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2077),
.B(n_864),
.Y(n_2179)
);

OAI221xp5_ASAP7_75t_L g2180 ( 
.A1(n_2083),
.A2(n_868),
.B1(n_881),
.B2(n_867),
.C(n_865),
.Y(n_2180)
);

OAI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2074),
.A2(n_1830),
.B1(n_1793),
.B2(n_1833),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2138),
.Y(n_2182)
);

OAI21xp33_ASAP7_75t_L g2183 ( 
.A1(n_2084),
.A2(n_881),
.B(n_868),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_2076),
.Y(n_2184)
);

AOI21xp33_ASAP7_75t_L g2185 ( 
.A1(n_2151),
.A2(n_2152),
.B(n_2135),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_SL g2186 ( 
.A(n_2106),
.B(n_1706),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2130),
.B(n_883),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_2156),
.B(n_1802),
.Y(n_2188)
);

AOI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_2082),
.A2(n_1802),
.B1(n_1836),
.B2(n_1833),
.Y(n_2189)
);

INVxp67_ASAP7_75t_SL g2190 ( 
.A(n_2155),
.Y(n_2190)
);

INVx1_ASAP7_75t_SL g2191 ( 
.A(n_2085),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2103),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2093),
.B(n_1836),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2101),
.B(n_883),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2134),
.B(n_891),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_2111),
.B(n_891),
.Y(n_2196)
);

O2A1O1Ixp33_ASAP7_75t_SL g2197 ( 
.A1(n_2086),
.A2(n_2100),
.B(n_2088),
.C(n_2127),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2144),
.B(n_895),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2082),
.Y(n_2199)
);

AOI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_2080),
.A2(n_1802),
.B1(n_895),
.B2(n_898),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2137),
.Y(n_2201)
);

OR2x2_ASAP7_75t_L g2202 ( 
.A(n_2104),
.B(n_897),
.Y(n_2202)
);

OAI221xp5_ASAP7_75t_L g2203 ( 
.A1(n_2116),
.A2(n_898),
.B1(n_902),
.B2(n_900),
.C(n_897),
.Y(n_2203)
);

OAI21xp5_ASAP7_75t_L g2204 ( 
.A1(n_2158),
.A2(n_902),
.B(n_900),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2087),
.B(n_905),
.Y(n_2205)
);

AOI32xp33_ASAP7_75t_L g2206 ( 
.A1(n_2097),
.A2(n_910),
.A3(n_920),
.B1(n_913),
.B2(n_905),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2143),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2139),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2148),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2072),
.B(n_910),
.Y(n_2210)
);

AOI21xp33_ASAP7_75t_L g2211 ( 
.A1(n_2097),
.A2(n_920),
.B(n_913),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2117),
.B(n_932),
.Y(n_2212)
);

AOI21xp5_ASAP7_75t_L g2213 ( 
.A1(n_2096),
.A2(n_934),
.B(n_932),
.Y(n_2213)
);

OAI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_2098),
.A2(n_2094),
.B(n_2150),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2131),
.Y(n_2215)
);

AOI21xp5_ASAP7_75t_L g2216 ( 
.A1(n_2146),
.A2(n_935),
.B(n_934),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2121),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2147),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2114),
.Y(n_2219)
);

NAND2x1_ASAP7_75t_L g2220 ( 
.A(n_2154),
.B(n_2123),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2114),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2110),
.B(n_935),
.Y(n_2222)
);

NAND3xp33_ASAP7_75t_L g2223 ( 
.A(n_2094),
.B(n_940),
.C(n_937),
.Y(n_2223)
);

AOI221xp5_ASAP7_75t_L g2224 ( 
.A1(n_2140),
.A2(n_956),
.B1(n_958),
.B2(n_940),
.C(n_937),
.Y(n_2224)
);

INVx1_ASAP7_75t_SL g2225 ( 
.A(n_2126),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2149),
.B(n_956),
.Y(n_2226)
);

NAND2xp33_ASAP7_75t_SL g2227 ( 
.A(n_2108),
.B(n_647),
.Y(n_2227)
);

AOI21xp5_ASAP7_75t_L g2228 ( 
.A1(n_2098),
.A2(n_967),
.B(n_958),
.Y(n_2228)
);

NAND3xp33_ASAP7_75t_L g2229 ( 
.A(n_2149),
.B(n_2113),
.C(n_2128),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_2099),
.A2(n_1802),
.B1(n_888),
.B2(n_960),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2129),
.Y(n_2231)
);

NAND2xp33_ASAP7_75t_SL g2232 ( 
.A(n_2154),
.B(n_649),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2102),
.Y(n_2233)
);

AO221x1_ASAP7_75t_L g2234 ( 
.A1(n_2124),
.A2(n_1802),
.B1(n_974),
.B2(n_975),
.C(n_973),
.Y(n_2234)
);

AO22x1_ASAP7_75t_L g2235 ( 
.A1(n_2133),
.A2(n_672),
.B1(n_688),
.B2(n_651),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2133),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2133),
.Y(n_2237)
);

INVx1_ASAP7_75t_SL g2238 ( 
.A(n_2157),
.Y(n_2238)
);

OAI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_2073),
.A2(n_1802),
.B1(n_1828),
.B2(n_1820),
.Y(n_2239)
);

AOI21xp33_ASAP7_75t_SL g2240 ( 
.A1(n_2073),
.A2(n_973),
.B(n_967),
.Y(n_2240)
);

AOI32xp33_ASAP7_75t_L g2241 ( 
.A1(n_2157),
.A2(n_987),
.A3(n_1002),
.B1(n_975),
.B2(n_974),
.Y(n_2241)
);

OA21x2_ASAP7_75t_L g2242 ( 
.A1(n_2095),
.A2(n_1002),
.B(n_987),
.Y(n_2242)
);

NOR2xp33_ASAP7_75t_L g2243 ( 
.A(n_2073),
.B(n_1006),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2119),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2133),
.Y(n_2245)
);

AOI222xp33_ASAP7_75t_L g2246 ( 
.A1(n_2091),
.A2(n_1007),
.B1(n_1009),
.B2(n_1006),
.C1(n_990),
.C2(n_904),
.Y(n_2246)
);

OAI221xp5_ASAP7_75t_SL g2247 ( 
.A1(n_2091),
.A2(n_1009),
.B1(n_922),
.B2(n_928),
.C(n_923),
.Y(n_2247)
);

OAI221xp5_ASAP7_75t_L g2248 ( 
.A1(n_2091),
.A2(n_928),
.B1(n_941),
.B2(n_923),
.C(n_871),
.Y(n_2248)
);

INVx1_ASAP7_75t_SL g2249 ( 
.A(n_2157),
.Y(n_2249)
);

OAI21xp5_ASAP7_75t_L g2250 ( 
.A1(n_2095),
.A2(n_977),
.B(n_941),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2133),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2109),
.B(n_1805),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_2073),
.B(n_642),
.Y(n_2253)
);

OAI21xp33_ASAP7_75t_SL g2254 ( 
.A1(n_2115),
.A2(n_1819),
.B(n_1826),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2133),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2133),
.Y(n_2256)
);

AOI211xp5_ASAP7_75t_L g2257 ( 
.A1(n_2091),
.A2(n_1003),
.B(n_1011),
.C(n_977),
.Y(n_2257)
);

O2A1O1Ixp33_ASAP7_75t_SL g2258 ( 
.A1(n_2133),
.A2(n_1011),
.B(n_1003),
.C(n_1775),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2133),
.Y(n_2259)
);

OAI32xp33_ASAP7_75t_L g2260 ( 
.A1(n_2073),
.A2(n_1820),
.A3(n_1835),
.B1(n_1829),
.B2(n_1828),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2133),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2133),
.Y(n_2262)
);

AOI31xp33_ASAP7_75t_L g2263 ( 
.A1(n_2157),
.A2(n_644),
.A3(n_646),
.B(n_643),
.Y(n_2263)
);

INVx2_ASAP7_75t_SL g2264 ( 
.A(n_2119),
.Y(n_2264)
);

O2A1O1Ixp33_ASAP7_75t_L g2265 ( 
.A1(n_2158),
.A2(n_960),
.B(n_978),
.C(n_904),
.Y(n_2265)
);

OAI21xp33_ASAP7_75t_L g2266 ( 
.A1(n_2091),
.A2(n_656),
.B(n_653),
.Y(n_2266)
);

OAI22xp33_ASAP7_75t_L g2267 ( 
.A1(n_2073),
.A2(n_1802),
.B1(n_1828),
.B2(n_1820),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2073),
.B(n_662),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_2073),
.B(n_1802),
.Y(n_2269)
);

OAI21xp33_ASAP7_75t_L g2270 ( 
.A1(n_2091),
.A2(n_667),
.B(n_666),
.Y(n_2270)
);

AOI222xp33_ASAP7_75t_L g2271 ( 
.A1(n_2091),
.A2(n_990),
.B1(n_960),
.B2(n_1004),
.C1(n_978),
.C2(n_904),
.Y(n_2271)
);

OAI22xp33_ASAP7_75t_L g2272 ( 
.A1(n_2073),
.A2(n_1802),
.B1(n_1828),
.B2(n_1820),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2133),
.Y(n_2273)
);

AOI222xp33_ASAP7_75t_L g2274 ( 
.A1(n_2091),
.A2(n_990),
.B1(n_960),
.B2(n_1004),
.C1(n_978),
.C2(n_904),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2109),
.B(n_1805),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2133),
.Y(n_2276)
);

INVxp67_ASAP7_75t_L g2277 ( 
.A(n_2153),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2109),
.B(n_1805),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2109),
.B(n_1806),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2109),
.B(n_1806),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2133),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2073),
.B(n_671),
.Y(n_2282)
);

AOI221xp5_ASAP7_75t_SL g2283 ( 
.A1(n_2091),
.A2(n_768),
.B1(n_804),
.B2(n_693),
.C(n_660),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2073),
.B(n_675),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2073),
.B(n_676),
.Y(n_2285)
);

NOR2xp67_ASAP7_75t_SL g2286 ( 
.A(n_2073),
.B(n_677),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2133),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2109),
.B(n_1806),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2133),
.Y(n_2289)
);

OAI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2095),
.A2(n_682),
.B(n_680),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2133),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_SL g2292 ( 
.A(n_2073),
.B(n_1706),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2133),
.Y(n_2293)
);

OAI21xp33_ASAP7_75t_L g2294 ( 
.A1(n_2091),
.A2(n_687),
.B(n_683),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2073),
.B(n_691),
.Y(n_2295)
);

O2A1O1Ixp33_ASAP7_75t_SL g2296 ( 
.A1(n_2133),
.A2(n_990),
.B(n_1004),
.C(n_978),
.Y(n_2296)
);

OAI21xp33_ASAP7_75t_L g2297 ( 
.A1(n_2091),
.A2(n_695),
.B(n_694),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2073),
.A2(n_1004),
.B1(n_1808),
.B2(n_1829),
.Y(n_2298)
);

INVxp67_ASAP7_75t_SL g2299 ( 
.A(n_2133),
.Y(n_2299)
);

OAI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2073),
.A2(n_1849),
.B1(n_1794),
.B2(n_1835),
.Y(n_2300)
);

INVx2_ASAP7_75t_SL g2301 ( 
.A(n_2119),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2133),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2133),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2109),
.B(n_1787),
.Y(n_2304)
);

INVx1_ASAP7_75t_SL g2305 ( 
.A(n_2157),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2133),
.Y(n_2306)
);

OAI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_2073),
.A2(n_1794),
.B1(n_1835),
.B2(n_1829),
.Y(n_2307)
);

NAND3xp33_ASAP7_75t_L g2308 ( 
.A(n_2095),
.B(n_693),
.C(n_660),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2220),
.Y(n_2309)
);

OAI21xp33_ASAP7_75t_SL g2310 ( 
.A1(n_2299),
.A2(n_1866),
.B(n_1826),
.Y(n_2310)
);

NOR4xp25_ASAP7_75t_L g2311 ( 
.A(n_2161),
.B(n_3),
.C(n_1),
.D(n_2),
.Y(n_2311)
);

OAI21xp33_ASAP7_75t_L g2312 ( 
.A1(n_2164),
.A2(n_1815),
.B(n_1784),
.Y(n_2312)
);

AOI22xp33_ASAP7_75t_L g2313 ( 
.A1(n_2238),
.A2(n_1815),
.B1(n_693),
.B2(n_768),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_L g2314 ( 
.A(n_2249),
.B(n_700),
.Y(n_2314)
);

OAI21xp33_ASAP7_75t_L g2315 ( 
.A1(n_2305),
.A2(n_1815),
.B(n_1784),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2160),
.Y(n_2316)
);

INVxp33_ASAP7_75t_L g2317 ( 
.A(n_2286),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2264),
.Y(n_2318)
);

AOI221xp5_ASAP7_75t_L g2319 ( 
.A1(n_2197),
.A2(n_702),
.B1(n_713),
.B2(n_707),
.C(n_706),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2301),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2184),
.Y(n_2321)
);

AOI32xp33_ASAP7_75t_L g2322 ( 
.A1(n_2182),
.A2(n_751),
.A3(n_767),
.B1(n_733),
.B2(n_718),
.Y(n_2322)
);

AOI211xp5_ASAP7_75t_L g2323 ( 
.A1(n_2168),
.A2(n_739),
.B(n_755),
.C(n_721),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2184),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2263),
.B(n_714),
.Y(n_2325)
);

NAND4xp25_ASAP7_75t_SL g2326 ( 
.A(n_2163),
.B(n_1815),
.C(n_1787),
.D(n_1827),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2190),
.B(n_715),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2244),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2236),
.Y(n_2329)
);

NAND3xp33_ASAP7_75t_L g2330 ( 
.A(n_2292),
.B(n_722),
.C(n_717),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2171),
.Y(n_2331)
);

AOI21xp33_ASAP7_75t_SL g2332 ( 
.A1(n_2253),
.A2(n_2),
.B(n_3),
.Y(n_2332)
);

AOI21xp33_ASAP7_75t_L g2333 ( 
.A1(n_2243),
.A2(n_725),
.B(n_723),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2172),
.B(n_728),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2159),
.B(n_730),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2277),
.B(n_732),
.Y(n_2336)
);

NAND3xp33_ASAP7_75t_SL g2337 ( 
.A(n_2271),
.B(n_741),
.C(n_737),
.Y(n_2337)
);

INVx1_ASAP7_75t_SL g2338 ( 
.A(n_2191),
.Y(n_2338)
);

AOI221xp5_ASAP7_75t_L g2339 ( 
.A1(n_2195),
.A2(n_2214),
.B1(n_2247),
.B2(n_2245),
.C(n_2237),
.Y(n_2339)
);

OAI21xp5_ASAP7_75t_L g2340 ( 
.A1(n_2209),
.A2(n_777),
.B(n_753),
.Y(n_2340)
);

AOI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2233),
.A2(n_744),
.B1(n_745),
.B2(n_742),
.Y(n_2341)
);

AND2x4_ASAP7_75t_L g2342 ( 
.A(n_2251),
.B(n_1809),
.Y(n_2342)
);

OAI221xp5_ASAP7_75t_L g2343 ( 
.A1(n_2225),
.A2(n_746),
.B1(n_760),
.B2(n_758),
.C(n_752),
.Y(n_2343)
);

OAI32xp33_ASAP7_75t_L g2344 ( 
.A1(n_2254),
.A2(n_1814),
.A3(n_1811),
.B1(n_1796),
.B2(n_772),
.Y(n_2344)
);

AOI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2186),
.A2(n_763),
.B1(n_775),
.B2(n_761),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2255),
.Y(n_2346)
);

INVxp67_ASAP7_75t_L g2347 ( 
.A(n_2174),
.Y(n_2347)
);

OAI322xp33_ASAP7_75t_L g2348 ( 
.A1(n_2256),
.A2(n_778),
.A3(n_786),
.B1(n_780),
.B2(n_790),
.C1(n_788),
.C2(n_783),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2259),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2261),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2219),
.A2(n_794),
.B1(n_796),
.B2(n_793),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2262),
.B(n_800),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2273),
.Y(n_2353)
);

OAI221xp5_ASAP7_75t_L g2354 ( 
.A1(n_2266),
.A2(n_807),
.B1(n_808),
.B2(n_806),
.C(n_802),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2199),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2276),
.Y(n_2356)
);

AOI221xp5_ASAP7_75t_SL g2357 ( 
.A1(n_2281),
.A2(n_768),
.B1(n_804),
.B2(n_693),
.C(n_660),
.Y(n_2357)
);

OAI31xp33_ASAP7_75t_L g2358 ( 
.A1(n_2232),
.A2(n_1811),
.A3(n_1702),
.B(n_1827),
.Y(n_2358)
);

AOI221xp5_ASAP7_75t_L g2359 ( 
.A1(n_2287),
.A2(n_2289),
.B1(n_2302),
.B2(n_2293),
.C(n_2291),
.Y(n_2359)
);

NOR4xp25_ASAP7_75t_L g2360 ( 
.A(n_2303),
.B(n_7),
.C(n_4),
.D(n_6),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2306),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2242),
.Y(n_2362)
);

OR2x2_ASAP7_75t_L g2363 ( 
.A(n_2207),
.B(n_4),
.Y(n_2363)
);

OAI21xp33_ASAP7_75t_L g2364 ( 
.A1(n_2169),
.A2(n_810),
.B(n_809),
.Y(n_2364)
);

OAI21xp5_ASAP7_75t_L g2365 ( 
.A1(n_2229),
.A2(n_851),
.B(n_825),
.Y(n_2365)
);

OAI221xp5_ASAP7_75t_L g2366 ( 
.A1(n_2266),
.A2(n_2297),
.B1(n_2294),
.B2(n_2270),
.C(n_2200),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2242),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2221),
.B(n_1787),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2178),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2252),
.A2(n_815),
.B1(n_817),
.B2(n_814),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2192),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2275),
.Y(n_2372)
);

INVxp67_ASAP7_75t_SL g2373 ( 
.A(n_2268),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2194),
.B(n_819),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2201),
.Y(n_2375)
);

AOI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2278),
.A2(n_827),
.B1(n_830),
.B2(n_820),
.Y(n_2376)
);

OAI22xp33_ASAP7_75t_L g2377 ( 
.A1(n_2282),
.A2(n_1818),
.B1(n_1796),
.B2(n_1785),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2215),
.B(n_833),
.Y(n_2378)
);

OAI221xp5_ASAP7_75t_SL g2379 ( 
.A1(n_2206),
.A2(n_2175),
.B1(n_2241),
.B2(n_2208),
.C(n_2246),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2170),
.Y(n_2380)
);

AOI21xp33_ASAP7_75t_L g2381 ( 
.A1(n_2274),
.A2(n_842),
.B(n_839),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_2296),
.A2(n_882),
.B(n_861),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2222),
.Y(n_2383)
);

A2O1A1Ixp33_ASAP7_75t_L g2384 ( 
.A1(n_2270),
.A2(n_847),
.B(n_854),
.C(n_846),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2196),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2162),
.Y(n_2386)
);

OAI221xp5_ASAP7_75t_L g2387 ( 
.A1(n_2294),
.A2(n_862),
.B1(n_863),
.B2(n_860),
.C(n_858),
.Y(n_2387)
);

AOI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_2297),
.A2(n_870),
.B1(n_873),
.B2(n_869),
.Y(n_2388)
);

AOI22xp33_ASAP7_75t_L g2389 ( 
.A1(n_2304),
.A2(n_768),
.B1(n_804),
.B2(n_660),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2187),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2179),
.Y(n_2391)
);

OAI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_2284),
.A2(n_1818),
.B1(n_1791),
.B2(n_1792),
.Y(n_2392)
);

AOI21xp33_ASAP7_75t_L g2393 ( 
.A1(n_2285),
.A2(n_879),
.B(n_876),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2295),
.B(n_884),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2173),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2212),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_2218),
.B(n_2185),
.Y(n_2397)
);

AOI21xp33_ASAP7_75t_SL g2398 ( 
.A1(n_2235),
.A2(n_6),
.B(n_8),
.Y(n_2398)
);

OAI221xp5_ASAP7_75t_L g2399 ( 
.A1(n_2230),
.A2(n_887),
.B1(n_889),
.B2(n_886),
.C(n_885),
.Y(n_2399)
);

AO221x1_ASAP7_75t_L g2400 ( 
.A1(n_2240),
.A2(n_768),
.B1(n_804),
.B2(n_693),
.C(n_660),
.Y(n_2400)
);

INVx1_ASAP7_75t_SL g2401 ( 
.A(n_2227),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2202),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2193),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2231),
.B(n_890),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2217),
.B(n_2290),
.Y(n_2405)
);

OAI32xp33_ASAP7_75t_L g2406 ( 
.A1(n_2269),
.A2(n_896),
.A3(n_899),
.B1(n_893),
.B2(n_892),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2250),
.B(n_2176),
.Y(n_2407)
);

OR2x2_ASAP7_75t_L g2408 ( 
.A(n_2205),
.B(n_9),
.Y(n_2408)
);

OR4x1_ASAP7_75t_L g2409 ( 
.A(n_2234),
.B(n_1058),
.C(n_1818),
.D(n_1791),
.Y(n_2409)
);

AOI322xp5_ASAP7_75t_L g2410 ( 
.A1(n_2283),
.A2(n_901),
.A3(n_907),
.B1(n_903),
.B2(n_914),
.C1(n_908),
.C2(n_906),
.Y(n_2410)
);

NOR2x1_ASAP7_75t_L g2411 ( 
.A(n_2308),
.B(n_693),
.Y(n_2411)
);

OAI31xp33_ASAP7_75t_L g2412 ( 
.A1(n_2165),
.A2(n_1827),
.A3(n_1728),
.B(n_14),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_2198),
.B(n_918),
.Y(n_2413)
);

OAI21xp5_ASAP7_75t_L g2414 ( 
.A1(n_2298),
.A2(n_948),
.B(n_927),
.Y(n_2414)
);

INVxp67_ASAP7_75t_L g2415 ( 
.A(n_2210),
.Y(n_2415)
);

NOR2xp33_ASAP7_75t_L g2416 ( 
.A(n_2183),
.B(n_925),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_2279),
.B(n_1809),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2226),
.Y(n_2418)
);

NAND3xp33_ASAP7_75t_SL g2419 ( 
.A(n_2257),
.B(n_929),
.C(n_926),
.Y(n_2419)
);

AOI221xp5_ASAP7_75t_L g2420 ( 
.A1(n_2248),
.A2(n_942),
.B1(n_944),
.B2(n_939),
.C(n_933),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2183),
.B(n_946),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2216),
.B(n_949),
.Y(n_2422)
);

OAI22xp33_ASAP7_75t_L g2423 ( 
.A1(n_2189),
.A2(n_1785),
.B1(n_1795),
.B2(n_1783),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2223),
.Y(n_2424)
);

AOI22xp33_ASAP7_75t_L g2425 ( 
.A1(n_2280),
.A2(n_804),
.B1(n_919),
.B2(n_768),
.Y(n_2425)
);

OAI21xp33_ASAP7_75t_L g2426 ( 
.A1(n_2288),
.A2(n_952),
.B(n_951),
.Y(n_2426)
);

AOI221xp5_ASAP7_75t_L g2427 ( 
.A1(n_2166),
.A2(n_959),
.B1(n_963),
.B2(n_955),
.C(n_954),
.Y(n_2427)
);

AOI21xp5_ASAP7_75t_L g2428 ( 
.A1(n_2317),
.A2(n_2258),
.B(n_2180),
.Y(n_2428)
);

OAI221xp5_ASAP7_75t_L g2429 ( 
.A1(n_2311),
.A2(n_2224),
.B1(n_2203),
.B2(n_2177),
.C(n_2211),
.Y(n_2429)
);

AOI211xp5_ASAP7_75t_SL g2430 ( 
.A1(n_2347),
.A2(n_2267),
.B(n_2272),
.C(n_2239),
.Y(n_2430)
);

OAI211xp5_ASAP7_75t_SL g2431 ( 
.A1(n_2339),
.A2(n_2265),
.B(n_2204),
.C(n_2228),
.Y(n_2431)
);

HB1xp67_ASAP7_75t_L g2432 ( 
.A(n_2309),
.Y(n_2432)
);

NOR2x1_ASAP7_75t_L g2433 ( 
.A(n_2316),
.B(n_2213),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_L g2434 ( 
.A(n_2338),
.B(n_2181),
.Y(n_2434)
);

NOR3xp33_ASAP7_75t_L g2435 ( 
.A(n_2379),
.B(n_2188),
.C(n_2300),
.Y(n_2435)
);

AOI22xp33_ASAP7_75t_L g2436 ( 
.A1(n_2318),
.A2(n_2307),
.B1(n_2167),
.B2(n_919),
.Y(n_2436)
);

OAI221xp5_ASAP7_75t_SL g2437 ( 
.A1(n_2359),
.A2(n_2412),
.B1(n_2320),
.B2(n_2328),
.C(n_2358),
.Y(n_2437)
);

AOI322xp5_ASAP7_75t_L g2438 ( 
.A1(n_2397),
.A2(n_2260),
.A3(n_964),
.B1(n_965),
.B2(n_970),
.C1(n_980),
.C2(n_972),
.Y(n_2438)
);

AOI22xp33_ASAP7_75t_L g2439 ( 
.A1(n_2331),
.A2(n_919),
.B1(n_930),
.B2(n_804),
.Y(n_2439)
);

NAND2x1_ASAP7_75t_SL g2440 ( 
.A(n_2362),
.B(n_1801),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2324),
.B(n_968),
.Y(n_2441)
);

AOI21xp5_ASAP7_75t_L g2442 ( 
.A1(n_2319),
.A2(n_983),
.B(n_982),
.Y(n_2442)
);

OAI211xp5_ASAP7_75t_L g2443 ( 
.A1(n_2360),
.A2(n_985),
.B(n_986),
.C(n_984),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2321),
.Y(n_2444)
);

AOI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_2365),
.A2(n_991),
.B(n_989),
.Y(n_2445)
);

NAND4xp25_ASAP7_75t_SL g2446 ( 
.A(n_2401),
.B(n_1832),
.C(n_1785),
.D(n_1795),
.Y(n_2446)
);

OAI211xp5_ASAP7_75t_SL g2447 ( 
.A1(n_2415),
.A2(n_995),
.B(n_996),
.C(n_992),
.Y(n_2447)
);

OAI222xp33_ASAP7_75t_L g2448 ( 
.A1(n_2329),
.A2(n_1010),
.B1(n_999),
.B2(n_1012),
.C1(n_1005),
.C2(n_997),
.Y(n_2448)
);

OAI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2355),
.A2(n_1791),
.B1(n_1792),
.B2(n_1790),
.Y(n_2449)
);

AOI211x1_ASAP7_75t_L g2450 ( 
.A1(n_2366),
.A2(n_1817),
.B(n_1792),
.C(n_1790),
.Y(n_2450)
);

OAI221xp5_ASAP7_75t_SL g2451 ( 
.A1(n_2341),
.A2(n_1712),
.B1(n_1832),
.B2(n_1724),
.C(n_1785),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2346),
.B(n_1013),
.Y(n_2452)
);

OA21x2_ASAP7_75t_L g2453 ( 
.A1(n_2367),
.A2(n_1014),
.B(n_1866),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2363),
.Y(n_2454)
);

AOI22xp5_ASAP7_75t_L g2455 ( 
.A1(n_2326),
.A2(n_930),
.B1(n_998),
.B2(n_919),
.Y(n_2455)
);

AOI322xp5_ASAP7_75t_L g2456 ( 
.A1(n_2349),
.A2(n_1783),
.A3(n_1795),
.B1(n_1798),
.B2(n_1810),
.C1(n_1807),
.C2(n_1801),
.Y(n_2456)
);

AOI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2372),
.A2(n_930),
.B1(n_998),
.B2(n_919),
.Y(n_2457)
);

NOR3xp33_ASAP7_75t_L g2458 ( 
.A(n_2337),
.B(n_1826),
.C(n_1817),
.Y(n_2458)
);

INVxp67_ASAP7_75t_L g2459 ( 
.A(n_2325),
.Y(n_2459)
);

AOI211xp5_ASAP7_75t_L g2460 ( 
.A1(n_2350),
.A2(n_930),
.B(n_998),
.C(n_919),
.Y(n_2460)
);

OAI21xp5_ASAP7_75t_SL g2461 ( 
.A1(n_2353),
.A2(n_998),
.B(n_930),
.Y(n_2461)
);

AOI21xp5_ASAP7_75t_L g2462 ( 
.A1(n_2374),
.A2(n_998),
.B(n_930),
.Y(n_2462)
);

AOI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2422),
.A2(n_2327),
.B(n_2382),
.Y(n_2463)
);

NOR3xp33_ASAP7_75t_L g2464 ( 
.A(n_2419),
.B(n_1817),
.C(n_10),
.Y(n_2464)
);

INVxp33_ASAP7_75t_SL g2465 ( 
.A(n_2314),
.Y(n_2465)
);

OAI22xp5_ASAP7_75t_L g2466 ( 
.A1(n_2356),
.A2(n_1807),
.B1(n_1810),
.B2(n_1801),
.Y(n_2466)
);

NAND2x1_ASAP7_75t_L g2467 ( 
.A(n_2403),
.B(n_998),
.Y(n_2467)
);

OAI221xp5_ASAP7_75t_L g2468 ( 
.A1(n_2361),
.A2(n_2322),
.B1(n_2345),
.B2(n_2364),
.C(n_2373),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2332),
.B(n_10),
.Y(n_2469)
);

OAI221xp5_ASAP7_75t_L g2470 ( 
.A1(n_2426),
.A2(n_1712),
.B1(n_1810),
.B2(n_1807),
.C(n_1783),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2408),
.Y(n_2471)
);

OAI211xp5_ASAP7_75t_L g2472 ( 
.A1(n_2410),
.A2(n_16),
.B(n_11),
.C(n_15),
.Y(n_2472)
);

AOI21xp33_ASAP7_75t_L g2473 ( 
.A1(n_2334),
.A2(n_15),
.B(n_16),
.Y(n_2473)
);

OAI21xp5_ASAP7_75t_L g2474 ( 
.A1(n_2330),
.A2(n_1728),
.B(n_1783),
.Y(n_2474)
);

AOI221xp5_ASAP7_75t_L g2475 ( 
.A1(n_2344),
.A2(n_2375),
.B1(n_2424),
.B2(n_2369),
.C(n_2398),
.Y(n_2475)
);

NAND3xp33_ASAP7_75t_L g2476 ( 
.A(n_2323),
.B(n_17),
.C(n_19),
.Y(n_2476)
);

OAI31xp33_ASAP7_75t_L g2477 ( 
.A1(n_2371),
.A2(n_20),
.A3(n_17),
.B(n_19),
.Y(n_2477)
);

O2A1O1Ixp33_ASAP7_75t_L g2478 ( 
.A1(n_2384),
.A2(n_23),
.B(n_20),
.C(n_21),
.Y(n_2478)
);

O2A1O1Ixp33_ASAP7_75t_L g2479 ( 
.A1(n_2381),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_2479)
);

AOI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2368),
.A2(n_1808),
.B1(n_1816),
.B2(n_1795),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2383),
.B(n_1809),
.Y(n_2481)
);

AOI221xp5_ASAP7_75t_L g2482 ( 
.A1(n_2409),
.A2(n_1808),
.B1(n_1798),
.B2(n_27),
.C(n_24),
.Y(n_2482)
);

NAND3xp33_ASAP7_75t_L g2483 ( 
.A(n_2313),
.B(n_26),
.C(n_29),
.Y(n_2483)
);

AOI21xp5_ASAP7_75t_L g2484 ( 
.A1(n_2343),
.A2(n_1808),
.B(n_1816),
.Y(n_2484)
);

NOR3x1_ASAP7_75t_L g2485 ( 
.A(n_2400),
.B(n_30),
.C(n_31),
.Y(n_2485)
);

AOI211xp5_ASAP7_75t_L g2486 ( 
.A1(n_2399),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2386),
.B(n_1809),
.Y(n_2487)
);

AOI21xp5_ASAP7_75t_L g2488 ( 
.A1(n_2404),
.A2(n_1816),
.B(n_1798),
.Y(n_2488)
);

OAI21xp5_ASAP7_75t_SL g2489 ( 
.A1(n_2405),
.A2(n_33),
.B(n_35),
.Y(n_2489)
);

NOR3xp33_ASAP7_75t_L g2490 ( 
.A(n_2418),
.B(n_35),
.C(n_36),
.Y(n_2490)
);

OAI221xp5_ASAP7_75t_L g2491 ( 
.A1(n_2395),
.A2(n_2385),
.B1(n_2340),
.B2(n_2376),
.C(n_2370),
.Y(n_2491)
);

AOI21xp5_ASAP7_75t_L g2492 ( 
.A1(n_2352),
.A2(n_1816),
.B(n_1798),
.Y(n_2492)
);

OAI221xp5_ASAP7_75t_L g2493 ( 
.A1(n_2351),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.C(n_40),
.Y(n_2493)
);

AOI21xp33_ASAP7_75t_L g2494 ( 
.A1(n_2335),
.A2(n_37),
.B(n_39),
.Y(n_2494)
);

NOR4xp25_ASAP7_75t_L g2495 ( 
.A(n_2348),
.B(n_43),
.C(n_41),
.D(n_42),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2378),
.Y(n_2496)
);

AOI21xp5_ASAP7_75t_L g2497 ( 
.A1(n_2336),
.A2(n_1816),
.B(n_1831),
.Y(n_2497)
);

AOI211xp5_ASAP7_75t_SL g2498 ( 
.A1(n_2402),
.A2(n_44),
.B(n_41),
.C(n_42),
.Y(n_2498)
);

OAI21xp33_ASAP7_75t_L g2499 ( 
.A1(n_2380),
.A2(n_1804),
.B(n_1800),
.Y(n_2499)
);

NAND3xp33_ASAP7_75t_L g2500 ( 
.A(n_2420),
.B(n_46),
.C(n_47),
.Y(n_2500)
);

OAI221xp5_ASAP7_75t_L g2501 ( 
.A1(n_2351),
.A2(n_49),
.B1(n_46),
.B2(n_48),
.C(n_50),
.Y(n_2501)
);

AOI322xp5_ASAP7_75t_L g2502 ( 
.A1(n_2391),
.A2(n_1804),
.A3(n_1800),
.B1(n_55),
.B2(n_52),
.C1(n_54),
.C2(n_50),
.Y(n_2502)
);

O2A1O1Ixp33_ASAP7_75t_L g2503 ( 
.A1(n_2414),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_2503)
);

NAND3xp33_ASAP7_75t_L g2504 ( 
.A(n_2389),
.B(n_51),
.C(n_53),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2413),
.B(n_54),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2390),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2396),
.B(n_55),
.Y(n_2507)
);

OAI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2407),
.A2(n_1789),
.B(n_56),
.Y(n_2508)
);

AOI322xp5_ASAP7_75t_L g2509 ( 
.A1(n_2411),
.A2(n_1804),
.A3(n_1800),
.B1(n_64),
.B2(n_61),
.C1(n_63),
.C2(n_59),
.Y(n_2509)
);

AOI221x1_ASAP7_75t_L g2510 ( 
.A1(n_2421),
.A2(n_63),
.B1(n_60),
.B2(n_62),
.C(n_66),
.Y(n_2510)
);

AOI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_2406),
.A2(n_1831),
.B(n_60),
.Y(n_2511)
);

AOI211xp5_ASAP7_75t_SL g2512 ( 
.A1(n_2315),
.A2(n_67),
.B(n_62),
.C(n_66),
.Y(n_2512)
);

AOI22xp33_ASAP7_75t_SL g2513 ( 
.A1(n_2342),
.A2(n_1831),
.B1(n_1800),
.B2(n_1804),
.Y(n_2513)
);

AOI221xp5_ASAP7_75t_L g2514 ( 
.A1(n_2357),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.C(n_70),
.Y(n_2514)
);

AO21x1_ASAP7_75t_L g2515 ( 
.A1(n_2342),
.A2(n_70),
.B(n_71),
.Y(n_2515)
);

OAI21xp33_ASAP7_75t_L g2516 ( 
.A1(n_2425),
.A2(n_1789),
.B(n_71),
.Y(n_2516)
);

AO22x2_ASAP7_75t_L g2517 ( 
.A1(n_2392),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_2517)
);

AOI211xp5_ASAP7_75t_L g2518 ( 
.A1(n_2427),
.A2(n_75),
.B(n_72),
.C(n_73),
.Y(n_2518)
);

AOI321xp33_ASAP7_75t_L g2519 ( 
.A1(n_2312),
.A2(n_78),
.A3(n_80),
.B1(n_76),
.B2(n_77),
.C(n_79),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2394),
.Y(n_2520)
);

AOI21xp33_ASAP7_75t_SL g2521 ( 
.A1(n_2416),
.A2(n_76),
.B(n_78),
.Y(n_2521)
);

AOI21x1_ASAP7_75t_L g2522 ( 
.A1(n_2417),
.A2(n_2333),
.B(n_2393),
.Y(n_2522)
);

AOI221xp5_ASAP7_75t_L g2523 ( 
.A1(n_2377),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.C(n_82),
.Y(n_2523)
);

AOI21xp33_ASAP7_75t_L g2524 ( 
.A1(n_2388),
.A2(n_83),
.B(n_84),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2354),
.A2(n_1831),
.B(n_84),
.Y(n_2525)
);

NOR3xp33_ASAP7_75t_L g2526 ( 
.A(n_2387),
.B(n_85),
.C(n_86),
.Y(n_2526)
);

O2A1O1Ixp33_ASAP7_75t_L g2527 ( 
.A1(n_2310),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_2527)
);

NOR3xp33_ASAP7_75t_L g2528 ( 
.A(n_2388),
.B(n_88),
.C(n_89),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2417),
.B(n_2423),
.Y(n_2529)
);

AOI22xp33_ASAP7_75t_SL g2530 ( 
.A1(n_2310),
.A2(n_1831),
.B1(n_1721),
.B2(n_1747),
.Y(n_2530)
);

INVx2_ASAP7_75t_SL g2531 ( 
.A(n_2324),
.Y(n_2531)
);

OAI211xp5_ASAP7_75t_SL g2532 ( 
.A1(n_2339),
.A2(n_91),
.B(n_88),
.C(n_89),
.Y(n_2532)
);

OAI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2338),
.A2(n_1721),
.B1(n_1756),
.B2(n_1680),
.Y(n_2533)
);

NAND3xp33_ASAP7_75t_L g2534 ( 
.A(n_2359),
.B(n_92),
.C(n_93),
.Y(n_2534)
);

OAI222xp33_ASAP7_75t_L g2535 ( 
.A1(n_2338),
.A2(n_96),
.B1(n_98),
.B2(n_94),
.C1(n_95),
.C2(n_97),
.Y(n_2535)
);

AOI321xp33_ASAP7_75t_L g2536 ( 
.A1(n_2359),
.A2(n_100),
.A3(n_102),
.B1(n_94),
.B2(n_99),
.C(n_101),
.Y(n_2536)
);

OA22x2_ASAP7_75t_L g2537 ( 
.A1(n_2309),
.A2(n_104),
.B1(n_101),
.B2(n_102),
.Y(n_2537)
);

AOI21xp5_ASAP7_75t_L g2538 ( 
.A1(n_2317),
.A2(n_104),
.B(n_105),
.Y(n_2538)
);

NOR3xp33_ASAP7_75t_L g2539 ( 
.A(n_2379),
.B(n_107),
.C(n_108),
.Y(n_2539)
);

NOR2x1_ASAP7_75t_L g2540 ( 
.A(n_2309),
.B(n_109),
.Y(n_2540)
);

AOI21xp5_ASAP7_75t_L g2541 ( 
.A1(n_2317),
.A2(n_110),
.B(n_111),
.Y(n_2541)
);

OAI21xp33_ASAP7_75t_L g2542 ( 
.A1(n_2338),
.A2(n_1789),
.B(n_110),
.Y(n_2542)
);

O2A1O1Ixp33_ASAP7_75t_L g2543 ( 
.A1(n_2311),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_2543)
);

OAI322xp33_ASAP7_75t_L g2544 ( 
.A1(n_2338),
.A2(n_117),
.A3(n_116),
.B1(n_114),
.B2(n_112),
.C1(n_113),
.C2(n_115),
.Y(n_2544)
);

OAI21xp33_ASAP7_75t_SL g2545 ( 
.A1(n_2362),
.A2(n_1789),
.B(n_115),
.Y(n_2545)
);

AOI21xp33_ASAP7_75t_SL g2546 ( 
.A1(n_2347),
.A2(n_117),
.B(n_119),
.Y(n_2546)
);

AOI221xp5_ASAP7_75t_L g2547 ( 
.A1(n_2311),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.C(n_123),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2338),
.B(n_120),
.Y(n_2548)
);

OAI221xp5_ASAP7_75t_L g2549 ( 
.A1(n_2311),
.A2(n_124),
.B1(n_121),
.B2(n_122),
.C(n_125),
.Y(n_2549)
);

AOI22xp5_ASAP7_75t_L g2550 ( 
.A1(n_2338),
.A2(n_1747),
.B1(n_1756),
.B2(n_127),
.Y(n_2550)
);

AOI21xp33_ASAP7_75t_L g2551 ( 
.A1(n_2317),
.A2(n_124),
.B(n_126),
.Y(n_2551)
);

OAI21xp33_ASAP7_75t_SL g2552 ( 
.A1(n_2362),
.A2(n_126),
.B(n_127),
.Y(n_2552)
);

XNOR2xp5_ASAP7_75t_L g2553 ( 
.A(n_2338),
.B(n_128),
.Y(n_2553)
);

AOI22xp33_ASAP7_75t_L g2554 ( 
.A1(n_2318),
.A2(n_1747),
.B1(n_1756),
.B2(n_131),
.Y(n_2554)
);

NOR3xp33_ASAP7_75t_L g2555 ( 
.A(n_2379),
.B(n_129),
.C(n_130),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2318),
.Y(n_2556)
);

AOI211xp5_ASAP7_75t_SL g2557 ( 
.A1(n_2347),
.A2(n_136),
.B(n_132),
.C(n_134),
.Y(n_2557)
);

OAI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2311),
.A2(n_132),
.B(n_136),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2318),
.B(n_137),
.Y(n_2559)
);

AOI221xp5_ASAP7_75t_L g2560 ( 
.A1(n_2311),
.A2(n_141),
.B1(n_137),
.B2(n_138),
.C(n_142),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_L g2561 ( 
.A(n_2317),
.B(n_143),
.Y(n_2561)
);

AOI221xp5_ASAP7_75t_L g2562 ( 
.A1(n_2311),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.C(n_148),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2338),
.B(n_147),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_2317),
.B(n_149),
.Y(n_2564)
);

OAI221xp5_ASAP7_75t_L g2565 ( 
.A1(n_2311),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.C(n_152),
.Y(n_2565)
);

AOI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2338),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_2566)
);

OAI21xp33_ASAP7_75t_L g2567 ( 
.A1(n_2338),
.A2(n_153),
.B(n_154),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2338),
.B(n_154),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2338),
.B(n_155),
.Y(n_2569)
);

OAI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2311),
.A2(n_155),
.B(n_156),
.Y(n_2570)
);

AOI21xp5_ASAP7_75t_L g2571 ( 
.A1(n_2317),
.A2(n_156),
.B(n_157),
.Y(n_2571)
);

OAI221xp5_ASAP7_75t_L g2572 ( 
.A1(n_2311),
.A2(n_162),
.B1(n_159),
.B2(n_161),
.C(n_163),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2318),
.Y(n_2573)
);

NAND4xp25_ASAP7_75t_L g2574 ( 
.A(n_2359),
.B(n_163),
.C(n_161),
.D(n_162),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2318),
.B(n_164),
.Y(n_2575)
);

OAI22xp33_ASAP7_75t_L g2576 ( 
.A1(n_2338),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2540),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2432),
.Y(n_2578)
);

OAI211xp5_ASAP7_75t_SL g2579 ( 
.A1(n_2475),
.A2(n_167),
.B(n_165),
.C(n_166),
.Y(n_2579)
);

INVxp67_ASAP7_75t_L g2580 ( 
.A(n_2469),
.Y(n_2580)
);

O2A1O1Ixp33_ASAP7_75t_L g2581 ( 
.A1(n_2543),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_2581)
);

OAI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2534),
.A2(n_168),
.B(n_169),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2515),
.Y(n_2583)
);

AOI221xp5_ASAP7_75t_L g2584 ( 
.A1(n_2539),
.A2(n_173),
.B1(n_170),
.B2(n_171),
.C(n_174),
.Y(n_2584)
);

BUFx2_ASAP7_75t_L g2585 ( 
.A(n_2552),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2536),
.B(n_171),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2498),
.B(n_2557),
.Y(n_2587)
);

AOI221xp5_ASAP7_75t_L g2588 ( 
.A1(n_2555),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.C(n_177),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_SL g2589 ( 
.A(n_2535),
.B(n_176),
.Y(n_2589)
);

OAI21xp5_ASAP7_75t_SL g2590 ( 
.A1(n_2434),
.A2(n_178),
.B(n_179),
.Y(n_2590)
);

AOI22xp33_ASAP7_75t_L g2591 ( 
.A1(n_2435),
.A2(n_2532),
.B1(n_2573),
.B2(n_2556),
.Y(n_2591)
);

AOI221xp5_ASAP7_75t_L g2592 ( 
.A1(n_2495),
.A2(n_183),
.B1(n_179),
.B2(n_181),
.C(n_184),
.Y(n_2592)
);

A2O1A1Ixp33_ASAP7_75t_L g2593 ( 
.A1(n_2547),
.A2(n_187),
.B(n_184),
.C(n_186),
.Y(n_2593)
);

AOI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2531),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_2594)
);

INVxp67_ASAP7_75t_L g2595 ( 
.A(n_2561),
.Y(n_2595)
);

OAI22xp33_ASAP7_75t_SL g2596 ( 
.A1(n_2437),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2559),
.B(n_189),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2440),
.Y(n_2598)
);

AOI221xp5_ASAP7_75t_L g2599 ( 
.A1(n_2558),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.C(n_194),
.Y(n_2599)
);

NAND4xp25_ASAP7_75t_L g2600 ( 
.A(n_2428),
.B(n_197),
.C(n_195),
.D(n_196),
.Y(n_2600)
);

OAI22xp5_ASAP7_75t_L g2601 ( 
.A1(n_2549),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_2601)
);

AOI221x1_ASAP7_75t_L g2602 ( 
.A1(n_2574),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.C(n_202),
.Y(n_2602)
);

AOI21xp5_ASAP7_75t_L g2603 ( 
.A1(n_2565),
.A2(n_200),
.B(n_201),
.Y(n_2603)
);

OAI22xp5_ASAP7_75t_L g2604 ( 
.A1(n_2572),
.A2(n_205),
.B1(n_202),
.B2(n_204),
.Y(n_2604)
);

A2O1A1Ixp33_ASAP7_75t_L g2605 ( 
.A1(n_2560),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_2605)
);

OAI21xp33_ASAP7_75t_L g2606 ( 
.A1(n_2465),
.A2(n_206),
.B(n_207),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2553),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_SL g2608 ( 
.A(n_2477),
.B(n_208),
.Y(n_2608)
);

OAI222xp33_ASAP7_75t_L g2609 ( 
.A1(n_2429),
.A2(n_211),
.B1(n_217),
.B2(n_209),
.C1(n_210),
.C2(n_216),
.Y(n_2609)
);

AOI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2564),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2610)
);

OAI211xp5_ASAP7_75t_L g2611 ( 
.A1(n_2570),
.A2(n_219),
.B(n_216),
.C(n_218),
.Y(n_2611)
);

OA21x2_ASAP7_75t_L g2612 ( 
.A1(n_2548),
.A2(n_218),
.B(n_222),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2454),
.Y(n_2613)
);

OAI21xp5_ASAP7_75t_SL g2614 ( 
.A1(n_2431),
.A2(n_2512),
.B(n_2443),
.Y(n_2614)
);

AOI22xp33_ASAP7_75t_L g2615 ( 
.A1(n_2464),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_2615)
);

AOI22xp33_ASAP7_75t_L g2616 ( 
.A1(n_2471),
.A2(n_228),
.B1(n_224),
.B2(n_225),
.Y(n_2616)
);

AOI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2527),
.A2(n_225),
.B(n_228),
.Y(n_2617)
);

AOI221xp5_ASAP7_75t_L g2618 ( 
.A1(n_2562),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.C(n_232),
.Y(n_2618)
);

O2A1O1Ixp33_ASAP7_75t_L g2619 ( 
.A1(n_2546),
.A2(n_2489),
.B(n_2576),
.C(n_2544),
.Y(n_2619)
);

AOI211xp5_ASAP7_75t_L g2620 ( 
.A1(n_2542),
.A2(n_234),
.B(n_231),
.C(n_233),
.Y(n_2620)
);

NAND4xp25_ASAP7_75t_L g2621 ( 
.A(n_2468),
.B(n_237),
.C(n_235),
.D(n_236),
.Y(n_2621)
);

AOI22xp5_ASAP7_75t_L g2622 ( 
.A1(n_2575),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_2622)
);

OAI21xp5_ASAP7_75t_L g2623 ( 
.A1(n_2511),
.A2(n_2430),
.B(n_2479),
.Y(n_2623)
);

O2A1O1Ixp33_ASAP7_75t_L g2624 ( 
.A1(n_2477),
.A2(n_241),
.B(n_238),
.C(n_240),
.Y(n_2624)
);

OAI221xp5_ASAP7_75t_L g2625 ( 
.A1(n_2519),
.A2(n_244),
.B1(n_241),
.B2(n_243),
.C(n_246),
.Y(n_2625)
);

NOR2x1_ASAP7_75t_L g2626 ( 
.A(n_2476),
.B(n_243),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2537),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2538),
.A2(n_2571),
.B(n_2541),
.Y(n_2628)
);

OAI22xp33_ASAP7_75t_L g2629 ( 
.A1(n_2563),
.A2(n_248),
.B1(n_244),
.B2(n_247),
.Y(n_2629)
);

NOR2xp67_ASAP7_75t_SL g2630 ( 
.A(n_2568),
.B(n_247),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2569),
.Y(n_2631)
);

AOI21xp33_ASAP7_75t_L g2632 ( 
.A1(n_2433),
.A2(n_248),
.B(n_249),
.Y(n_2632)
);

AOI322xp5_ASAP7_75t_L g2633 ( 
.A1(n_2459),
.A2(n_250),
.A3(n_251),
.B1(n_252),
.B2(n_253),
.C1(n_254),
.C2(n_255),
.Y(n_2633)
);

OAI22xp5_ASAP7_75t_L g2634 ( 
.A1(n_2566),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_2634)
);

AOI221xp5_ASAP7_75t_L g2635 ( 
.A1(n_2444),
.A2(n_257),
.B1(n_254),
.B2(n_256),
.C(n_258),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2496),
.B(n_256),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_SL g2637 ( 
.A(n_2545),
.B(n_257),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2505),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2567),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2441),
.Y(n_2640)
);

NAND5xp2_ASAP7_75t_L g2641 ( 
.A(n_2436),
.B(n_261),
.C(n_259),
.D(n_260),
.E(n_262),
.Y(n_2641)
);

OAI21xp5_ASAP7_75t_L g2642 ( 
.A1(n_2500),
.A2(n_259),
.B(n_260),
.Y(n_2642)
);

AOI222xp33_ASAP7_75t_L g2643 ( 
.A1(n_2516),
.A2(n_263),
.B1(n_264),
.B2(n_267),
.C1(n_270),
.C2(n_271),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2518),
.A2(n_272),
.B1(n_263),
.B2(n_271),
.Y(n_2644)
);

AOI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_2526),
.A2(n_276),
.B1(n_273),
.B2(n_274),
.Y(n_2645)
);

OAI322xp33_ASAP7_75t_L g2646 ( 
.A1(n_2529),
.A2(n_273),
.A3(n_276),
.B1(n_277),
.B2(n_278),
.C1(n_279),
.C2(n_280),
.Y(n_2646)
);

AO21x1_ASAP7_75t_L g2647 ( 
.A1(n_2467),
.A2(n_2452),
.B(n_2507),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2517),
.Y(n_2648)
);

NOR2xp67_ASAP7_75t_L g2649 ( 
.A(n_2521),
.B(n_2472),
.Y(n_2649)
);

OAI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_2486),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2517),
.Y(n_2651)
);

OAI22xp5_ASAP7_75t_L g2652 ( 
.A1(n_2491),
.A2(n_2451),
.B1(n_2470),
.B2(n_2455),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2522),
.Y(n_2653)
);

OAI322xp33_ASAP7_75t_L g2654 ( 
.A1(n_2506),
.A2(n_281),
.A3(n_282),
.B1(n_283),
.B2(n_284),
.C1(n_285),
.C2(n_286),
.Y(n_2654)
);

AOI211x1_ASAP7_75t_L g2655 ( 
.A1(n_2508),
.A2(n_284),
.B(n_281),
.C(n_282),
.Y(n_2655)
);

INVx1_ASAP7_75t_SL g2656 ( 
.A(n_2551),
.Y(n_2656)
);

OAI22xp5_ASAP7_75t_L g2657 ( 
.A1(n_2483),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_2657)
);

AOI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2528),
.A2(n_291),
.B1(n_288),
.B2(n_290),
.Y(n_2658)
);

XNOR2x1_ASAP7_75t_L g2659 ( 
.A(n_2520),
.B(n_290),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_2502),
.B(n_293),
.Y(n_2660)
);

OAI22xp5_ASAP7_75t_L g2661 ( 
.A1(n_2550),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_2661)
);

AOI21xp33_ASAP7_75t_L g2662 ( 
.A1(n_2503),
.A2(n_294),
.B(n_296),
.Y(n_2662)
);

AOI211xp5_ASAP7_75t_L g2663 ( 
.A1(n_2523),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_2663)
);

AOI211xp5_ASAP7_75t_L g2664 ( 
.A1(n_2514),
.A2(n_2482),
.B(n_2525),
.C(n_2524),
.Y(n_2664)
);

O2A1O1Ixp33_ASAP7_75t_L g2665 ( 
.A1(n_2596),
.A2(n_2490),
.B(n_2478),
.C(n_2448),
.Y(n_2665)
);

NOR2xp33_ASAP7_75t_L g2666 ( 
.A(n_2585),
.B(n_2473),
.Y(n_2666)
);

AOI32xp33_ASAP7_75t_L g2667 ( 
.A1(n_2579),
.A2(n_2487),
.A3(n_2447),
.B1(n_2458),
.B2(n_2481),
.Y(n_2667)
);

AND2x4_ASAP7_75t_L g2668 ( 
.A(n_2577),
.B(n_2463),
.Y(n_2668)
);

NAND3xp33_ASAP7_75t_SL g2669 ( 
.A(n_2592),
.B(n_2509),
.C(n_2460),
.Y(n_2669)
);

AOI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2589),
.A2(n_2504),
.B1(n_2446),
.B2(n_2554),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2648),
.Y(n_2671)
);

NOR2xp33_ASAP7_75t_R g2672 ( 
.A(n_2613),
.B(n_2485),
.Y(n_2672)
);

OAI321xp33_ASAP7_75t_L g2673 ( 
.A1(n_2623),
.A2(n_2457),
.A3(n_2439),
.B1(n_2462),
.B2(n_2501),
.C(n_2493),
.Y(n_2673)
);

AOI322xp5_ASAP7_75t_L g2674 ( 
.A1(n_2591),
.A2(n_2653),
.A3(n_2660),
.B1(n_2583),
.B2(n_2586),
.C1(n_2587),
.C2(n_2627),
.Y(n_2674)
);

NAND2xp33_ASAP7_75t_SL g2675 ( 
.A(n_2630),
.B(n_2510),
.Y(n_2675)
);

O2A1O1Ixp5_ASAP7_75t_L g2676 ( 
.A1(n_2637),
.A2(n_2488),
.B(n_2492),
.C(n_2497),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2651),
.Y(n_2677)
);

O2A1O1Ixp33_ASAP7_75t_L g2678 ( 
.A1(n_2609),
.A2(n_2494),
.B(n_2461),
.C(n_2442),
.Y(n_2678)
);

NAND3xp33_ASAP7_75t_SL g2679 ( 
.A(n_2608),
.B(n_2438),
.C(n_2445),
.Y(n_2679)
);

OAI211xp5_ASAP7_75t_SL g2680 ( 
.A1(n_2614),
.A2(n_2474),
.B(n_2484),
.C(n_2530),
.Y(n_2680)
);

OAI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2615),
.A2(n_2625),
.B1(n_2645),
.B2(n_2649),
.Y(n_2681)
);

AOI31xp33_ASAP7_75t_R g2682 ( 
.A1(n_2641),
.A2(n_2453),
.A3(n_2450),
.B(n_2499),
.Y(n_2682)
);

NAND3xp33_ASAP7_75t_L g2683 ( 
.A(n_2599),
.B(n_2453),
.C(n_2449),
.Y(n_2683)
);

NOR2xp33_ASAP7_75t_L g2684 ( 
.A(n_2613),
.B(n_2466),
.Y(n_2684)
);

OAI21xp5_ASAP7_75t_SL g2685 ( 
.A1(n_2590),
.A2(n_2513),
.B(n_2480),
.Y(n_2685)
);

INVx2_ASAP7_75t_SL g2686 ( 
.A(n_2578),
.Y(n_2686)
);

AOI21xp33_ASAP7_75t_L g2687 ( 
.A1(n_2619),
.A2(n_2533),
.B(n_298),
.Y(n_2687)
);

INVx1_ASAP7_75t_SL g2688 ( 
.A(n_2659),
.Y(n_2688)
);

OAI22xp5_ASAP7_75t_L g2689 ( 
.A1(n_2658),
.A2(n_2456),
.B1(n_301),
.B2(n_299),
.Y(n_2689)
);

CKINVDCx16_ASAP7_75t_R g2690 ( 
.A(n_2626),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2612),
.Y(n_2691)
);

INVxp67_ASAP7_75t_L g2692 ( 
.A(n_2636),
.Y(n_2692)
);

AOI221xp5_ASAP7_75t_L g2693 ( 
.A1(n_2632),
.A2(n_300),
.B1(n_302),
.B2(n_303),
.C(n_304),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2617),
.B(n_302),
.Y(n_2694)
);

AOI221xp5_ASAP7_75t_L g2695 ( 
.A1(n_2581),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.C(n_307),
.Y(n_2695)
);

AOI221xp5_ASAP7_75t_L g2696 ( 
.A1(n_2662),
.A2(n_308),
.B1(n_309),
.B2(n_311),
.C(n_312),
.Y(n_2696)
);

AO21x1_ASAP7_75t_L g2697 ( 
.A1(n_2624),
.A2(n_308),
.B(n_309),
.Y(n_2697)
);

OAI21xp33_ASAP7_75t_L g2698 ( 
.A1(n_2639),
.A2(n_312),
.B(n_313),
.Y(n_2698)
);

OA21x2_ASAP7_75t_L g2699 ( 
.A1(n_2602),
.A2(n_313),
.B(n_315),
.Y(n_2699)
);

OAI221xp5_ASAP7_75t_L g2700 ( 
.A1(n_2582),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.C(n_319),
.Y(n_2700)
);

AOI21xp33_ASAP7_75t_L g2701 ( 
.A1(n_2656),
.A2(n_317),
.B(n_319),
.Y(n_2701)
);

NOR4xp25_ASAP7_75t_SL g2702 ( 
.A(n_2607),
.B(n_323),
.C(n_320),
.D(n_322),
.Y(n_2702)
);

AOI21xp33_ASAP7_75t_SL g2703 ( 
.A1(n_2612),
.A2(n_320),
.B(n_322),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2628),
.B(n_323),
.Y(n_2704)
);

AOI21xp33_ASAP7_75t_SL g2705 ( 
.A1(n_2601),
.A2(n_324),
.B(n_326),
.Y(n_2705)
);

A2O1A1Ixp33_ASAP7_75t_L g2706 ( 
.A1(n_2584),
.A2(n_328),
.B(n_324),
.C(n_326),
.Y(n_2706)
);

O2A1O1Ixp33_ASAP7_75t_L g2707 ( 
.A1(n_2593),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_2707)
);

OAI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2603),
.A2(n_329),
.B(n_331),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2655),
.B(n_331),
.Y(n_2709)
);

NAND2xp33_ASAP7_75t_R g2710 ( 
.A(n_2597),
.B(n_332),
.Y(n_2710)
);

INVxp67_ASAP7_75t_L g2711 ( 
.A(n_2604),
.Y(n_2711)
);

NOR2x1_ASAP7_75t_L g2712 ( 
.A(n_2600),
.B(n_332),
.Y(n_2712)
);

AOI22xp5_ASAP7_75t_L g2713 ( 
.A1(n_2621),
.A2(n_336),
.B1(n_333),
.B2(n_334),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2598),
.Y(n_2714)
);

AOI221x1_ASAP7_75t_SL g2715 ( 
.A1(n_2664),
.A2(n_333),
.B1(n_336),
.B2(n_337),
.C(n_338),
.Y(n_2715)
);

AOI21xp33_ASAP7_75t_SL g2716 ( 
.A1(n_2644),
.A2(n_337),
.B(n_339),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2622),
.Y(n_2717)
);

NOR2x1_ASAP7_75t_L g2718 ( 
.A(n_2646),
.B(n_339),
.Y(n_2718)
);

AOI221x1_ASAP7_75t_SL g2719 ( 
.A1(n_2652),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.C(n_343),
.Y(n_2719)
);

BUFx6f_ASAP7_75t_L g2720 ( 
.A(n_2631),
.Y(n_2720)
);

AND2x6_ASAP7_75t_L g2721 ( 
.A(n_2638),
.B(n_340),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2588),
.B(n_343),
.Y(n_2722)
);

NAND4xp25_ASAP7_75t_L g2723 ( 
.A(n_2674),
.B(n_2580),
.C(n_2595),
.D(n_2620),
.Y(n_2723)
);

HB1xp67_ASAP7_75t_L g2724 ( 
.A(n_2691),
.Y(n_2724)
);

AO21x1_ASAP7_75t_L g2725 ( 
.A1(n_2675),
.A2(n_2629),
.B(n_2650),
.Y(n_2725)
);

AOI221xp5_ASAP7_75t_L g2726 ( 
.A1(n_2719),
.A2(n_2611),
.B1(n_2618),
.B2(n_2661),
.C(n_2605),
.Y(n_2726)
);

NAND3xp33_ASAP7_75t_L g2727 ( 
.A(n_2703),
.B(n_2643),
.C(n_2663),
.Y(n_2727)
);

INVxp33_ASAP7_75t_L g2728 ( 
.A(n_2672),
.Y(n_2728)
);

AOI22xp5_ASAP7_75t_L g2729 ( 
.A1(n_2666),
.A2(n_2634),
.B1(n_2657),
.B2(n_2640),
.Y(n_2729)
);

NAND2x1p5_ASAP7_75t_L g2730 ( 
.A(n_2668),
.B(n_2686),
.Y(n_2730)
);

AOI211xp5_ASAP7_75t_L g2731 ( 
.A1(n_2687),
.A2(n_2642),
.B(n_2647),
.C(n_2654),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2712),
.B(n_2606),
.Y(n_2732)
);

OAI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2670),
.A2(n_2610),
.B1(n_2594),
.B2(n_2616),
.Y(n_2733)
);

NOR2xp33_ASAP7_75t_L g2734 ( 
.A(n_2690),
.B(n_2635),
.Y(n_2734)
);

NOR4xp75_ASAP7_75t_L g2735 ( 
.A(n_2697),
.B(n_2633),
.C(n_348),
.D(n_345),
.Y(n_2735)
);

AOI22xp5_ASAP7_75t_L g2736 ( 
.A1(n_2671),
.A2(n_350),
.B1(n_347),
.B2(n_349),
.Y(n_2736)
);

XOR2x2_ASAP7_75t_L g2737 ( 
.A(n_2718),
.B(n_352),
.Y(n_2737)
);

AOI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2704),
.A2(n_352),
.B(n_353),
.Y(n_2738)
);

NOR2xp33_ASAP7_75t_L g2739 ( 
.A(n_2688),
.B(n_354),
.Y(n_2739)
);

CKINVDCx20_ASAP7_75t_R g2740 ( 
.A(n_2681),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2677),
.B(n_355),
.Y(n_2741)
);

AOI221x1_ASAP7_75t_L g2742 ( 
.A1(n_2714),
.A2(n_356),
.B1(n_357),
.B2(n_359),
.C(n_360),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2721),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2721),
.Y(n_2744)
);

AOI21xp5_ASAP7_75t_L g2745 ( 
.A1(n_2665),
.A2(n_360),
.B(n_361),
.Y(n_2745)
);

OAI22xp5_ASAP7_75t_L g2746 ( 
.A1(n_2713),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_2746)
);

OAI221xp5_ASAP7_75t_SL g2747 ( 
.A1(n_2667),
.A2(n_362),
.B1(n_364),
.B2(n_366),
.C(n_367),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_L g2748 ( 
.A(n_2698),
.B(n_364),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2721),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2699),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2715),
.B(n_368),
.Y(n_2751)
);

OAI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2711),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_2752)
);

OAI221xp5_ASAP7_75t_L g2753 ( 
.A1(n_2685),
.A2(n_369),
.B1(n_370),
.B2(n_371),
.C(n_372),
.Y(n_2753)
);

OAI211xp5_ASAP7_75t_L g2754 ( 
.A1(n_2708),
.A2(n_374),
.B(n_371),
.C(n_372),
.Y(n_2754)
);

INVx1_ASAP7_75t_SL g2755 ( 
.A(n_2694),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_SL g2756 ( 
.A(n_2720),
.B(n_374),
.Y(n_2756)
);

AOI22x1_ASAP7_75t_L g2757 ( 
.A1(n_2720),
.A2(n_2717),
.B1(n_2692),
.B2(n_2682),
.Y(n_2757)
);

CKINVDCx6p67_ASAP7_75t_R g2758 ( 
.A(n_2709),
.Y(n_2758)
);

OR2x2_ASAP7_75t_L g2759 ( 
.A(n_2750),
.B(n_2722),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2732),
.B(n_2730),
.Y(n_2760)
);

NOR2x1_ASAP7_75t_L g2761 ( 
.A(n_2743),
.B(n_2679),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2724),
.Y(n_2762)
);

AOI22xp5_ASAP7_75t_L g2763 ( 
.A1(n_2740),
.A2(n_2710),
.B1(n_2669),
.B2(n_2680),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2744),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2749),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2737),
.Y(n_2766)
);

INVxp33_ASAP7_75t_L g2767 ( 
.A(n_2739),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2725),
.Y(n_2768)
);

AOI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2734),
.A2(n_2696),
.B1(n_2695),
.B2(n_2684),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2741),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2758),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2752),
.Y(n_2772)
);

NOR2xp33_ASAP7_75t_L g2773 ( 
.A(n_2728),
.B(n_2705),
.Y(n_2773)
);

NOR2x1_ASAP7_75t_SL g2774 ( 
.A(n_2754),
.B(n_2683),
.Y(n_2774)
);

NOR2x1_ASAP7_75t_L g2775 ( 
.A(n_2723),
.B(n_2700),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2751),
.Y(n_2776)
);

NOR2x1_ASAP7_75t_L g2777 ( 
.A(n_2756),
.B(n_2707),
.Y(n_2777)
);

NOR2x1_ASAP7_75t_L g2778 ( 
.A(n_2727),
.B(n_2706),
.Y(n_2778)
);

NOR2x1_ASAP7_75t_L g2779 ( 
.A(n_2768),
.B(n_2738),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_L g2780 ( 
.A(n_2762),
.B(n_2747),
.Y(n_2780)
);

NOR2x1_ASAP7_75t_L g2781 ( 
.A(n_2760),
.B(n_2745),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2774),
.Y(n_2782)
);

OAI22xp5_ASAP7_75t_L g2783 ( 
.A1(n_2763),
.A2(n_2753),
.B1(n_2769),
.B2(n_2729),
.Y(n_2783)
);

NOR2x1_ASAP7_75t_L g2784 ( 
.A(n_2761),
.B(n_2748),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2759),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2764),
.B(n_2702),
.Y(n_2786)
);

XNOR2xp5_ASAP7_75t_L g2787 ( 
.A(n_2775),
.B(n_2735),
.Y(n_2787)
);

INVxp67_ASAP7_75t_L g2788 ( 
.A(n_2773),
.Y(n_2788)
);

NAND2x1p5_ASAP7_75t_L g2789 ( 
.A(n_2777),
.B(n_2757),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2765),
.Y(n_2790)
);

NOR2x1_ASAP7_75t_L g2791 ( 
.A(n_2778),
.B(n_2755),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2771),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2766),
.Y(n_2793)
);

INVx3_ASAP7_75t_L g2794 ( 
.A(n_2770),
.Y(n_2794)
);

CKINVDCx20_ASAP7_75t_R g2795 ( 
.A(n_2769),
.Y(n_2795)
);

OAI22xp5_ASAP7_75t_L g2796 ( 
.A1(n_2795),
.A2(n_2731),
.B1(n_2772),
.B2(n_2767),
.Y(n_2796)
);

NAND3xp33_ASAP7_75t_SL g2797 ( 
.A(n_2789),
.B(n_2726),
.C(n_2693),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2790),
.Y(n_2798)
);

OAI322xp33_ASAP7_75t_L g2799 ( 
.A1(n_2782),
.A2(n_2733),
.A3(n_2776),
.B1(n_2689),
.B2(n_2678),
.C1(n_2716),
.C2(n_2746),
.Y(n_2799)
);

NAND4xp75_ASAP7_75t_L g2800 ( 
.A(n_2781),
.B(n_2742),
.C(n_2701),
.D(n_2736),
.Y(n_2800)
);

OAI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2792),
.A2(n_2736),
.B1(n_2673),
.B2(n_2676),
.Y(n_2801)
);

AOI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2780),
.A2(n_2793),
.B1(n_2791),
.B2(n_2783),
.Y(n_2802)
);

A2O1A1Ixp33_ASAP7_75t_L g2803 ( 
.A1(n_2785),
.A2(n_377),
.B(n_375),
.C(n_376),
.Y(n_2803)
);

NAND4xp25_ASAP7_75t_L g2804 ( 
.A(n_2784),
.B(n_378),
.C(n_376),
.D(n_377),
.Y(n_2804)
);

OAI211xp5_ASAP7_75t_L g2805 ( 
.A1(n_2786),
.A2(n_378),
.B(n_379),
.C(n_381),
.Y(n_2805)
);

AOI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2787),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_2806)
);

OR2x2_ASAP7_75t_L g2807 ( 
.A(n_2794),
.B(n_2788),
.Y(n_2807)
);

AOI21xp33_ASAP7_75t_L g2808 ( 
.A1(n_2779),
.A2(n_382),
.B(n_383),
.Y(n_2808)
);

AOI221xp5_ASAP7_75t_L g2809 ( 
.A1(n_2783),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.C(n_386),
.Y(n_2809)
);

OAI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2795),
.A2(n_384),
.B1(n_387),
.B2(n_388),
.Y(n_2810)
);

XOR2xp5_ASAP7_75t_L g2811 ( 
.A(n_2787),
.B(n_388),
.Y(n_2811)
);

NOR3xp33_ASAP7_75t_L g2812 ( 
.A(n_2783),
.B(n_389),
.C(n_391),
.Y(n_2812)
);

AO22x2_ASAP7_75t_L g2813 ( 
.A1(n_2783),
.A2(n_389),
.B1(n_391),
.B2(n_392),
.Y(n_2813)
);

NOR3x2_ASAP7_75t_L g2814 ( 
.A(n_2781),
.B(n_392),
.C(n_393),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2811),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2813),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2814),
.Y(n_2817)
);

NAND3xp33_ASAP7_75t_SL g2818 ( 
.A(n_2812),
.B(n_393),
.C(n_394),
.Y(n_2818)
);

NAND3xp33_ASAP7_75t_L g2819 ( 
.A(n_2802),
.B(n_395),
.C(n_396),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2813),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2800),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2798),
.Y(n_2822)
);

XOR2xp5_ASAP7_75t_L g2823 ( 
.A(n_2796),
.B(n_396),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2807),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2806),
.Y(n_2825)
);

NOR2xp33_ASAP7_75t_L g2826 ( 
.A(n_2804),
.B(n_398),
.Y(n_2826)
);

AND2x4_ASAP7_75t_L g2827 ( 
.A(n_2803),
.B(n_398),
.Y(n_2827)
);

AO22x2_ASAP7_75t_L g2828 ( 
.A1(n_2801),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.Y(n_2828)
);

HB1xp67_ASAP7_75t_L g2829 ( 
.A(n_2810),
.Y(n_2829)
);

NOR2x1_ASAP7_75t_L g2830 ( 
.A(n_2805),
.B(n_400),
.Y(n_2830)
);

OR2x2_ASAP7_75t_L g2831 ( 
.A(n_2797),
.B(n_401),
.Y(n_2831)
);

XNOR2xp5_ASAP7_75t_L g2832 ( 
.A(n_2809),
.B(n_402),
.Y(n_2832)
);

NAND3x1_ASAP7_75t_L g2833 ( 
.A(n_2799),
.B(n_403),
.C(n_405),
.Y(n_2833)
);

AND2x4_ASAP7_75t_L g2834 ( 
.A(n_2808),
.B(n_405),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2813),
.Y(n_2835)
);

OAI22xp5_ASAP7_75t_L g2836 ( 
.A1(n_2831),
.A2(n_406),
.B1(n_407),
.B2(n_409),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2822),
.B(n_406),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2828),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2828),
.Y(n_2839)
);

XNOR2x1_ASAP7_75t_SL g2840 ( 
.A(n_2820),
.B(n_407),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2816),
.B(n_409),
.Y(n_2841)
);

XOR2xp5_ASAP7_75t_L g2842 ( 
.A(n_2823),
.B(n_410),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2835),
.Y(n_2843)
);

HB1xp67_ASAP7_75t_L g2844 ( 
.A(n_2830),
.Y(n_2844)
);

NOR3xp33_ASAP7_75t_L g2845 ( 
.A(n_2821),
.B(n_2824),
.C(n_2819),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2833),
.Y(n_2846)
);

INVx3_ASAP7_75t_L g2847 ( 
.A(n_2817),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2826),
.Y(n_2848)
);

XNOR2xp5_ASAP7_75t_L g2849 ( 
.A(n_2832),
.B(n_410),
.Y(n_2849)
);

XNOR2xp5_ASAP7_75t_L g2850 ( 
.A(n_2815),
.B(n_411),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2837),
.Y(n_2851)
);

OAI22x1_ASAP7_75t_L g2852 ( 
.A1(n_2842),
.A2(n_2834),
.B1(n_2827),
.B2(n_2825),
.Y(n_2852)
);

OAI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2842),
.A2(n_2829),
.B1(n_2818),
.B2(n_413),
.Y(n_2853)
);

INVxp67_ASAP7_75t_L g2854 ( 
.A(n_2841),
.Y(n_2854)
);

OR4x1_ASAP7_75t_L g2855 ( 
.A(n_2843),
.B(n_411),
.C(n_412),
.D(n_413),
.Y(n_2855)
);

NOR4xp25_ASAP7_75t_L g2856 ( 
.A(n_2838),
.B(n_412),
.C(n_414),
.D(n_416),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2840),
.Y(n_2857)
);

OAI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2849),
.A2(n_414),
.B(n_416),
.Y(n_2858)
);

OAI22xp5_ASAP7_75t_SL g2859 ( 
.A1(n_2846),
.A2(n_417),
.B1(n_418),
.B2(n_420),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2850),
.Y(n_2860)
);

AND2x4_ASAP7_75t_L g2861 ( 
.A(n_2845),
.B(n_421),
.Y(n_2861)
);

OAI22xp5_ASAP7_75t_SL g2862 ( 
.A1(n_2839),
.A2(n_421),
.B1(n_422),
.B2(n_423),
.Y(n_2862)
);

AOI22xp5_ASAP7_75t_L g2863 ( 
.A1(n_2847),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.Y(n_2863)
);

AOI211xp5_ASAP7_75t_SL g2864 ( 
.A1(n_2844),
.A2(n_2848),
.B(n_2836),
.C(n_426),
.Y(n_2864)
);

CKINVDCx5p33_ASAP7_75t_R g2865 ( 
.A(n_2852),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2861),
.Y(n_2866)
);

AOI21x1_ASAP7_75t_L g2867 ( 
.A1(n_2857),
.A2(n_424),
.B(n_425),
.Y(n_2867)
);

AOI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2853),
.A2(n_426),
.B1(n_428),
.B2(n_429),
.Y(n_2868)
);

HB1xp67_ASAP7_75t_L g2869 ( 
.A(n_2862),
.Y(n_2869)
);

OAI22xp5_ASAP7_75t_SL g2870 ( 
.A1(n_2855),
.A2(n_2856),
.B1(n_2858),
.B2(n_2859),
.Y(n_2870)
);

AOI22xp5_ASAP7_75t_L g2871 ( 
.A1(n_2860),
.A2(n_428),
.B1(n_430),
.B2(n_431),
.Y(n_2871)
);

AO221x2_ASAP7_75t_L g2872 ( 
.A1(n_2851),
.A2(n_430),
.B1(n_435),
.B2(n_436),
.C(n_438),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2863),
.Y(n_2873)
);

XNOR2xp5_ASAP7_75t_L g2874 ( 
.A(n_2854),
.B(n_436),
.Y(n_2874)
);

XNOR2xp5_ASAP7_75t_L g2875 ( 
.A(n_2864),
.B(n_438),
.Y(n_2875)
);

OAI21xp5_ASAP7_75t_L g2876 ( 
.A1(n_2853),
.A2(n_439),
.B(n_441),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2861),
.Y(n_2877)
);

INVxp67_ASAP7_75t_L g2878 ( 
.A(n_2861),
.Y(n_2878)
);

AOI22x1_ASAP7_75t_L g2879 ( 
.A1(n_2852),
.A2(n_442),
.B1(n_443),
.B2(n_444),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2867),
.Y(n_2880)
);

OAI22xp5_ASAP7_75t_SL g2881 ( 
.A1(n_2870),
.A2(n_442),
.B1(n_443),
.B2(n_445),
.Y(n_2881)
);

OAI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2865),
.A2(n_446),
.B1(n_447),
.B2(n_448),
.Y(n_2882)
);

CKINVDCx5p33_ASAP7_75t_R g2883 ( 
.A(n_2875),
.Y(n_2883)
);

BUFx2_ASAP7_75t_L g2884 ( 
.A(n_2876),
.Y(n_2884)
);

OAI22xp5_ASAP7_75t_SL g2885 ( 
.A1(n_2869),
.A2(n_446),
.B1(n_447),
.B2(n_449),
.Y(n_2885)
);

CKINVDCx20_ASAP7_75t_R g2886 ( 
.A(n_2878),
.Y(n_2886)
);

OAI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2868),
.A2(n_451),
.B1(n_452),
.B2(n_454),
.Y(n_2887)
);

AOI22xp5_ASAP7_75t_L g2888 ( 
.A1(n_2866),
.A2(n_454),
.B1(n_455),
.B2(n_456),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2879),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2874),
.Y(n_2890)
);

AO22x2_ASAP7_75t_L g2891 ( 
.A1(n_2877),
.A2(n_456),
.B1(n_457),
.B2(n_458),
.Y(n_2891)
);

OAI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_2886),
.A2(n_2873),
.B(n_2871),
.Y(n_2892)
);

AOI22xp33_ASAP7_75t_L g2893 ( 
.A1(n_2889),
.A2(n_2872),
.B1(n_460),
.B2(n_462),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2880),
.A2(n_2872),
.B(n_460),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2882),
.B(n_2887),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_L g2896 ( 
.A1(n_2883),
.A2(n_459),
.B1(n_463),
.B2(n_464),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2891),
.Y(n_2897)
);

BUFx3_ASAP7_75t_L g2898 ( 
.A(n_2884),
.Y(n_2898)
);

AOI22xp33_ASAP7_75t_L g2899 ( 
.A1(n_2890),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_2899)
);

OAI21xp5_ASAP7_75t_L g2900 ( 
.A1(n_2888),
.A2(n_465),
.B(n_466),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2891),
.Y(n_2901)
);

AOI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2881),
.A2(n_468),
.B(n_469),
.Y(n_2902)
);

OA21x2_ASAP7_75t_L g2903 ( 
.A1(n_2892),
.A2(n_2897),
.B(n_2901),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2902),
.Y(n_2904)
);

AOI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2894),
.A2(n_2885),
.B(n_470),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2898),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2893),
.B(n_468),
.Y(n_2907)
);

NAND3xp33_ASAP7_75t_L g2908 ( 
.A(n_2900),
.B(n_2895),
.C(n_2899),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2896),
.Y(n_2909)
);

XNOR2xp5_ASAP7_75t_L g2910 ( 
.A(n_2898),
.B(n_470),
.Y(n_2910)
);

AOI21xp5_ASAP7_75t_L g2911 ( 
.A1(n_2894),
.A2(n_471),
.B(n_472),
.Y(n_2911)
);

A2O1A1Ixp33_ASAP7_75t_L g2912 ( 
.A1(n_2902),
.A2(n_472),
.B(n_474),
.C(n_475),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2912),
.B(n_2911),
.Y(n_2913)
);

AOI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2906),
.A2(n_475),
.B1(n_476),
.B2(n_477),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2905),
.A2(n_2903),
.B(n_2908),
.Y(n_2915)
);

AOI22xp33_ASAP7_75t_SL g2916 ( 
.A1(n_2907),
.A2(n_476),
.B1(n_477),
.B2(n_478),
.Y(n_2916)
);

AOI322xp5_ASAP7_75t_L g2917 ( 
.A1(n_2913),
.A2(n_2904),
.A3(n_2909),
.B1(n_2903),
.B2(n_2910),
.C1(n_483),
.C2(n_484),
.Y(n_2917)
);

OR2x6_ASAP7_75t_L g2918 ( 
.A(n_2917),
.B(n_2915),
.Y(n_2918)
);

AOI221xp5_ASAP7_75t_L g2919 ( 
.A1(n_2918),
.A2(n_2916),
.B1(n_2914),
.B2(n_480),
.C(n_481),
.Y(n_2919)
);

AOI211xp5_ASAP7_75t_L g2920 ( 
.A1(n_2919),
.A2(n_478),
.B(n_479),
.C(n_483),
.Y(n_2920)
);


endmodule