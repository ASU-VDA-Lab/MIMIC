module fake_netlist_5_1984_n_993 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_46, n_233, n_21, n_94, n_203, n_245, n_205, n_113, n_38, n_123, n_139, n_105, n_246, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_258, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_247, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_243, n_239, n_175, n_252, n_169, n_59, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_253, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_204, n_50, n_250, n_52, n_88, n_110, n_216, n_993);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_258;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_175;
input n_252;
input n_169;
input n_59;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_88;
input n_110;
input n_216;

output n_993;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_419;
wire n_318;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_785;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_525;
wire n_397;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_677;
wire n_859;
wire n_864;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_449;
wire n_325;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_942;
wire n_381;
wire n_291;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_570;
wire n_457;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_839;
wire n_727;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_388;
wire n_761;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_338;
wire n_571;
wire n_477;
wire n_333;
wire n_461;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_283;
wire n_383;
wire n_711;
wire n_834;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_891;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_699;
wire n_632;
wire n_979;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_846;
wire n_586;
wire n_748;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_966;
wire n_987;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_647;
wire n_710;
wire n_707;
wire n_795;
wire n_832;
wire n_857;
wire n_695;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_327;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_352;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_222),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_30),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_51),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_255),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_89),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_214),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_121),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_147),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_111),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_162),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_165),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_81),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_174),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_199),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_106),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_49),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_41),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_85),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_135),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_187),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_28),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_71),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_142),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_70),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_143),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_141),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_90),
.Y(n_289)
);

BUFx8_ASAP7_75t_SL g290 ( 
.A(n_18),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_160),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_6),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_212),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_77),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_208),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_149),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_130),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_231),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_36),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_154),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_168),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_123),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_118),
.Y(n_305)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_227),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_32),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_205),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_236),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_196),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_218),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_1),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_115),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_8),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_117),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_140),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_114),
.Y(n_318)
);

INVx4_ASAP7_75t_R g319 ( 
.A(n_210),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_202),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_44),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_150),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_152),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_251),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_103),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_15),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_244),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_3),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_75),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_241),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_158),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_217),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_195),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_84),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_40),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_234),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_124),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_228),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_151),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_79),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_119),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_224),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_24),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_69),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_39),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_248),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_164),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_52),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_109),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_166),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_148),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_60),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_133),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_99),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_68),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_50),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_181),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_87),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_98),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_129),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_144),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_92),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_43),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_190),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_5),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_250),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_42),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_65),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_215),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_107),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_167),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_53),
.Y(n_372)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_86),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_206),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_122),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_178),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_180),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_155),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_136),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_145),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_24),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_156),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_8),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_242),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_235),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_204),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_116),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_16),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_237),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_11),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_9),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_74),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_58),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_246),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_108),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_100),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_229),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_226),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_112),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_230),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_110),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_225),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_193),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_2),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_189),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_258),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_243),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_4),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_17),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_169),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_223),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_163),
.Y(n_412)
);

BUFx2_ASAP7_75t_SL g413 ( 
.A(n_57),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_59),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_240),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_159),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_153),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_127),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_177),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_207),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_194),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_120),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_252),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_173),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_76),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_138),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_34),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_171),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_211),
.Y(n_429)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_54),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_221),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_21),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_26),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_16),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_83),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_268),
.B(n_0),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_306),
.B(n_0),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_408),
.B(n_1),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_276),
.B(n_2),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_3),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_263),
.B(n_4),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_304),
.B(n_5),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_6),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_373),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_373),
.Y(n_446)
);

BUFx12f_ASAP7_75t_L g447 ( 
.A(n_266),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_263),
.B(n_7),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_269),
.B(n_7),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_269),
.B(n_9),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_290),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_285),
.B(n_10),
.Y(n_453)
);

INVx5_ASAP7_75t_L g454 ( 
.A(n_353),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_266),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_353),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_285),
.B(n_10),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_373),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_294),
.B(n_12),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_422),
.B(n_12),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_373),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_294),
.B(n_302),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_279),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_264),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_302),
.B(n_13),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_13),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_391),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_261),
.B(n_14),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_292),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_265),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_329),
.B(n_14),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_329),
.B(n_15),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_279),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_367),
.B(n_17),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_367),
.B(n_19),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_267),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_395),
.B(n_19),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_308),
.Y(n_483)
);

BUFx12f_ASAP7_75t_L g484 ( 
.A(n_262),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_274),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_321),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_271),
.Y(n_487)
);

BUFx8_ASAP7_75t_SL g488 ( 
.A(n_343),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_313),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_373),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_272),
.Y(n_491)
);

CKINVDCx6p67_ASAP7_75t_R g492 ( 
.A(n_345),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_326),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_395),
.B(n_402),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_402),
.B(n_20),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_414),
.B(n_20),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_414),
.B(n_21),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_373),
.B(n_22),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_260),
.B(n_22),
.Y(n_499)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_413),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_434),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_270),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_273),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_275),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_278),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_282),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_283),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_277),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_293),
.B(n_23),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_289),
.B(n_425),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_296),
.B(n_298),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_300),
.B(n_25),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_315),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_301),
.B(n_26),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_303),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_280),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_307),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_319),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_312),
.B(n_37),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_322),
.B(n_27),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_409),
.B(n_27),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_328),
.B(n_28),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_365),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_330),
.B(n_29),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_381),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_388),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_332),
.B(n_29),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_390),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_404),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_333),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_335),
.B(n_38),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_427),
.B(n_31),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_432),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_337),
.B(n_31),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_433),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_510),
.A2(n_378),
.B1(n_406),
.B2(n_377),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_485),
.B(n_338),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_518),
.B(n_281),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_436),
.Y(n_539)
);

AO22x2_ASAP7_75t_L g540 ( 
.A1(n_439),
.A2(n_348),
.B1(n_349),
.B2(n_344),
.Y(n_540)
);

AO22x2_ASAP7_75t_L g541 ( 
.A1(n_462),
.A2(n_360),
.B1(n_363),
.B2(n_355),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_521),
.A2(n_420),
.B1(n_374),
.B2(n_375),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_444),
.A2(n_286),
.B1(n_287),
.B2(n_284),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_436),
.Y(n_544)
);

OAI22xp33_ASAP7_75t_L g545 ( 
.A1(n_473),
.A2(n_382),
.B1(n_385),
.B2(n_369),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_463),
.A2(n_291),
.B1(n_295),
.B2(n_288),
.Y(n_546)
);

OA22x2_ASAP7_75t_L g547 ( 
.A1(n_513),
.A2(n_398),
.B1(n_400),
.B2(n_392),
.Y(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_462),
.A2(n_423),
.B1(n_417),
.B2(n_418),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_518),
.B(n_485),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_L g550 ( 
.A1(n_496),
.A2(n_412),
.B1(n_419),
.B2(n_424),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_518),
.Y(n_551)
);

AO22x2_ASAP7_75t_L g552 ( 
.A1(n_497),
.A2(n_428),
.B1(n_33),
.B2(n_35),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_469),
.A2(n_438),
.B1(n_484),
.B2(n_443),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_522),
.A2(n_362),
.B1(n_431),
.B2(n_429),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_485),
.B(n_297),
.Y(n_555)
);

AO22x2_ASAP7_75t_L g556 ( 
.A1(n_497),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_486),
.B(n_299),
.Y(n_557)
);

AO22x2_ASAP7_75t_L g558 ( 
.A1(n_499),
.A2(n_435),
.B1(n_426),
.B2(n_421),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_478),
.A2(n_416),
.B1(n_415),
.B2(n_411),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_449),
.Y(n_560)
);

OA22x2_ASAP7_75t_L g561 ( 
.A1(n_523),
.A2(n_410),
.B1(n_407),
.B2(n_405),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_449),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_532),
.A2(n_529),
.B1(n_535),
.B2(n_525),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_525),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_467),
.B(n_401),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_529),
.A2(n_399),
.B1(n_397),
.B2(n_396),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_535),
.A2(n_351),
.B1(n_394),
.B2(n_393),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_447),
.B(n_305),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_460),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_507),
.A2(n_389),
.B1(n_387),
.B2(n_386),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_456),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_460),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_521),
.A2(n_452),
.B1(n_466),
.B2(n_455),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_478),
.B(n_309),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_437),
.A2(n_441),
.B1(n_440),
.B2(n_498),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_486),
.B(n_310),
.Y(n_576)
);

AO22x2_ASAP7_75t_L g577 ( 
.A1(n_499),
.A2(n_384),
.B1(n_380),
.B2(n_379),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_502),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_533),
.B(n_311),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_514),
.A2(n_342),
.B1(n_371),
.B2(n_370),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_478),
.B(n_481),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_527),
.A2(n_376),
.B1(n_368),
.B2(n_366),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_491),
.B(n_503),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_475),
.A2(n_339),
.B1(n_361),
.B2(n_359),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_470),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_487),
.B(n_314),
.Y(n_586)
);

AO22x2_ASAP7_75t_L g587 ( 
.A1(n_509),
.A2(n_364),
.B1(n_358),
.B2(n_357),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_516),
.B(n_316),
.Y(n_588)
);

AO22x2_ASAP7_75t_L g589 ( 
.A1(n_509),
.A2(n_524),
.B1(n_442),
.B2(n_448),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_503),
.B(n_317),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_517),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_504),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_459),
.B(n_318),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_459),
.B(n_320),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_508),
.B(n_323),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_450),
.A2(n_356),
.B1(n_354),
.B2(n_352),
.Y(n_596)
);

AO22x2_ASAP7_75t_L g597 ( 
.A1(n_524),
.A2(n_350),
.B1(n_347),
.B2(n_346),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_L g598 ( 
.A1(n_451),
.A2(n_341),
.B1(n_340),
.B2(n_336),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_504),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_465),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_526),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_471),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_504),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_530),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_482),
.A2(n_331),
.B1(n_327),
.B2(n_325),
.Y(n_605)
);

AO22x2_ASAP7_75t_L g606 ( 
.A1(n_453),
.A2(n_479),
.B1(n_495),
.B2(n_458),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_512),
.A2(n_334),
.B1(n_324),
.B2(n_47),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_530),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_539),
.Y(n_609)
);

INVxp33_ASAP7_75t_SL g610 ( 
.A(n_536),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_600),
.B(n_508),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_544),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_585),
.Y(n_613)
);

BUFx8_ASAP7_75t_L g614 ( 
.A(n_588),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_526),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_602),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_592),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_560),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_599),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_604),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_608),
.Y(n_621)
);

XNOR2x2_ASAP7_75t_L g622 ( 
.A(n_556),
.B(n_468),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_603),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_569),
.Y(n_624)
);

NOR2xp67_ASAP7_75t_L g625 ( 
.A(n_551),
.B(n_500),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_571),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_594),
.B(n_564),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_573),
.B(n_492),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_581),
.B(n_526),
.Y(n_629)
);

OR2x6_ASAP7_75t_L g630 ( 
.A(n_556),
.B(n_520),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_545),
.B(n_500),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g632 ( 
.A(n_542),
.B(n_561),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_553),
.B(n_563),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_584),
.B(n_500),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_572),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_565),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_562),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_579),
.B(n_528),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_578),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_606),
.B(n_445),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_591),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_562),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_589),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_589),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_575),
.B(n_511),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_547),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_586),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_550),
.B(n_528),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_537),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_541),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_543),
.A2(n_477),
.B(n_476),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_541),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_566),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g654 ( 
.A(n_606),
.B(n_488),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_596),
.B(n_480),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_548),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_567),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_548),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_540),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_R g660 ( 
.A(n_568),
.B(n_494),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_555),
.B(n_472),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_540),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_557),
.B(n_494),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_549),
.B(n_446),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_576),
.B(n_595),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_583),
.B(n_601),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_538),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_570),
.B(n_493),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_552),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_605),
.B(n_530),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_552),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_574),
.B(n_493),
.Y(n_672)
);

XOR2x2_ASAP7_75t_L g673 ( 
.A(n_580),
.B(n_534),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_607),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_590),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_582),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_546),
.Y(n_677)
);

XOR2x2_ASAP7_75t_L g678 ( 
.A(n_554),
.B(n_45),
.Y(n_678)
);

INVxp67_ASAP7_75t_SL g679 ( 
.A(n_598),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_558),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_559),
.B(n_505),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_558),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_577),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_568),
.A2(n_531),
.B(n_519),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_577),
.B(n_505),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_587),
.B(n_506),
.Y(n_686)
);

XOR2xp5_ASAP7_75t_L g687 ( 
.A(n_587),
.B(n_46),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_597),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_645),
.B(n_597),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_639),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_645),
.B(n_457),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_641),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_663),
.B(n_457),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_663),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_665),
.B(n_519),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_646),
.B(n_519),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_661),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_655),
.B(n_461),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_643),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_640),
.A2(n_531),
.B(n_490),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_655),
.B(n_464),
.Y(n_701)
);

INVxp33_ASAP7_75t_L g702 ( 
.A(n_627),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_649),
.B(n_474),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_676),
.B(n_454),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_623),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_617),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_666),
.B(n_474),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_640),
.A2(n_531),
.B(n_454),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_672),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_619),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_620),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_621),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_609),
.Y(n_713)
);

AND2x2_ASAP7_75t_SL g714 ( 
.A(n_644),
.B(n_674),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_664),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_611),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_659),
.B(n_483),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_613),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_616),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_664),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_670),
.B(n_515),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_612),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_675),
.B(n_515),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_667),
.B(n_48),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_650),
.B(n_55),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_651),
.B(n_483),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_618),
.Y(n_727)
);

AND2x2_ASAP7_75t_SL g728 ( 
.A(n_662),
.B(n_489),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_651),
.B(n_489),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_679),
.B(n_677),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_679),
.B(n_501),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_670),
.B(n_454),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_672),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_647),
.B(n_501),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_668),
.B(n_56),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_636),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_637),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_668),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_638),
.B(n_61),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_626),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_615),
.B(n_62),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_671),
.B(n_63),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_652),
.B(n_259),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_630),
.B(n_64),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_635),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_624),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_610),
.B(n_66),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_642),
.Y(n_748)
);

NAND2x1p5_ASAP7_75t_L g749 ( 
.A(n_656),
.B(n_67),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_658),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_629),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_631),
.B(n_72),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_669),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_614),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_648),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_631),
.B(n_73),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_681),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_685),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_684),
.B(n_78),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_688),
.B(n_80),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_734),
.Y(n_761)
);

HB1xp67_ASAP7_75t_SL g762 ( 
.A(n_754),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_694),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_694),
.Y(n_764)
);

BUFx12f_ASAP7_75t_L g765 ( 
.A(n_754),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_706),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_725),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_SL g768 ( 
.A(n_747),
.B(n_684),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_702),
.B(n_633),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_699),
.Y(n_770)
);

NAND2x1_ASAP7_75t_SL g771 ( 
.A(n_696),
.B(n_685),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_694),
.B(n_682),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_710),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_698),
.B(n_673),
.Y(n_774)
);

NAND2x1p5_ASAP7_75t_L g775 ( 
.A(n_709),
.B(n_743),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_733),
.B(n_634),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_709),
.B(n_680),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_733),
.B(n_683),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_736),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_755),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_755),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_718),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_698),
.B(n_701),
.Y(n_783)
);

NOR2x1_ASAP7_75t_R g784 ( 
.A(n_709),
.B(n_622),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_738),
.B(n_686),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_731),
.B(n_686),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_693),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_718),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_738),
.B(n_653),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_701),
.B(n_632),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_750),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_SL g792 ( 
.A(n_749),
.B(n_657),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_693),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_731),
.B(n_678),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_753),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_753),
.B(n_697),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_690),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_707),
.B(n_628),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_743),
.B(n_625),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_692),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_758),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_759),
.B(n_614),
.Y(n_802)
);

BUFx12f_ASAP7_75t_L g803 ( 
.A(n_730),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_755),
.Y(n_804)
);

BUFx12f_ASAP7_75t_L g805 ( 
.A(n_717),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_SL g806 ( 
.A(n_749),
.B(n_687),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_710),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_724),
.B(n_751),
.Y(n_808)
);

NAND2x1p5_ASAP7_75t_L g809 ( 
.A(n_764),
.B(n_724),
.Y(n_809)
);

BUFx24_ASAP7_75t_L g810 ( 
.A(n_789),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_779),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_796),
.Y(n_812)
);

BUFx4f_ASAP7_75t_L g813 ( 
.A(n_765),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_796),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_805),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_764),
.B(n_724),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_803),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_762),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_780),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_795),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_783),
.B(n_715),
.Y(n_821)
);

BUFx12f_ASAP7_75t_L g822 ( 
.A(n_789),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_797),
.Y(n_823)
);

BUFx8_ASAP7_75t_L g824 ( 
.A(n_798),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_800),
.Y(n_825)
);

INVx5_ASAP7_75t_L g826 ( 
.A(n_780),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_763),
.B(n_735),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_774),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_786),
.B(n_715),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_767),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_770),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_766),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_780),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_775),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_768),
.A2(n_691),
.B1(n_689),
.B2(n_714),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_767),
.Y(n_836)
);

INVx5_ASAP7_75t_L g837 ( 
.A(n_780),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_835),
.A2(n_768),
.B1(n_794),
.B2(n_689),
.Y(n_838)
);

BUFx10_ASAP7_75t_L g839 ( 
.A(n_831),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_823),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_826),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_825),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_828),
.A2(n_769),
.B1(n_806),
.B2(n_790),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_821),
.A2(n_806),
.B1(n_691),
.B2(n_792),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_829),
.A2(n_792),
.B1(n_726),
.B2(n_729),
.Y(n_845)
);

CKINVDCx11_ASAP7_75t_R g846 ( 
.A(n_822),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_L g847 ( 
.A1(n_828),
.A2(n_790),
.B1(n_702),
.B2(n_757),
.Y(n_847)
);

CKINVDCx11_ASAP7_75t_R g848 ( 
.A(n_815),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_811),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_832),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_812),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_814),
.Y(n_852)
);

INVx8_ASAP7_75t_L g853 ( 
.A(n_826),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_820),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_830),
.A2(n_726),
.B1(n_729),
.B2(n_714),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_818),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_819),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_824),
.A2(n_769),
.B1(n_716),
.B2(n_723),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_838),
.B(n_744),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_856),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_844),
.A2(n_843),
.B1(n_858),
.B2(n_845),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_844),
.A2(n_838),
.B1(n_847),
.B2(n_654),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_842),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_845),
.B(n_744),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_855),
.A2(n_801),
.B1(n_809),
.B2(n_816),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_855),
.A2(n_809),
.B1(n_816),
.B2(n_808),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_840),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_847),
.A2(n_802),
.B1(n_752),
.B2(n_756),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_850),
.Y(n_869)
);

BUFx12f_ASAP7_75t_L g870 ( 
.A(n_848),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_852),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_851),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_849),
.A2(n_785),
.B1(n_760),
.B2(n_732),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_854),
.A2(n_732),
.B1(n_761),
.B2(n_707),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_857),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_846),
.A2(n_739),
.B1(n_704),
.B2(n_776),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_841),
.Y(n_877)
);

BUFx12f_ASAP7_75t_SL g878 ( 
.A(n_841),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_853),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_846),
.A2(n_739),
.B1(n_704),
.B2(n_776),
.Y(n_880)
);

OAI22xp33_ASAP7_75t_SL g881 ( 
.A1(n_839),
.A2(n_721),
.B1(n_827),
.B2(n_777),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_839),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_861),
.A2(n_848),
.B1(n_720),
.B2(n_712),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_862),
.A2(n_703),
.B1(n_793),
.B2(n_787),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_867),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_863),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_860),
.B(n_784),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_859),
.A2(n_712),
.B1(n_711),
.B2(n_745),
.Y(n_888)
);

OAI22xp33_ASAP7_75t_L g889 ( 
.A1(n_859),
.A2(n_660),
.B1(n_810),
.B2(n_834),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_864),
.A2(n_711),
.B1(n_745),
.B2(n_703),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_868),
.A2(n_773),
.B1(n_807),
.B2(n_817),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_L g892 ( 
.A(n_881),
.B(n_741),
.C(n_751),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_876),
.A2(n_660),
.B1(n_799),
.B2(n_815),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_880),
.A2(n_836),
.B1(n_740),
.B2(n_713),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_875),
.B(n_778),
.Y(n_895)
);

OAI222xp33_ASAP7_75t_L g896 ( 
.A1(n_865),
.A2(n_717),
.B1(n_742),
.B2(n_748),
.C1(n_778),
.C2(n_772),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_873),
.A2(n_728),
.B1(n_791),
.B2(n_813),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_SL g898 ( 
.A1(n_870),
.A2(n_813),
.B1(n_708),
.B2(n_853),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_870),
.A2(n_705),
.B1(n_722),
.B2(n_772),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_866),
.A2(n_799),
.B1(n_742),
.B2(n_695),
.Y(n_900)
);

OAI22xp33_ASAP7_75t_L g901 ( 
.A1(n_871),
.A2(n_700),
.B1(n_781),
.B2(n_804),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_869),
.B(n_771),
.Y(n_902)
);

AOI221xp5_ASAP7_75t_L g903 ( 
.A1(n_874),
.A2(n_746),
.B1(n_755),
.B2(n_737),
.C(n_727),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_872),
.A2(n_804),
.B1(n_737),
.B2(n_727),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_882),
.A2(n_804),
.B1(n_696),
.B2(n_719),
.Y(n_905)
);

NAND3xp33_ASAP7_75t_L g906 ( 
.A(n_877),
.B(n_719),
.C(n_833),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_L g907 ( 
.A(n_897),
.B(n_879),
.C(n_763),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_886),
.B(n_879),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_885),
.B(n_879),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_895),
.B(n_833),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_889),
.B(n_892),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_889),
.B(n_826),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_887),
.B(n_82),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_883),
.B(n_782),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_893),
.A2(n_837),
.B1(n_788),
.B2(n_782),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_902),
.B(n_788),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_L g917 ( 
.A1(n_884),
.A2(n_878),
.B(n_88),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_898),
.B(n_891),
.C(n_899),
.Y(n_918)
);

OA21x2_ASAP7_75t_L g919 ( 
.A1(n_896),
.A2(n_837),
.B(n_93),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_890),
.B(n_91),
.Y(n_920)
);

OAI22xp33_ASAP7_75t_L g921 ( 
.A1(n_900),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_894),
.B(n_97),
.C(n_101),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_888),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_923)
);

NOR2xp67_ASAP7_75t_L g924 ( 
.A(n_906),
.B(n_113),
.Y(n_924)
);

INVxp67_ASAP7_75t_SL g925 ( 
.A(n_901),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_909),
.B(n_904),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_SL g927 ( 
.A(n_917),
.B(n_918),
.C(n_911),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_L g928 ( 
.A(n_911),
.B(n_905),
.C(n_903),
.Y(n_928)
);

AO21x2_ASAP7_75t_L g929 ( 
.A1(n_907),
.A2(n_916),
.B(n_912),
.Y(n_929)
);

AO21x2_ASAP7_75t_L g930 ( 
.A1(n_912),
.A2(n_125),
.B(n_126),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_908),
.B(n_128),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_922),
.B(n_131),
.C(n_132),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_910),
.B(n_134),
.Y(n_933)
);

NOR3xp33_ASAP7_75t_L g934 ( 
.A(n_921),
.B(n_137),
.C(n_139),
.Y(n_934)
);

INVx3_ASAP7_75t_SL g935 ( 
.A(n_913),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_925),
.B(n_146),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_935),
.B(n_919),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_929),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_926),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_930),
.Y(n_940)
);

XNOR2x2_ASAP7_75t_L g941 ( 
.A(n_927),
.B(n_915),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_931),
.B(n_919),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_930),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_936),
.Y(n_944)
);

INVx5_ASAP7_75t_L g945 ( 
.A(n_932),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_933),
.B(n_920),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_932),
.B(n_924),
.Y(n_947)
);

AO22x2_ASAP7_75t_L g948 ( 
.A1(n_928),
.A2(n_914),
.B1(n_923),
.B2(n_161),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_928),
.Y(n_949)
);

XOR2x2_ASAP7_75t_L g950 ( 
.A(n_941),
.B(n_934),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_939),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_938),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_949),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_937),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_944),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_938),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_945),
.Y(n_957)
);

XNOR2xp5_ASAP7_75t_L g958 ( 
.A(n_946),
.B(n_948),
.Y(n_958)
);

XOR2xp5_ASAP7_75t_L g959 ( 
.A(n_948),
.B(n_157),
.Y(n_959)
);

OA22x2_ASAP7_75t_L g960 ( 
.A1(n_958),
.A2(n_947),
.B1(n_943),
.B2(n_940),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_951),
.Y(n_961)
);

OA22x2_ASAP7_75t_L g962 ( 
.A1(n_959),
.A2(n_947),
.B1(n_940),
.B2(n_945),
.Y(n_962)
);

OA22x2_ASAP7_75t_SL g963 ( 
.A1(n_950),
.A2(n_945),
.B1(n_942),
.B2(n_172),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_957),
.Y(n_964)
);

OA22x2_ASAP7_75t_L g965 ( 
.A1(n_953),
.A2(n_170),
.B1(n_175),
.B2(n_176),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_952),
.Y(n_966)
);

OA22x2_ASAP7_75t_L g967 ( 
.A1(n_955),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_954),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_956),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_966),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_961),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_962),
.Y(n_972)
);

NAND4xp75_ASAP7_75t_L g973 ( 
.A(n_972),
.B(n_963),
.C(n_964),
.D(n_960),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_970),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_970),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_971),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_974),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_973),
.A2(n_965),
.B1(n_967),
.B2(n_968),
.Y(n_978)
);

AND4x1_ASAP7_75t_L g979 ( 
.A(n_976),
.B(n_969),
.C(n_966),
.D(n_188),
.Y(n_979)
);

XNOR2x1_ASAP7_75t_L g980 ( 
.A(n_978),
.B(n_975),
.Y(n_980)
);

OAI211xp5_ASAP7_75t_L g981 ( 
.A1(n_977),
.A2(n_184),
.B(n_185),
.C(n_191),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_979),
.A2(n_192),
.B1(n_198),
.B2(n_200),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_980),
.Y(n_983)
);

AND4x1_ASAP7_75t_L g984 ( 
.A(n_983),
.B(n_982),
.C(n_981),
.D(n_203),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_984),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_985),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_986),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_987),
.A2(n_201),
.B1(n_209),
.B2(n_213),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_988),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_989),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_990),
.Y(n_991)
);

OAI221xp5_ASAP7_75t_L g992 ( 
.A1(n_991),
.A2(n_232),
.B1(n_233),
.B2(n_238),
.C(n_239),
.Y(n_992)
);

AOI211xp5_ASAP7_75t_L g993 ( 
.A1(n_992),
.A2(n_247),
.B(n_254),
.C(n_256),
.Y(n_993)
);


endmodule