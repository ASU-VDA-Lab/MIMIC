module fake_jpeg_9211_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_24),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_48),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_64),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_21),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_32),
.B1(n_30),
.B2(n_33),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_56),
.A2(n_25),
.B1(n_27),
.B2(n_19),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_32),
.B1(n_22),
.B2(n_30),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_68),
.B1(n_31),
.B2(n_26),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_32),
.B1(n_33),
.B2(n_30),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_25),
.B1(n_31),
.B2(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_70),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_39),
.A2(n_33),
.B(n_15),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_16),
.B(n_17),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_26),
.B1(n_35),
.B2(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_77),
.B(n_80),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_81),
.B(n_100),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_26),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_83),
.A2(n_107),
.B(n_41),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_88),
.B1(n_93),
.B2(n_95),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_45),
.B1(n_43),
.B2(n_42),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_108),
.B1(n_72),
.B2(n_23),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_82),
.C(n_84),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_64),
.A2(n_66),
.B1(n_55),
.B2(n_68),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_41),
.C(n_21),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_57),
.A2(n_43),
.B1(n_42),
.B2(n_46),
.Y(n_95)
);

AO22x1_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_46),
.B1(n_41),
.B2(n_37),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_96),
.A2(n_115),
.B1(n_41),
.B2(n_63),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_17),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_19),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx24_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_60),
.A2(n_46),
.B1(n_41),
.B2(n_37),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_49),
.B(n_12),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_18),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_63),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_49),
.B(n_12),
.Y(n_113)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_18),
.B1(n_35),
.B2(n_23),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_95),
.C(n_115),
.Y(n_156)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_123),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_133),
.B(n_84),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_85),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_129),
.B(n_78),
.Y(n_175)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_18),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_143),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_96),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_37),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_144),
.A2(n_96),
.B(n_87),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_145),
.A2(n_110),
.B1(n_109),
.B2(n_106),
.Y(n_154)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_1),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_147),
.A2(n_149),
.B(n_130),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_144),
.A2(n_93),
.B(n_82),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_151),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_83),
.B(n_104),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_153),
.A2(n_160),
.B(n_171),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_159),
.B1(n_121),
.B2(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_161),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_166),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_90),
.B1(n_107),
.B2(n_83),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_107),
.B1(n_86),
.B2(n_101),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_165),
.B1(n_173),
.B2(n_121),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_86),
.B1(n_114),
.B2(n_79),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_79),
.C(n_99),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_1),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_170),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_168),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_136),
.Y(n_170)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_127),
.B(n_1),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_177),
.B(n_179),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_127),
.A2(n_114),
.B1(n_63),
.B2(n_99),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_134),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_116),
.A2(n_58),
.B(n_74),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_120),
.A2(n_21),
.B(n_23),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_120),
.B(n_89),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_135),
.B(n_126),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_182),
.B(n_183),
.Y(n_226)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_145),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_177),
.C(n_166),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_193),
.B1(n_200),
.B2(n_154),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_189),
.A2(n_194),
.B(n_199),
.Y(n_221)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_190),
.B(n_192),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_161),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_191),
.A2(n_209),
.B(n_130),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_122),
.B1(n_135),
.B2(n_126),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_198),
.Y(n_223)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_89),
.A3(n_34),
.B1(n_13),
.B2(n_15),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_130),
.B(n_124),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_173),
.A2(n_131),
.B1(n_78),
.B2(n_139),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_205),
.B(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_8),
.B(n_14),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g209 ( 
.A1(n_153),
.A2(n_130),
.B(n_3),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_241),
.B1(n_206),
.B2(n_209),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_219),
.Y(n_247)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_169),
.B1(n_159),
.B2(n_163),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_220),
.A2(n_222),
.B1(n_206),
.B2(n_212),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_156),
.B1(n_172),
.B2(n_147),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_224),
.Y(n_252)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_150),
.C(n_186),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_235),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_234),
.C(n_240),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_189),
.A2(n_164),
.B1(n_155),
.B2(n_158),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_233),
.B1(n_239),
.B2(n_190),
.Y(n_243)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_153),
.A3(n_149),
.B1(n_150),
.B2(n_179),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_238),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_201),
.A2(n_160),
.B1(n_166),
.B2(n_174),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_151),
.C(n_178),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_237),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_193),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_182),
.A2(n_162),
.B1(n_167),
.B2(n_157),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_167),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_215),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_194),
.B1(n_183),
.B2(n_198),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_245),
.A2(n_214),
.B1(n_219),
.B2(n_10),
.Y(n_278)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_256),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_221),
.A2(n_195),
.B(n_209),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_250),
.A2(n_263),
.B(n_2),
.Y(n_281)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_258),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_195),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_254),
.C(n_264),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_191),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_259),
.B1(n_260),
.B2(n_216),
.Y(n_273)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_222),
.A2(n_191),
.B1(n_181),
.B2(n_211),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_220),
.A2(n_181),
.B1(n_212),
.B2(n_204),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_228),
.B(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_197),
.C(n_3),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_240),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_273),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_221),
.B(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_270),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_241),
.B(n_235),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_275),
.B(n_281),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_247),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_228),
.B(n_218),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_283),
.B1(n_264),
.B2(n_243),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_224),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_279),
.C(n_282),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_214),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_2),
.C(n_3),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_R g283 ( 
.A(n_245),
.B(n_9),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_251),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_285),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_255),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_296),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_4),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_248),
.B1(n_263),
.B2(n_246),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_8),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_3),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_299),
.Y(n_310)
);

BUFx12_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_276),
.B1(n_283),
.B2(n_269),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_300),
.A2(n_302),
.B1(n_290),
.B2(n_293),
.Y(n_313)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_282),
.B(n_281),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_301),
.A2(n_287),
.B(n_285),
.Y(n_318)
);

OAI211xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_272),
.B(n_279),
.C(n_265),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_272),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_306),
.C(n_305),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_4),
.C(n_5),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_308),
.B1(n_312),
.B2(n_298),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_288),
.B(n_6),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_309),
.B(n_296),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_292),
.A2(n_6),
.B1(n_7),
.B2(n_290),
.Y(n_312)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_294),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_319),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_316),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_306),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_318),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_286),
.C(n_297),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_321),
.B(n_310),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_286),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_311),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_319),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_326),
.B(n_314),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_321),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_299),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_327),
.B(n_328),
.Y(n_335)
);

OAI211xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_325),
.B(n_334),
.C(n_322),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_298),
.B1(n_308),
.B2(n_299),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_7),
.C(n_326),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_7),
.Y(n_339)
);


endmodule