module fake_jpeg_5328_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_34),
.Y(n_48)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_46),
.Y(n_61)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_27),
.B1(n_30),
.B2(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_51),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_63),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_55),
.B1(n_44),
.B2(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_56),
.B1(n_64),
.B2(n_22),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_27),
.B1(n_30),
.B2(n_23),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_23),
.B1(n_33),
.B2(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_23),
.B1(n_33),
.B2(n_17),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_22),
.C(n_26),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_24),
.C(n_34),
.Y(n_89)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_40),
.Y(n_94)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_45),
.B1(n_37),
.B2(n_35),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_72),
.A2(n_73),
.B1(n_89),
.B2(n_75),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_41),
.B(n_38),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_76),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_82),
.Y(n_114)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_86),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_43),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_35),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_43),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_43),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_37),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_36),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_36),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_86),
.B(n_84),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_129),
.B1(n_91),
.B2(n_96),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_48),
.B(n_45),
.C(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_101),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_46),
.C(n_47),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_46),
.C(n_25),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_132),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_40),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_115),
.B(n_119),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_73),
.A2(n_62),
.B1(n_59),
.B2(n_69),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_62),
.B1(n_59),
.B2(n_69),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_85),
.A2(n_69),
.B1(n_41),
.B2(n_40),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_17),
.B1(n_29),
.B2(n_71),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_129),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_140),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_146),
.B1(n_165),
.B2(n_122),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_139),
.A2(n_155),
.B(n_25),
.Y(n_198)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_147),
.Y(n_166)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_76),
.B1(n_80),
.B2(n_102),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_150),
.B1(n_127),
.B2(n_133),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_80),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_153),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_145),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_97),
.B1(n_81),
.B2(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_81),
.B1(n_87),
.B2(n_83),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_88),
.Y(n_151)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_29),
.B1(n_82),
.B2(n_50),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_158),
.B1(n_120),
.B2(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_46),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_109),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_154),
.Y(n_200)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_161),
.Y(n_184)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_104),
.B1(n_100),
.B2(n_98),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_71),
.Y(n_159)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_50),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_126),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_164),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_115),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_111),
.A2(n_16),
.B1(n_28),
.B2(n_20),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_160),
.B1(n_142),
.B2(n_28),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_109),
.C(n_118),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_173),
.B(n_176),
.Y(n_226)
);

AOI31xp67_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_108),
.A3(n_118),
.B(n_122),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_161),
.B(n_159),
.C(n_165),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_156),
.A2(n_148),
.B(n_145),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_111),
.B1(n_118),
.B2(n_114),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_177),
.A2(n_136),
.B1(n_162),
.B2(n_137),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_133),
.B1(n_127),
.B2(n_116),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_134),
.A2(n_105),
.B1(n_114),
.B2(n_16),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_134),
.A2(n_105),
.B1(n_16),
.B2(n_95),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_191),
.B1(n_197),
.B2(n_182),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_157),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_139),
.B(n_138),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_157),
.B1(n_20),
.B2(n_10),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_25),
.B(n_32),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_198),
.B(n_199),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_16),
.B1(n_77),
.B2(n_95),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_151),
.B(n_153),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_195),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_140),
.A2(n_25),
.B(n_32),
.Y(n_195)
);

HAxp5_ASAP7_75t_SL g196 ( 
.A(n_146),
.B(n_25),
.CON(n_196),
.SN(n_196)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_32),
.B(n_28),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_28),
.B1(n_20),
.B2(n_25),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_136),
.A2(n_32),
.B(n_1),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_202),
.B(n_206),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_207),
.B1(n_183),
.B2(n_181),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_222),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_228),
.B(n_229),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

CKINVDCx12_ASAP7_75t_R g209 ( 
.A(n_174),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_211),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_214),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_20),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_191),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_216),
.B(n_218),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_217),
.Y(n_233)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_168),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_220),
.Y(n_251)
);

AO22x1_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_95),
.B1(n_77),
.B2(n_2),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_169),
.B1(n_178),
.B2(n_172),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_170),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_170),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_172),
.C(n_169),
.Y(n_238)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_77),
.B1(n_9),
.B2(n_10),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_189),
.B1(n_188),
.B2(n_194),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_192),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_230),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_173),
.C(n_185),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_236),
.C(n_252),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_192),
.C(n_190),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_238),
.A2(n_249),
.B(n_15),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_171),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_243),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_219),
.CI(n_211),
.CON(n_263),
.SN(n_263)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_166),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_196),
.C(n_193),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_248),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_0),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_201),
.B(n_195),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_201),
.A2(n_178),
.B(n_189),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_203),
.B(n_200),
.Y(n_252)
);

INVxp33_ASAP7_75t_SL g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_228),
.C(n_229),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_259),
.C(n_236),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_208),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_216),
.B1(n_204),
.B2(n_213),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_271),
.B1(n_275),
.B2(n_276),
.Y(n_278)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_221),
.C(n_214),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_261),
.B(n_262),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_205),
.C(n_213),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_239),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_224),
.B1(n_218),
.B2(n_200),
.Y(n_264)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_265),
.A2(n_274),
.B(n_249),
.Y(n_289)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_232),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_273),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_234),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_230),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_281),
.C(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_239),
.C(n_244),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_254),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_284),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_260),
.B1(n_267),
.B2(n_263),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_286),
.A2(n_12),
.B1(n_14),
.B2(n_13),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_244),
.C(n_241),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_289),
.B(n_291),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_253),
.C(n_248),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_293),
.C(n_12),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_266),
.B(n_247),
.CI(n_231),
.CON(n_291),
.SN(n_291)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_263),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_243),
.C(n_7),
.Y(n_293)
);

INVx11_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_306),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_259),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_297),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_256),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_282),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_301),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_287),
.B(n_277),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_272),
.B1(n_262),
.B2(n_275),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_266),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_297),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_276),
.B(n_12),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g308 ( 
.A1(n_304),
.A2(n_289),
.B(n_15),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_307),
.C(n_290),
.Y(n_313)
);

AO21x1_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_15),
.B(n_11),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_312),
.C(n_315),
.Y(n_328)
);

XNOR2x1_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_302),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_314),
.C(n_317),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_279),
.C(n_293),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_292),
.C(n_283),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_277),
.C(n_284),
.Y(n_319)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_312),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_320),
.A2(n_322),
.B1(n_6),
.B2(n_7),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_298),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_324),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_318),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_294),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_327),
.B(n_278),
.C(n_311),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_310),
.B(n_306),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_334),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_323),
.A2(n_316),
.B1(n_278),
.B2(n_314),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_331),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_328),
.A2(n_295),
.B1(n_310),
.B2(n_11),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_326),
.C(n_7),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_337),
.C(n_335),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_6),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_8),
.C(n_329),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_8),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_8),
.Y(n_342)
);


endmodule