module fake_netlist_6_4739_n_2199 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2199);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2199;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_2083;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_2149;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_98),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_81),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_162),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_27),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_16),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_30),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_41),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_1),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_19),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_10),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_63),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_70),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_108),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_94),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_105),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_177),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_146),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_115),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_61),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_55),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_213),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_28),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_80),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_128),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_14),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_138),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_145),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_79),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_68),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_164),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_103),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_22),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_205),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_61),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_166),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_72),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_93),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_1),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_40),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_179),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_72),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_157),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_121),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_102),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_172),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_89),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_150),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_44),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_2),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_37),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_8),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_14),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_12),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_12),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_17),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_135),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_48),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_9),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_191),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_68),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_197),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_214),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_106),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_175),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_184),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_74),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_173),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_189),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_203),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_29),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_130),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_156),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_38),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_45),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_207),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_133),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_170),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_86),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_148),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_6),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_154),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_54),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_66),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_20),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_25),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_62),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_69),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_41),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_149),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_208),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_83),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_3),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_74),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_20),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_155),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_101),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_47),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_26),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_82),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_79),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_66),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_2),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_37),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_28),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_114),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_33),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_95),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_30),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_38),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_180),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_55),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_78),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_13),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_29),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_70),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_118),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_4),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_152),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_88),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_5),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_161),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_65),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_54),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_181),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_107),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_22),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_82),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_60),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_119),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_126),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_31),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_129),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_90),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_10),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_34),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_7),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_96),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_200),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_116),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_25),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_84),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_73),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_17),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_141),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_120),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_6),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_53),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_21),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_50),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_87),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_85),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_92),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_15),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_137),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_168),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_4),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_91),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_104),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_64),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_158),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_3),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_63),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_151),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_174),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_167),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_34),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_132),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_51),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_142),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_160),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_111),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_182),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_27),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_8),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_11),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_33),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_169),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_171),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_56),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_99),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_124),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_211),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_153),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_44),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_69),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_76),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_143),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_59),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_56),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_217),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_51),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_26),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_123),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_58),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_75),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_42),
.Y(n_418)
);

BUFx10_ASAP7_75t_L g419 ( 
.A(n_59),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_48),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_190),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_195),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_144),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_39),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_18),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_40),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_206),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_39),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_198),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_228),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_326),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_269),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_281),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_283),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_291),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_386),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_307),
.B(n_0),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_285),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_287),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_374),
.B(n_0),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_300),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_333),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_232),
.B(n_5),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_333),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_293),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_307),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_232),
.B(n_246),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_333),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_294),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_329),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_307),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_299),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_333),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_251),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_301),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_333),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_333),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_311),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_251),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_355),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_324),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_312),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_333),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_318),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_389),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_332),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_338),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_347),
.Y(n_469)
);

INVxp33_ASAP7_75t_SL g470 ( 
.A(n_273),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_351),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_231),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_352),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_391),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_231),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_231),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_231),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_241),
.B(n_7),
.Y(n_478)
);

INVxp33_ASAP7_75t_SL g479 ( 
.A(n_220),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_286),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_231),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_249),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_246),
.B(n_9),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_278),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_249),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_354),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_286),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_249),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_284),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_249),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_249),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_271),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_220),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_R g494 ( 
.A(n_363),
.B(n_97),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_271),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_366),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_272),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_271),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_263),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_271),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_222),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_271),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_261),
.B(n_11),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_219),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_306),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_274),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_279),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_219),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_316),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_306),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_263),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_263),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g513 ( 
.A(n_406),
.B(n_13),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_222),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_221),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_221),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_306),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_242),
.B(n_15),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_306),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_233),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_233),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_235),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_306),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_223),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_288),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_295),
.Y(n_526)
);

INVxp33_ASAP7_75t_SL g527 ( 
.A(n_223),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_308),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_308),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_265),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_235),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_308),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_308),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g534 ( 
.A(n_265),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_308),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_304),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_240),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_337),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_305),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_240),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_438),
.B(n_261),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_431),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_501),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_472),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_472),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_475),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_475),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_438),
.B(n_422),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_448),
.B(n_337),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_437),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_499),
.B(n_337),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_514),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_445),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_437),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_511),
.B(n_337),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_437),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_437),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_445),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_532),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_447),
.B(n_337),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_436),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_476),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_437),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_462),
.A2(n_398),
.B1(n_425),
.B2(n_323),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_433),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_532),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_433),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_512),
.B(n_477),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_477),
.B(n_422),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_481),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_481),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_482),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_482),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_485),
.B(n_267),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_485),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_488),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_443),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_513),
.B(n_265),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_488),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_478),
.B(n_386),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_490),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_490),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_497),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_491),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_449),
.Y(n_588)
);

AND3x2_ASAP7_75t_L g589 ( 
.A(n_444),
.B(n_289),
.C(n_267),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_452),
.B(n_350),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_491),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_449),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_492),
.B(n_289),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_492),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_430),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_495),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_455),
.B(n_480),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_495),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_483),
.B(n_350),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_454),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_487),
.B(n_350),
.Y(n_601)
);

OAI21x1_ASAP7_75t_L g602 ( 
.A1(n_454),
.A2(n_405),
.B(n_290),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_460),
.B(n_350),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_498),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_457),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_457),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_458),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_513),
.B(n_350),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_498),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_500),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_458),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_500),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_502),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_464),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_503),
.B(n_365),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_464),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_502),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_505),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_505),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_510),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_510),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_517),
.B(n_290),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_530),
.B(n_365),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_517),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_519),
.B(n_523),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_519),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_523),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_528),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_528),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_553),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_553),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_561),
.B(n_460),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_557),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_588),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_570),
.B(n_478),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_623),
.B(n_434),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_553),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_623),
.B(n_435),
.Y(n_638)
);

AO22x2_ASAP7_75t_L g639 ( 
.A1(n_565),
.A2(n_615),
.B1(n_541),
.B2(n_548),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_553),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_L g641 ( 
.A(n_583),
.B(n_439),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_588),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_588),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_616),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_557),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_583),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_616),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_557),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_569),
.B(n_440),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_542),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_616),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_583),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_607),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_607),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_597),
.B(n_446),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_599),
.A2(n_470),
.B1(n_441),
.B2(n_413),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_599),
.A2(n_413),
.B1(n_365),
.B2(n_406),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_607),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_559),
.Y(n_659)
);

BUFx4f_ASAP7_75t_L g660 ( 
.A(n_566),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_603),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_607),
.Y(n_662)
);

AND2x2_ASAP7_75t_SL g663 ( 
.A(n_541),
.B(n_405),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_566),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_569),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_586),
.B(n_530),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_607),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_586),
.B(n_224),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_569),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_559),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_561),
.A2(n_413),
.B1(n_365),
.B2(n_518),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_568),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_557),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_542),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_551),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_568),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_557),
.Y(n_677)
);

AND2x6_ASAP7_75t_L g678 ( 
.A(n_541),
.B(n_386),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_597),
.B(n_450),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_541),
.B(n_386),
.Y(n_680)
);

INVx6_ASAP7_75t_L g681 ( 
.A(n_605),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_543),
.A2(n_534),
.B1(n_226),
.B2(n_430),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_586),
.B(n_534),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_597),
.B(n_453),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_581),
.B(n_456),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_L g686 ( 
.A1(n_543),
.A2(n_581),
.B1(n_552),
.B2(n_583),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_541),
.A2(n_540),
.B1(n_508),
.B2(n_515),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_SL g688 ( 
.A(n_565),
.B(n_516),
.C(n_504),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_568),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_548),
.B(n_459),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_559),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_569),
.B(n_463),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_559),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_568),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_569),
.B(n_465),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_561),
.B(n_467),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_590),
.B(n_529),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_577),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_557),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_560),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_548),
.B(n_468),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_590),
.B(n_469),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_560),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_SL g704 ( 
.A1(n_615),
.A2(n_518),
.B1(n_479),
.B2(n_493),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_552),
.B(n_524),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_577),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_548),
.B(n_471),
.Y(n_707)
);

BUFx4f_ASAP7_75t_L g708 ( 
.A(n_566),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_590),
.B(n_473),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_557),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_548),
.B(n_486),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_589),
.Y(n_712)
);

INVx6_ASAP7_75t_L g713 ( 
.A(n_605),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_551),
.Y(n_714)
);

INVx5_ASAP7_75t_L g715 ( 
.A(n_566),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_589),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_566),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_577),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_570),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_595),
.B(n_496),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_557),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_603),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_560),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_562),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_560),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_625),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_577),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_580),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_595),
.B(n_506),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_570),
.B(n_507),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_580),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_556),
.B(n_525),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_625),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_556),
.B(n_526),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_601),
.B(n_527),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_625),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_580),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_566),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_566),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_625),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_625),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_601),
.A2(n_413),
.B1(n_365),
.B2(n_292),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_566),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_603),
.B(n_536),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_626),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_626),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_605),
.B(n_539),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_549),
.B(n_509),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_571),
.B(n_218),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_580),
.Y(n_750)
);

BUFx4f_ASAP7_75t_L g751 ( 
.A(n_600),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_587),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_605),
.B(n_529),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_592),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_592),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_608),
.Y(n_756)
);

INVxp33_ASAP7_75t_SL g757 ( 
.A(n_549),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_608),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_626),
.Y(n_759)
);

AOI22x1_ASAP7_75t_L g760 ( 
.A1(n_571),
.A2(n_277),
.B1(n_302),
.B2(n_292),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_592),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_571),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_605),
.B(n_520),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_592),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_606),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_587),
.B(n_533),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_562),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_571),
.B(n_533),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_606),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_571),
.B(n_260),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_587),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_600),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_606),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_606),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_544),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_544),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_600),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_600),
.Y(n_778)
);

INVx4_ASAP7_75t_L g779 ( 
.A(n_600),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_587),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_627),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_627),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_SL g783 ( 
.A1(n_627),
.A2(n_489),
.B1(n_484),
.B2(n_451),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_627),
.B(n_535),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_636),
.A2(n_522),
.B1(n_531),
.B2(n_521),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_661),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_SL g787 ( 
.A1(n_724),
.A2(n_461),
.B1(n_466),
.B2(n_442),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_L g788 ( 
.A(n_646),
.B(n_386),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_675),
.B(n_600),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_714),
.B(n_600),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_661),
.Y(n_791)
);

AOI221xp5_ASAP7_75t_L g792 ( 
.A1(n_682),
.A2(n_248),
.B1(n_388),
.B2(n_381),
.C(n_378),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_646),
.B(n_600),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_652),
.B(n_611),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_665),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_735),
.B(n_474),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_722),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_652),
.B(n_611),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_719),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_756),
.B(n_611),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_663),
.A2(n_576),
.B1(n_622),
.B2(n_593),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_663),
.B(n_611),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_663),
.B(n_611),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_756),
.B(n_611),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_758),
.B(n_611),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_638),
.B(n_763),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_632),
.B(n_576),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_668),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_757),
.A2(n_537),
.B1(n_429),
.B2(n_237),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_775),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_722),
.Y(n_811)
);

INVx8_ASAP7_75t_L g812 ( 
.A(n_749),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_665),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_776),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_665),
.B(n_611),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_758),
.B(n_757),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_776),
.Y(n_817)
);

OAI22xp33_ASAP7_75t_L g818 ( 
.A1(n_668),
.A2(n_303),
.B1(n_346),
.B2(n_236),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_639),
.A2(n_576),
.B1(n_622),
.B2(n_593),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_732),
.B(n_614),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_719),
.B(n_360),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_770),
.A2(n_538),
.B(n_535),
.C(n_302),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_705),
.B(n_225),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_734),
.B(n_614),
.Y(n_824)
);

AND2x6_ASAP7_75t_SL g825 ( 
.A(n_635),
.B(n_244),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_650),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_655),
.B(n_379),
.Y(n_827)
);

NAND2x1p5_ASAP7_75t_L g828 ( 
.A(n_752),
.B(n_602),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_697),
.B(n_614),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_665),
.B(n_614),
.Y(n_830)
);

AND2x2_ASAP7_75t_SL g831 ( 
.A(n_657),
.B(n_230),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_669),
.B(n_614),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_687),
.B(n_310),
.C(n_309),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_669),
.B(n_614),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_697),
.B(n_614),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_700),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_679),
.B(n_243),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_650),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_696),
.B(n_243),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_700),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_SL g841 ( 
.A(n_716),
.B(n_413),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_702),
.B(n_247),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_703),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_669),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_709),
.B(n_614),
.Y(n_845)
);

AND2x6_ASAP7_75t_L g846 ( 
.A(n_653),
.B(n_234),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_752),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_669),
.B(n_576),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_632),
.B(n_316),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_695),
.B(n_762),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_780),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_780),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_770),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_703),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_649),
.B(n_576),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_692),
.B(n_593),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_782),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_726),
.B(n_593),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_767),
.Y(n_859)
);

NOR2xp67_ASAP7_75t_L g860 ( 
.A(n_748),
.B(n_545),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_686),
.B(n_247),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_723),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_726),
.B(n_593),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_733),
.B(n_622),
.Y(n_864)
);

AND2x6_ASAP7_75t_L g865 ( 
.A(n_653),
.B(n_245),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_733),
.B(n_622),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_736),
.B(n_622),
.Y(n_867)
);

BUFx2_ASAP7_75t_SL g868 ( 
.A(n_767),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_736),
.B(n_545),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_748),
.B(n_250),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_684),
.B(n_250),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_740),
.B(n_741),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_740),
.B(n_546),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_741),
.B(n_546),
.Y(n_874)
);

NAND3xp33_ASAP7_75t_L g875 ( 
.A(n_656),
.B(n_315),
.C(n_314),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_747),
.B(n_547),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_723),
.Y(n_877)
);

OAI22xp33_ASAP7_75t_L g878 ( 
.A1(n_716),
.A2(n_256),
.B1(n_264),
.B2(n_253),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_704),
.B(n_297),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_768),
.B(n_547),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_768),
.B(n_555),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_639),
.A2(n_258),
.B1(n_266),
.B2(n_255),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_782),
.B(n_555),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_654),
.B(n_563),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_704),
.B(n_298),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_654),
.B(n_563),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_658),
.B(n_572),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_725),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_705),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_658),
.B(n_572),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_766),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_771),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_662),
.B(n_317),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_662),
.B(n_573),
.Y(n_894)
);

OAI22xp33_ASAP7_75t_L g895 ( 
.A1(n_674),
.A2(n_340),
.B1(n_341),
.B2(n_327),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_671),
.A2(n_602),
.B(n_319),
.C(n_320),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_771),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_743),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_667),
.B(n_573),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_667),
.B(n_574),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_784),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_688),
.B(n_574),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_744),
.B(n_325),
.C(n_321),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_749),
.B(n_575),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_L g905 ( 
.A(n_641),
.B(n_330),
.C(n_328),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_781),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_749),
.B(n_575),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_725),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_745),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_681),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_690),
.B(n_255),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_781),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_639),
.A2(n_602),
.B1(n_359),
.B2(n_361),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_745),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_678),
.B(n_343),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_701),
.B(n_258),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_749),
.B(n_578),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_742),
.A2(n_407),
.B(n_320),
.C(n_319),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_753),
.B(n_578),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_707),
.B(n_336),
.C(n_334),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_711),
.B(n_266),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_746),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_639),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_666),
.B(n_316),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_746),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_681),
.B(n_579),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_712),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_683),
.B(n_322),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_681),
.B(n_579),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_635),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_660),
.A2(n_619),
.B(n_584),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_759),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_712),
.B(n_743),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_712),
.B(n_367),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_759),
.Y(n_935)
);

BUFx12f_ASAP7_75t_L g936 ( 
.A(n_635),
.Y(n_936)
);

AOI221xp5_ASAP7_75t_L g937 ( 
.A1(n_685),
.A2(n_378),
.B1(n_259),
.B2(n_257),
.C(n_252),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_681),
.B(n_582),
.Y(n_938)
);

INVx4_ASAP7_75t_L g939 ( 
.A(n_713),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_634),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_713),
.B(n_582),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_712),
.B(n_376),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_713),
.B(n_584),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_633),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_743),
.B(n_377),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_713),
.A2(n_399),
.B1(n_421),
.B2(n_427),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_720),
.B(n_268),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_738),
.B(n_739),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_738),
.B(n_585),
.Y(n_949)
);

AO221x1_ASAP7_75t_L g950 ( 
.A1(n_645),
.A2(n_296),
.B1(n_262),
.B2(n_270),
.C(n_275),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_738),
.B(n_585),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_642),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_739),
.B(n_591),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_729),
.B(n_268),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_783),
.B(n_322),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_827),
.B(n_642),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_910),
.B(n_739),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_786),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_791),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_836),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_910),
.A2(n_708),
.B(n_660),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_797),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_910),
.A2(n_708),
.B(n_660),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_806),
.B(n_643),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_944),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_853),
.B(n_643),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_853),
.B(n_644),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_889),
.Y(n_968)
);

NOR2x1_ASAP7_75t_L g969 ( 
.A(n_816),
.B(n_730),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_870),
.B(n_635),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_808),
.B(n_635),
.Y(n_971)
);

AOI21x1_ASAP7_75t_L g972 ( 
.A1(n_794),
.A2(n_647),
.B(n_644),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_939),
.A2(n_751),
.B(n_708),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_861),
.A2(n_850),
.B1(n_837),
.B2(n_939),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_826),
.B(n_777),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_939),
.A2(n_751),
.B1(n_387),
.B2(n_393),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_811),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_844),
.B(n_777),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_789),
.A2(n_751),
.B(n_717),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_844),
.B(n_777),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_849),
.B(n_322),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_790),
.A2(n_717),
.B(n_664),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_844),
.B(n_743),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_838),
.B(n_647),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_860),
.B(n_651),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_931),
.A2(n_717),
.B(n_664),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_796),
.B(n_419),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_871),
.A2(n_842),
.B(n_839),
.C(n_937),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_807),
.A2(n_678),
.B1(n_680),
.B2(n_651),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_809),
.B(n_818),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_847),
.B(n_254),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_848),
.A2(n_772),
.B(n_664),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_923),
.A2(n_676),
.B(n_689),
.C(n_672),
.Y(n_993)
);

BUFx12f_ASAP7_75t_L g994 ( 
.A(n_825),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_807),
.B(n_672),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_891),
.B(n_676),
.Y(n_996)
);

O2A1O1Ixp5_ASAP7_75t_L g997 ( 
.A1(n_876),
.A2(n_769),
.B(n_765),
.C(n_694),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_848),
.A2(n_779),
.B(n_772),
.Y(n_998)
);

AO21x1_ASAP7_75t_L g999 ( 
.A1(n_802),
.A2(n_402),
.B(n_385),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_845),
.A2(n_779),
.B(n_772),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_794),
.A2(n_694),
.B(n_689),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_847),
.B(n_276),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_901),
.B(n_698),
.Y(n_1003)
);

NAND2x1p5_ASAP7_75t_L g1004 ( 
.A(n_844),
.B(n_779),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_927),
.B(n_778),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_793),
.A2(n_778),
.B(n_743),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_836),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_812),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_855),
.B(n_698),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_856),
.B(n_706),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_868),
.B(n_419),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_802),
.A2(n_718),
.B(n_706),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_924),
.B(n_419),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_798),
.A2(n_778),
.B(n_648),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_803),
.A2(n_778),
.B(n_648),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_803),
.A2(n_727),
.B(n_718),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_872),
.A2(n_830),
.B(n_815),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_892),
.B(n_727),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_902),
.A2(n_680),
.B1(n_678),
.B2(n_773),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_892),
.B(n_728),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_927),
.B(n_280),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_859),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_815),
.A2(n_778),
.B(n_648),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_830),
.A2(n_648),
.B(n_633),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_928),
.B(n_823),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_911),
.A2(n_921),
.B(n_916),
.C(n_792),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_955),
.B(n_728),
.Y(n_1027)
);

AOI33xp33_ASAP7_75t_L g1028 ( 
.A1(n_895),
.A2(n_368),
.A3(n_282),
.B1(n_313),
.B2(n_331),
.B3(n_335),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_785),
.B(n_821),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_933),
.A2(n_680),
.B1(n_678),
.B2(n_774),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_832),
.A2(n_648),
.B(n_633),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_875),
.B(n_731),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_906),
.B(n_731),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_912),
.B(n_370),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_897),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_851),
.B(n_737),
.Y(n_1036)
);

AOI21x1_ASAP7_75t_L g1037 ( 
.A1(n_832),
.A2(n_750),
.B(n_737),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_840),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_947),
.B(n_225),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_954),
.B(n_227),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_852),
.B(n_750),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_834),
.A2(n_699),
.B(n_633),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_795),
.B(n_633),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_795),
.B(n_699),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_833),
.B(n_227),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_810),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_834),
.A2(n_710),
.B(n_699),
.Y(n_1047)
);

AOI21x1_ASAP7_75t_L g1048 ( 
.A1(n_926),
.A2(n_755),
.B(n_754),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_829),
.A2(n_755),
.B(n_754),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_857),
.B(n_831),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_929),
.A2(n_764),
.B(n_761),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_810),
.Y(n_1052)
);

OAI22x1_ASAP7_75t_L g1053 ( 
.A1(n_799),
.A2(n_229),
.B1(n_238),
.B2(n_239),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_879),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_787),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_799),
.B(n_229),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_840),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_879),
.A2(n_774),
.B(n_773),
.C(n_761),
.Y(n_1058)
);

INVxp67_ASAP7_75t_R g1059 ( 
.A(n_814),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_835),
.A2(n_896),
.B(n_828),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_843),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_831),
.B(n_764),
.Y(n_1062)
);

NOR2x2_ASAP7_75t_L g1063 ( 
.A(n_814),
.B(n_277),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_897),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_897),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_938),
.A2(n_769),
.B(n_765),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_817),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_885),
.Y(n_1068)
);

AND2x6_ASAP7_75t_L g1069 ( 
.A(n_795),
.B(n_645),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_896),
.A2(n_631),
.B(n_630),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_934),
.B(n_645),
.Y(n_1071)
);

BUFx4f_ASAP7_75t_L g1072 ( 
.A(n_936),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_820),
.A2(n_710),
.B(n_699),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_817),
.B(n_673),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_824),
.A2(n_710),
.B(n_699),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_813),
.B(n_673),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_801),
.A2(n_412),
.B1(n_760),
.B2(n_372),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_843),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_936),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_788),
.A2(n_710),
.B(n_715),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_897),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_854),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_854),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_813),
.B(n_710),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_813),
.B(n_880),
.Y(n_1085)
);

BUFx12f_ASAP7_75t_L g1086 ( 
.A(n_930),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_944),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_882),
.A2(n_407),
.B(n_428),
.C(n_420),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_L g1089 ( 
.A(n_920),
.B(n_373),
.C(n_372),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_788),
.A2(n_715),
.B(n_677),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_828),
.A2(n_631),
.B(n_630),
.Y(n_1091)
);

OR2x6_ASAP7_75t_L g1092 ( 
.A(n_812),
.B(n_375),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_858),
.A2(n_715),
.B(n_677),
.Y(n_1093)
);

AND2x6_ASAP7_75t_L g1094 ( 
.A(n_862),
.B(n_673),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_934),
.B(n_677),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_863),
.A2(n_866),
.B(n_864),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_941),
.A2(n_715),
.B(n_721),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_862),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_867),
.A2(n_907),
.B(n_904),
.Y(n_1099)
);

AOI21xp33_ASAP7_75t_L g1100 ( 
.A1(n_905),
.A2(n_342),
.B(n_339),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_944),
.B(n_721),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_881),
.B(n_721),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_940),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_877),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_943),
.A2(n_715),
.B(n_640),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_885),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_822),
.A2(n_414),
.B(n_410),
.C(n_408),
.Y(n_1107)
);

OAI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_942),
.A2(n_239),
.B(n_238),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_942),
.B(n_344),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_867),
.A2(n_715),
.B(n_640),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_933),
.A2(n_760),
.B1(n_423),
.B2(n_415),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_952),
.B(n_637),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_898),
.A2(n_659),
.B(n_637),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_877),
.B(n_693),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_888),
.B(n_693),
.Y(n_1115)
);

AO21x1_ASAP7_75t_L g1116 ( 
.A1(n_945),
.A2(n_384),
.B(n_383),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_903),
.B(n_248),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_917),
.A2(n_670),
.B(n_659),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_800),
.A2(n_691),
.B(n_670),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_L g1120 ( 
.A(n_819),
.B(n_348),
.C(n_345),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_888),
.B(n_691),
.Y(n_1121)
);

NOR3xp33_ASAP7_75t_L g1122 ( 
.A(n_878),
.B(n_380),
.C(n_373),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_909),
.Y(n_1123)
);

INVxp67_ASAP7_75t_SL g1124 ( 
.A(n_944),
.Y(n_1124)
);

NOR2x1_ASAP7_75t_L g1125 ( 
.A(n_869),
.B(n_591),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_841),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_908),
.B(n_893),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_908),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_909),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_804),
.B(n_380),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_805),
.A2(n_554),
.B(n_558),
.Y(n_1131)
);

NAND2x1p5_ASAP7_75t_L g1132 ( 
.A(n_922),
.B(n_619),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_919),
.B(n_678),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_913),
.A2(n_409),
.B1(n_415),
.B2(n_404),
.Y(n_1134)
);

OAI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_918),
.A2(n_417),
.B(n_257),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_873),
.B(n_874),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_812),
.Y(n_1137)
);

OAI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_918),
.A2(n_418),
.B(n_259),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_841),
.A2(n_390),
.B(n_397),
.C(n_396),
.Y(n_1139)
);

BUFx4f_ASAP7_75t_L g1140 ( 
.A(n_812),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_948),
.A2(n_680),
.B(n_678),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_893),
.A2(n_594),
.B(n_629),
.C(n_628),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_914),
.B(n_680),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_935),
.B(n_680),
.Y(n_1144)
);

BUFx4f_ASAP7_75t_L g1145 ( 
.A(n_846),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1136),
.B(n_883),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_968),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1008),
.B(n_935),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1086),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1026),
.B(n_988),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1026),
.A2(n_946),
.B(n_945),
.C(n_884),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_965),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_961),
.A2(n_951),
.B(n_949),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1103),
.Y(n_1154)
);

OR2x6_ASAP7_75t_SL g1155 ( 
.A(n_1134),
.B(n_1050),
.Y(n_1155)
);

NAND2xp33_ASAP7_75t_L g1156 ( 
.A(n_988),
.B(n_846),
.Y(n_1156)
);

BUFx12f_ASAP7_75t_L g1157 ( 
.A(n_994),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_963),
.A2(n_973),
.B(n_1096),
.Y(n_1158)
);

NAND2x1p5_ASAP7_75t_L g1159 ( 
.A(n_1140),
.B(n_925),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1085),
.A2(n_953),
.B(n_915),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1027),
.A2(n_886),
.B1(n_887),
.B2(n_900),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1022),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1136),
.B(n_890),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1027),
.A2(n_894),
.B1(n_899),
.B2(n_932),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1035),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_965),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_974),
.A2(n_423),
.B1(n_409),
.B2(n_404),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_965),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_956),
.B(n_846),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_1035),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_960),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_965),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1007),
.Y(n_1173)
);

AO22x1_ASAP7_75t_L g1174 ( 
.A1(n_990),
.A2(n_1029),
.B1(n_1056),
.B2(n_969),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1008),
.B(n_846),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1038),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1087),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1057),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1039),
.B(n_1040),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_990),
.B(n_349),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1064),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1029),
.A2(n_846),
.B1(n_865),
.B2(n_950),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1054),
.A2(n_915),
.B(n_403),
.C(n_400),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1073),
.A2(n_1075),
.B(n_1066),
.Y(n_1184)
);

OAI22x1_ASAP7_75t_L g1185 ( 
.A1(n_971),
.A2(n_426),
.B1(n_424),
.B2(n_418),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1087),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1068),
.A2(n_403),
.B1(n_400),
.B2(n_394),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1063),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1061),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_970),
.A2(n_865),
.B1(n_846),
.B2(n_394),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1122),
.A2(n_865),
.B1(n_680),
.B2(n_252),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_984),
.B(n_865),
.Y(n_1192)
);

CKINVDCx16_ASAP7_75t_R g1193 ( 
.A(n_1055),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_SL g1194 ( 
.A1(n_1032),
.A2(n_1060),
.B(n_1095),
.C(n_1071),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1064),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1078),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1088),
.A2(n_610),
.B(n_629),
.C(n_628),
.Y(n_1197)
);

NAND3xp33_ASAP7_75t_SL g1198 ( 
.A(n_1045),
.B(n_494),
.C(n_381),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1099),
.B(n_382),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1025),
.B(n_353),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1088),
.A2(n_609),
.B(n_624),
.C(n_621),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1106),
.B(n_382),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1011),
.B(n_392),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1087),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1082),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1083),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_984),
.B(n_865),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1065),
.Y(n_1208)
);

BUFx12f_ASAP7_75t_L g1209 ( 
.A(n_1079),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_987),
.B(n_356),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_975),
.B(n_865),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1017),
.A2(n_624),
.B(n_621),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_986),
.A2(n_1010),
.B(n_1009),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1065),
.Y(n_1214)
);

BUFx10_ASAP7_75t_L g1215 ( 
.A(n_1109),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_975),
.B(n_966),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1062),
.A2(n_392),
.B1(n_358),
.B2(n_362),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_982),
.A2(n_550),
.B(n_554),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1046),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1139),
.A2(n_620),
.B(n_594),
.C(n_618),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1013),
.B(n_357),
.Y(n_1221)
);

BUFx12f_ASAP7_75t_L g1222 ( 
.A(n_991),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1140),
.B(n_1137),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_991),
.Y(n_1224)
);

AO32x1_ASAP7_75t_L g1225 ( 
.A1(n_1077),
.A2(n_538),
.A3(n_618),
.B1(n_617),
.B2(n_613),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_971),
.A2(n_620),
.B1(n_596),
.B2(n_617),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_981),
.B(n_364),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1052),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_958),
.B(n_369),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_996),
.A2(n_371),
.B1(n_395),
.B2(n_396),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1032),
.A2(n_609),
.B(n_613),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_967),
.B(n_596),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_959),
.B(n_388),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1089),
.A2(n_598),
.B1(n_612),
.B2(n_610),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1098),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1081),
.Y(n_1236)
);

BUFx5_ASAP7_75t_L g1237 ( 
.A(n_1069),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_SL g1238 ( 
.A1(n_1005),
.A2(n_604),
.B(n_598),
.C(n_619),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1002),
.B(n_395),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_962),
.B(n_397),
.Y(n_1240)
);

O2A1O1Ixp5_ASAP7_75t_L g1241 ( 
.A1(n_999),
.A2(n_619),
.B(n_567),
.C(n_564),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1067),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_R g1243 ( 
.A(n_1137),
.B(n_401),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_R g1244 ( 
.A(n_1137),
.B(n_401),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1137),
.B(n_619),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1002),
.B(n_411),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1127),
.B(n_550),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1003),
.A2(n_426),
.B1(n_416),
.B2(n_417),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1000),
.A2(n_979),
.B(n_1004),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1104),
.Y(n_1250)
);

NOR3xp33_ASAP7_75t_SL g1251 ( 
.A(n_1108),
.B(n_411),
.C(n_416),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1128),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1089),
.A2(n_424),
.B1(n_564),
.B2(n_558),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1129),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1087),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1122),
.A2(n_567),
.B1(n_564),
.B2(n_558),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1034),
.B(n_100),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1004),
.A2(n_564),
.B(n_558),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1123),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1124),
.A2(n_1120),
.B1(n_995),
.B2(n_1133),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_977),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1127),
.Y(n_1262)
);

NAND3xp33_ASAP7_75t_SL g1263 ( 
.A(n_1109),
.B(n_16),
.C(n_18),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1126),
.B(n_19),
.Y(n_1264)
);

OAI22x1_ASAP7_75t_L g1265 ( 
.A1(n_1021),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1071),
.A2(n_564),
.B(n_558),
.C(n_554),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_R g1267 ( 
.A(n_1072),
.B(n_109),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1117),
.B(n_23),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_SL g1269 ( 
.A1(n_1095),
.A2(n_567),
.B(n_554),
.C(n_550),
.Y(n_1269)
);

NOR3xp33_ASAP7_75t_SL g1270 ( 
.A(n_1139),
.B(n_24),
.C(n_31),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1145),
.B(n_554),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1001),
.Y(n_1272)
);

OAI21xp33_ASAP7_75t_L g1273 ( 
.A1(n_1028),
.A2(n_567),
.B(n_550),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1033),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1094),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1124),
.A2(n_550),
.B1(n_567),
.B2(n_113),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1081),
.B(n_32),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1072),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_964),
.A2(n_112),
.B1(n_215),
.B2(n_212),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1094),
.Y(n_1280)
);

NOR3xp33_ASAP7_75t_SL g1281 ( 
.A(n_1135),
.B(n_1138),
.C(n_1100),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1069),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_957),
.A2(n_216),
.B(n_210),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_972),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1021),
.A2(n_209),
.B1(n_201),
.B2(n_199),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1114),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_985),
.B(n_32),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_957),
.A2(n_193),
.B(n_188),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1112),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1102),
.B(n_35),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1049),
.A2(n_187),
.B1(n_186),
.B2(n_185),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1145),
.B(n_183),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_989),
.B(n_1019),
.Y(n_1293)
);

OR2x6_ASAP7_75t_L g1294 ( 
.A(n_1092),
.B(n_178),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1043),
.A2(n_176),
.B(n_165),
.Y(n_1295)
);

AOI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1044),
.A2(n_163),
.B(n_159),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1034),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_993),
.A2(n_35),
.B(n_36),
.C(n_42),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1018),
.B(n_36),
.Y(n_1299)
);

O2A1O1Ixp5_ASAP7_75t_SL g1300 ( 
.A1(n_1130),
.A2(n_1111),
.B(n_1005),
.C(n_1044),
.Y(n_1300)
);

O2A1O1Ixp5_ASAP7_75t_L g1301 ( 
.A1(n_1130),
.A2(n_147),
.B(n_140),
.C(n_139),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1107),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1053),
.B(n_43),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1092),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1058),
.A2(n_46),
.B(n_47),
.C(n_49),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1012),
.B(n_136),
.Y(n_1306)
);

OR2x6_ASAP7_75t_SL g1307 ( 
.A(n_1020),
.B(n_49),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1016),
.B(n_134),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1115),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1294),
.B(n_1092),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1162),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1180),
.B(n_1036),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1180),
.B(n_1041),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1213),
.A2(n_1091),
.B(n_998),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1158),
.A2(n_1070),
.B(n_1037),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1179),
.B(n_1121),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1249),
.A2(n_992),
.B(n_1084),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1261),
.Y(n_1318)
);

NOR2x1_ASAP7_75t_R g1319 ( 
.A(n_1278),
.B(n_978),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1146),
.A2(n_1059),
.B1(n_1030),
.B2(n_983),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1150),
.A2(n_1298),
.B1(n_1305),
.B2(n_1302),
.C(n_1167),
.Y(n_1321)
);

BUFx12f_ASAP7_75t_L g1322 ( 
.A(n_1209),
.Y(n_1322)
);

AO21x1_ASAP7_75t_L g1323 ( 
.A1(n_1306),
.A2(n_983),
.B(n_1084),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1163),
.A2(n_1076),
.B(n_1014),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1260),
.A2(n_1116),
.A3(n_1107),
.B(n_976),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1154),
.Y(n_1326)
);

BUFx12f_ASAP7_75t_L g1327 ( 
.A(n_1222),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1300),
.A2(n_997),
.B(n_1119),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1194),
.A2(n_978),
.B(n_980),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_SL g1330 ( 
.A1(n_1296),
.A2(n_1051),
.B(n_1048),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1184),
.A2(n_1006),
.B(n_1015),
.Y(n_1331)
);

INVx8_ASAP7_75t_L g1332 ( 
.A(n_1172),
.Y(n_1332)
);

AO21x2_ASAP7_75t_L g1333 ( 
.A1(n_1194),
.A2(n_980),
.B(n_1023),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1274),
.B(n_1174),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1147),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1263),
.A2(n_1125),
.B1(n_1069),
.B2(n_1144),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1289),
.B(n_1216),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1147),
.B(n_1074),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1223),
.B(n_1101),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1156),
.A2(n_1024),
.B(n_1047),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1161),
.A2(n_1031),
.A3(n_1042),
.B(n_1093),
.Y(n_1341)
);

INVx5_ASAP7_75t_L g1342 ( 
.A(n_1172),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1164),
.A2(n_1090),
.A3(n_1105),
.B(n_1131),
.Y(n_1343)
);

AO21x2_ASAP7_75t_L g1344 ( 
.A1(n_1269),
.A2(n_1141),
.B(n_1080),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1153),
.A2(n_997),
.B(n_1097),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1281),
.A2(n_1151),
.B(n_1221),
.C(n_1210),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1200),
.B(n_1028),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_SL g1348 ( 
.A(n_1193),
.B(n_1069),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1172),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1160),
.A2(n_1118),
.B(n_1113),
.Y(n_1350)
);

AOI31xp67_ASAP7_75t_L g1351 ( 
.A1(n_1306),
.A2(n_1308),
.A3(n_1199),
.B(n_1284),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1169),
.A2(n_1308),
.B(n_1293),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1286),
.B(n_1069),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1219),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1218),
.A2(n_1110),
.B(n_1132),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1309),
.B(n_1132),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1228),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1262),
.B(n_1143),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1266),
.A2(n_1094),
.A3(n_1142),
.B(n_53),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1297),
.B(n_1094),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1293),
.A2(n_1094),
.B(n_131),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1242),
.Y(n_1362)
);

AO31x2_ASAP7_75t_L g1363 ( 
.A1(n_1272),
.A2(n_50),
.A3(n_52),
.B(n_57),
.Y(n_1363)
);

NOR2x1_ASAP7_75t_SL g1364 ( 
.A(n_1275),
.B(n_127),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1211),
.A2(n_125),
.B(n_122),
.Y(n_1365)
);

INVx3_ASAP7_75t_SL g1366 ( 
.A(n_1149),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1172),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1188),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1221),
.B(n_1200),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1157),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1175),
.A2(n_117),
.B(n_110),
.Y(n_1371)
);

AOI221x1_ASAP7_75t_L g1372 ( 
.A1(n_1291),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.C(n_60),
.Y(n_1372)
);

BUFx10_ASAP7_75t_L g1373 ( 
.A(n_1264),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1192),
.A2(n_62),
.B(n_64),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1210),
.B(n_83),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1171),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1268),
.B(n_65),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1212),
.A2(n_1258),
.B(n_1241),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1264),
.A2(n_67),
.B1(n_71),
.B2(n_73),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1227),
.B(n_67),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1281),
.A2(n_71),
.B(n_75),
.C(n_76),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1227),
.B(n_77),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1224),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1165),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1229),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_1385)
);

NOR2x1_ASAP7_75t_SL g1386 ( 
.A(n_1275),
.B(n_81),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1223),
.B(n_1304),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1241),
.A2(n_1199),
.B(n_1207),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1232),
.A2(n_1271),
.B(n_1148),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1290),
.A2(n_1182),
.B(n_1301),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_SL g1391 ( 
.A1(n_1292),
.A2(n_1183),
.B(n_1271),
.C(n_1245),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1259),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1173),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1245),
.A2(n_1282),
.B(n_1159),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1165),
.B(n_1170),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1170),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1215),
.B(n_1203),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1148),
.A2(n_1231),
.B(n_1282),
.Y(n_1398)
);

AO21x1_ASAP7_75t_L g1399 ( 
.A1(n_1287),
.A2(n_1299),
.B(n_1279),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1269),
.A2(n_1247),
.B(n_1175),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1198),
.A2(n_1202),
.B(n_1251),
.C(n_1277),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1229),
.A2(n_1233),
.B1(n_1185),
.B2(n_1257),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1176),
.Y(n_1403)
);

AO31x2_ASAP7_75t_L g1404 ( 
.A1(n_1276),
.A2(n_1225),
.A3(n_1283),
.B(n_1288),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1247),
.A2(n_1225),
.B(n_1190),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1239),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1215),
.A2(n_1244),
.B1(n_1243),
.B2(n_1303),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1225),
.A2(n_1295),
.B(n_1301),
.Y(n_1408)
);

BUFx10_ASAP7_75t_L g1409 ( 
.A(n_1233),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1178),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1177),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1181),
.B(n_1236),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1181),
.B(n_1236),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1189),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1265),
.A2(n_1235),
.A3(n_1250),
.B(n_1252),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1275),
.A2(n_1280),
.B(n_1159),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1251),
.A2(n_1217),
.B(n_1230),
.C(n_1248),
.Y(n_1417)
);

AO31x2_ASAP7_75t_L g1418 ( 
.A1(n_1196),
.A2(n_1254),
.A3(n_1206),
.B(n_1205),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1220),
.A2(n_1197),
.B(n_1201),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_SL g1420 ( 
.A(n_1243),
.B(n_1244),
.C(n_1191),
.Y(n_1420)
);

AO31x2_ASAP7_75t_L g1421 ( 
.A1(n_1187),
.A2(n_1155),
.A3(n_1238),
.B(n_1226),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1275),
.A2(n_1280),
.B(n_1257),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1280),
.A2(n_1186),
.B(n_1177),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1280),
.A2(n_1294),
.B(n_1186),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1191),
.A2(n_1253),
.B(n_1285),
.C(n_1234),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1195),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1177),
.A2(n_1186),
.B(n_1237),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1195),
.Y(n_1428)
);

INVx4_ASAP7_75t_SL g1429 ( 
.A(n_1294),
.Y(n_1429)
);

NOR4xp25_ASAP7_75t_L g1430 ( 
.A(n_1273),
.B(n_1270),
.C(n_1240),
.D(n_1246),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1177),
.A2(n_1186),
.B(n_1237),
.Y(n_1431)
);

NAND2x1p5_ASAP7_75t_L g1432 ( 
.A(n_1152),
.B(n_1166),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1208),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1270),
.A2(n_1214),
.B(n_1208),
.C(n_1256),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1214),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1267),
.A2(n_1237),
.B(n_1256),
.Y(n_1436)
);

INVx3_ASAP7_75t_SL g1437 ( 
.A(n_1152),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1166),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1237),
.A2(n_1168),
.B(n_1204),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1168),
.B(n_1204),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1255),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1255),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1267),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1307),
.B(n_1237),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1162),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1146),
.B(n_1163),
.Y(n_1446)
);

CKINVDCx11_ASAP7_75t_R g1447 ( 
.A(n_1157),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1162),
.Y(n_1448)
);

CKINVDCx6p67_ASAP7_75t_R g1449 ( 
.A(n_1209),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1180),
.B(n_1026),
.C(n_988),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1158),
.A2(n_1249),
.B(n_1184),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1146),
.B(n_1180),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1150),
.A2(n_988),
.B(n_1026),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1180),
.A2(n_1026),
.B(n_988),
.C(n_990),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1158),
.A2(n_1249),
.B(n_1184),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1150),
.A2(n_988),
.B(n_1026),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1213),
.A2(n_939),
.B(n_910),
.Y(n_1457)
);

NAND3xp33_ASAP7_75t_L g1458 ( 
.A(n_1180),
.B(n_1026),
.C(n_988),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1146),
.B(n_1180),
.Y(n_1459)
);

BUFx8_ASAP7_75t_L g1460 ( 
.A(n_1157),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1213),
.A2(n_939),
.B(n_910),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1146),
.B(n_1180),
.Y(n_1462)
);

OAI22x1_ASAP7_75t_L g1463 ( 
.A1(n_1180),
.A2(n_990),
.B1(n_1029),
.B2(n_1150),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1180),
.B(n_1026),
.C(n_988),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1158),
.A2(n_1249),
.B(n_1184),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1158),
.A2(n_1249),
.B(n_1184),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1150),
.A2(n_988),
.B(n_1026),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1180),
.A2(n_1026),
.B(n_988),
.C(n_990),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1158),
.A2(n_1249),
.B(n_1184),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1162),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1158),
.A2(n_1249),
.B(n_1184),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1180),
.A2(n_1026),
.B(n_988),
.C(n_827),
.Y(n_1472)
);

AO31x2_ASAP7_75t_L g1473 ( 
.A1(n_1158),
.A2(n_999),
.A3(n_1213),
.B(n_1260),
.Y(n_1473)
);

A2O1A1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1180),
.A2(n_1026),
.B(n_988),
.C(n_990),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1180),
.A2(n_668),
.B1(n_785),
.B2(n_821),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1180),
.A2(n_1026),
.B(n_988),
.C(n_990),
.Y(n_1476)
);

AOI221x1_ASAP7_75t_L g1477 ( 
.A1(n_1180),
.A2(n_988),
.B1(n_1026),
.B2(n_990),
.C(n_1305),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1158),
.A2(n_1249),
.B(n_1184),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1146),
.B(n_1163),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1179),
.B(n_767),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1335),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1395),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1450),
.A2(n_1458),
.B1(n_1464),
.B2(n_1475),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1326),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1452),
.B(n_1459),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1462),
.A2(n_1454),
.B1(n_1468),
.B2(n_1474),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1450),
.A2(n_1458),
.B1(n_1464),
.B2(n_1369),
.Y(n_1487)
);

BUFx10_ASAP7_75t_L g1488 ( 
.A(n_1445),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1463),
.A2(n_1420),
.B1(n_1312),
.B2(n_1313),
.Y(n_1489)
);

BUFx8_ASAP7_75t_SL g1490 ( 
.A(n_1370),
.Y(n_1490)
);

BUFx2_ASAP7_75t_SL g1491 ( 
.A(n_1470),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1311),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1447),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1375),
.A2(n_1380),
.B1(n_1382),
.B2(n_1347),
.Y(n_1494)
);

BUFx12f_ASAP7_75t_L g1495 ( 
.A(n_1460),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1318),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1342),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1476),
.A2(n_1479),
.B1(n_1446),
.B2(n_1472),
.Y(n_1498)
);

AOI21xp33_ASAP7_75t_L g1499 ( 
.A1(n_1346),
.A2(n_1456),
.B(n_1453),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1376),
.Y(n_1500)
);

INVx11_ASAP7_75t_L g1501 ( 
.A(n_1460),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1366),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1443),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1402),
.A2(n_1397),
.B1(n_1406),
.B2(n_1444),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1393),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1395),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1410),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1354),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1387),
.A2(n_1334),
.B1(n_1448),
.B2(n_1377),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1322),
.Y(n_1510)
);

CKINVDCx11_ASAP7_75t_R g1511 ( 
.A(n_1327),
.Y(n_1511)
);

INVx6_ASAP7_75t_L g1512 ( 
.A(n_1342),
.Y(n_1512)
);

NAND2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1384),
.B(n_1396),
.Y(n_1513)
);

INVx6_ASAP7_75t_L g1514 ( 
.A(n_1332),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1453),
.A2(n_1467),
.B1(n_1456),
.B2(n_1402),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1357),
.Y(n_1516)
);

INVx6_ASAP7_75t_L g1517 ( 
.A(n_1332),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1467),
.A2(n_1399),
.B1(n_1409),
.B2(n_1379),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1362),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1418),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1409),
.A2(n_1373),
.B1(n_1385),
.B2(n_1310),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1429),
.B(n_1387),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1373),
.A2(n_1385),
.B1(n_1310),
.B2(n_1480),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1477),
.A2(n_1407),
.B(n_1425),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1446),
.B(n_1479),
.Y(n_1525)
);

INVx6_ASAP7_75t_L g1526 ( 
.A(n_1349),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1448),
.A2(n_1310),
.B1(n_1348),
.B2(n_1429),
.Y(n_1527)
);

CKINVDCx11_ASAP7_75t_R g1528 ( 
.A(n_1449),
.Y(n_1528)
);

INVx6_ASAP7_75t_L g1529 ( 
.A(n_1349),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1383),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_SL g1531 ( 
.A1(n_1386),
.A2(n_1348),
.B1(n_1436),
.B2(n_1372),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1337),
.A2(n_1434),
.B1(n_1381),
.B2(n_1316),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1392),
.Y(n_1533)
);

AOI22x1_ASAP7_75t_SL g1534 ( 
.A1(n_1428),
.A2(n_1438),
.B1(n_1403),
.B2(n_1414),
.Y(n_1534)
);

CKINVDCx6p67_ASAP7_75t_R g1535 ( 
.A(n_1437),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1433),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1435),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1415),
.Y(n_1538)
);

CKINVDCx11_ASAP7_75t_R g1539 ( 
.A(n_1426),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1338),
.Y(n_1540)
);

INVx4_ASAP7_75t_L g1541 ( 
.A(n_1367),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1412),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1430),
.B(n_1321),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1413),
.Y(n_1544)
);

CKINVDCx20_ASAP7_75t_R g1545 ( 
.A(n_1368),
.Y(n_1545)
);

INVx6_ASAP7_75t_L g1546 ( 
.A(n_1367),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1430),
.B(n_1321),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1415),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1411),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_SL g1550 ( 
.A1(n_1374),
.A2(n_1339),
.B1(n_1390),
.B2(n_1336),
.Y(n_1550)
);

INVxp67_ASAP7_75t_SL g1551 ( 
.A(n_1398),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1363),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1352),
.B(n_1389),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1411),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1363),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1440),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1363),
.Y(n_1557)
);

NAND2x1p5_ASAP7_75t_L g1558 ( 
.A(n_1394),
.B(n_1360),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1390),
.A2(n_1436),
.B1(n_1323),
.B2(n_1320),
.Y(n_1559)
);

OAI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1336),
.A2(n_1356),
.B1(n_1353),
.B2(n_1320),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1360),
.A2(n_1422),
.B1(n_1358),
.B2(n_1391),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_1432),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1442),
.Y(n_1563)
);

BUFx8_ASAP7_75t_L g1564 ( 
.A(n_1319),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1358),
.A2(n_1388),
.B1(n_1361),
.B2(n_1405),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1319),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1441),
.Y(n_1567)
);

BUFx12f_ASAP7_75t_L g1568 ( 
.A(n_1371),
.Y(n_1568)
);

CKINVDCx11_ASAP7_75t_R g1569 ( 
.A(n_1424),
.Y(n_1569)
);

CKINVDCx6p67_ASAP7_75t_R g1570 ( 
.A(n_1364),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1416),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1417),
.B(n_1401),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1365),
.A2(n_1423),
.B1(n_1439),
.B2(n_1400),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1388),
.A2(n_1329),
.B1(n_1419),
.B2(n_1333),
.Y(n_1574)
);

INVx6_ASAP7_75t_L g1575 ( 
.A(n_1427),
.Y(n_1575)
);

BUFx2_ASAP7_75t_SL g1576 ( 
.A(n_1431),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1333),
.A2(n_1408),
.B1(n_1324),
.B2(n_1340),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1344),
.Y(n_1578)
);

OAI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1317),
.A2(n_1314),
.B1(n_1461),
.B2(n_1457),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1359),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1328),
.A2(n_1350),
.B1(n_1378),
.B2(n_1315),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1359),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1344),
.A2(n_1330),
.B1(n_1328),
.B2(n_1355),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1451),
.A2(n_1478),
.B1(n_1465),
.B2(n_1471),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1359),
.Y(n_1585)
);

INVx6_ASAP7_75t_L g1586 ( 
.A(n_1421),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1421),
.Y(n_1587)
);

BUFx12f_ASAP7_75t_L g1588 ( 
.A(n_1351),
.Y(n_1588)
);

BUFx12f_ASAP7_75t_L g1589 ( 
.A(n_1325),
.Y(n_1589)
);

OAI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1325),
.A2(n_1404),
.B1(n_1473),
.B2(n_1341),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1343),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1345),
.Y(n_1592)
);

CKINVDCx6p67_ASAP7_75t_R g1593 ( 
.A(n_1325),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1455),
.A2(n_1466),
.B1(n_1469),
.B2(n_1331),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1404),
.A2(n_1473),
.B1(n_1341),
.B2(n_1343),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1341),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_SL g1597 ( 
.A1(n_1404),
.A2(n_668),
.B1(n_1180),
.B2(n_990),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1343),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1473),
.A2(n_990),
.B1(n_1458),
.B2(n_1450),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1452),
.A2(n_1459),
.B1(n_1462),
.B2(n_1454),
.Y(n_1600)
);

INVx6_ASAP7_75t_L g1601 ( 
.A(n_1342),
.Y(n_1601)
);

AO22x1_ASAP7_75t_L g1602 ( 
.A1(n_1312),
.A2(n_990),
.B1(n_1180),
.B2(n_1029),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1450),
.A2(n_990),
.B1(n_1464),
.B2(n_1458),
.Y(n_1603)
);

OAI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1369),
.A2(n_668),
.B1(n_1459),
.B2(n_1452),
.Y(n_1604)
);

CKINVDCx6p67_ASAP7_75t_R g1605 ( 
.A(n_1366),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1326),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1452),
.A2(n_1459),
.B1(n_1462),
.B2(n_1454),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1450),
.A2(n_990),
.B1(n_1464),
.B2(n_1458),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1326),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1450),
.A2(n_990),
.B1(n_1464),
.B2(n_1458),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1326),
.Y(n_1611)
);

BUFx8_ASAP7_75t_L g1612 ( 
.A(n_1370),
.Y(n_1612)
);

BUFx2_ASAP7_75t_SL g1613 ( 
.A(n_1470),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_SL g1614 ( 
.A1(n_1450),
.A2(n_668),
.B1(n_1180),
.B2(n_990),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1369),
.A2(n_668),
.B1(n_1459),
.B2(n_1452),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1452),
.A2(n_1459),
.B1(n_1462),
.B2(n_1454),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1326),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1450),
.A2(n_990),
.B1(n_1464),
.B2(n_1458),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1450),
.A2(n_990),
.B1(n_1464),
.B2(n_1458),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1452),
.B(n_1459),
.Y(n_1620)
);

INVx3_ASAP7_75t_SL g1621 ( 
.A(n_1445),
.Y(n_1621)
);

OAI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1369),
.A2(n_668),
.B1(n_1459),
.B2(n_1452),
.Y(n_1622)
);

CKINVDCx11_ASAP7_75t_R g1623 ( 
.A(n_1447),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1326),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1475),
.A2(n_1180),
.B1(n_1029),
.B2(n_990),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1335),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1326),
.Y(n_1627)
);

BUFx2_ASAP7_75t_R g1628 ( 
.A(n_1445),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1450),
.A2(n_668),
.B1(n_1180),
.B2(n_990),
.Y(n_1629)
);

INVx6_ASAP7_75t_L g1630 ( 
.A(n_1342),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1335),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1452),
.B(n_1459),
.Y(n_1632)
);

BUFx10_ASAP7_75t_L g1633 ( 
.A(n_1445),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1452),
.B(n_1459),
.Y(n_1634)
);

INVx6_ASAP7_75t_L g1635 ( 
.A(n_1342),
.Y(n_1635)
);

BUFx8_ASAP7_75t_L g1636 ( 
.A(n_1370),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1326),
.Y(n_1637)
);

OAI22x1_ASAP7_75t_SL g1638 ( 
.A1(n_1443),
.A2(n_562),
.B1(n_724),
.B2(n_719),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1326),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1335),
.Y(n_1640)
);

INVx5_ASAP7_75t_L g1641 ( 
.A(n_1332),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1326),
.Y(n_1642)
);

BUFx10_ASAP7_75t_L g1643 ( 
.A(n_1445),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1452),
.A2(n_1459),
.B1(n_1462),
.B2(n_1454),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1538),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1512),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1551),
.B(n_1522),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1548),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1585),
.B(n_1515),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1614),
.A2(n_1629),
.B1(n_1625),
.B2(n_1572),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1551),
.B(n_1522),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1520),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1485),
.B(n_1620),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1552),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1575),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1591),
.B(n_1598),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1555),
.Y(n_1657)
);

AO21x2_ASAP7_75t_L g1658 ( 
.A1(n_1579),
.A2(n_1594),
.B(n_1590),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1557),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1599),
.B(n_1483),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1580),
.Y(n_1661)
);

AO21x2_ASAP7_75t_L g1662 ( 
.A1(n_1553),
.A2(n_1499),
.B(n_1592),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1569),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1485),
.B(n_1620),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1580),
.Y(n_1665)
);

OA21x2_ASAP7_75t_L g1666 ( 
.A1(n_1577),
.A2(n_1559),
.B(n_1574),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1632),
.B(n_1634),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1582),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1512),
.Y(n_1669)
);

INVx3_ASAP7_75t_SL g1670 ( 
.A(n_1535),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1602),
.B(n_1556),
.Y(n_1671)
);

NAND2x1p5_ASAP7_75t_L g1672 ( 
.A(n_1573),
.B(n_1582),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1575),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1614),
.A2(n_1629),
.B1(n_1489),
.B2(n_1523),
.Y(n_1674)
);

CKINVDCx20_ASAP7_75t_R g1675 ( 
.A(n_1623),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1575),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1558),
.Y(n_1677)
);

NAND2x1_ASAP7_75t_L g1678 ( 
.A(n_1561),
.B(n_1586),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1508),
.Y(n_1679)
);

OAI21x1_ASAP7_75t_L g1680 ( 
.A1(n_1584),
.A2(n_1553),
.B(n_1583),
.Y(n_1680)
);

INVx4_ASAP7_75t_L g1681 ( 
.A(n_1497),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1516),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1487),
.B(n_1603),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1558),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1512),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1519),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1589),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1601),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1542),
.Y(n_1689)
);

NAND2x1_ASAP7_75t_L g1690 ( 
.A(n_1586),
.B(n_1565),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1596),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1533),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_1492),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1486),
.A2(n_1509),
.B1(n_1532),
.B2(n_1607),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1632),
.B(n_1634),
.Y(n_1695)
);

AO21x1_ASAP7_75t_L g1696 ( 
.A1(n_1524),
.A2(n_1486),
.B(n_1550),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1600),
.B(n_1607),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1571),
.A2(n_1494),
.B1(n_1616),
.B2(n_1600),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1481),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1587),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1626),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1593),
.B(n_1543),
.Y(n_1702)
);

OAI21xp33_ASAP7_75t_SL g1703 ( 
.A1(n_1543),
.A2(n_1547),
.B(n_1619),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1578),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1616),
.B(n_1644),
.Y(n_1705)
);

OA21x2_ASAP7_75t_L g1706 ( 
.A1(n_1578),
.A2(n_1592),
.B(n_1547),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1609),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1499),
.A2(n_1608),
.B(n_1610),
.Y(n_1708)
);

AO21x2_ASAP7_75t_L g1709 ( 
.A1(n_1560),
.A2(n_1622),
.B(n_1615),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1644),
.B(n_1525),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1487),
.B(n_1618),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1498),
.B(n_1540),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1601),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1588),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_SL g1715 ( 
.A(n_1576),
.B(n_1498),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1544),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1497),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1611),
.Y(n_1718)
);

BUFx2_ASAP7_75t_SL g1719 ( 
.A(n_1497),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1597),
.B(n_1525),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1539),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1530),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1544),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1624),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1627),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1637),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1604),
.B(n_1536),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1639),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1642),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1484),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1532),
.B(n_1482),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1597),
.B(n_1606),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1527),
.B(n_1617),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1568),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1504),
.A2(n_1521),
.B1(n_1545),
.B2(n_1518),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1595),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1482),
.B(n_1595),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1506),
.B(n_1537),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1513),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1496),
.B(n_1505),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1500),
.B(n_1507),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1531),
.B(n_1563),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1513),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_SL g1744 ( 
.A(n_1628),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1567),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1581),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1581),
.B(n_1531),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1630),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1631),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1630),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1630),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1640),
.B(n_1613),
.Y(n_1752)
);

OAI21x1_ASAP7_75t_L g1753 ( 
.A1(n_1534),
.A2(n_1570),
.B(n_1635),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1635),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1562),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1566),
.B(n_1491),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1549),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1546),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1546),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1546),
.Y(n_1760)
);

AO21x2_ASAP7_75t_L g1761 ( 
.A1(n_1541),
.A2(n_1554),
.B(n_1526),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1529),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1564),
.B(n_1621),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1641),
.A2(n_1638),
.B(n_1517),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1514),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1517),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1628),
.B(n_1488),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1564),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1701),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1700),
.B(n_1488),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1694),
.A2(n_1503),
.B(n_1502),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1695),
.B(n_1643),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1674),
.A2(n_1605),
.B1(n_1495),
.B2(n_1510),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_L g1774 ( 
.A(n_1698),
.B(n_1636),
.C(n_1612),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1703),
.B(n_1643),
.Y(n_1775)
);

INVx4_ASAP7_75t_L g1776 ( 
.A(n_1734),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1710),
.B(n_1633),
.Y(n_1777)
);

A2O1A1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1697),
.A2(n_1493),
.B(n_1633),
.C(n_1501),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1712),
.B(n_1700),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1743),
.B(n_1528),
.Y(n_1780)
);

OAI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1735),
.A2(n_1511),
.B1(n_1612),
.B2(n_1636),
.Y(n_1781)
);

INVx4_ASAP7_75t_L g1782 ( 
.A(n_1734),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1743),
.B(n_1490),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1689),
.B(n_1742),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1732),
.B(n_1739),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1653),
.B(n_1664),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1667),
.B(n_1716),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1705),
.B(n_1712),
.Y(n_1788)
);

OA21x2_ASAP7_75t_L g1789 ( 
.A1(n_1680),
.A2(n_1746),
.B(n_1696),
.Y(n_1789)
);

AOI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1650),
.A2(n_1711),
.B1(n_1683),
.B2(n_1696),
.C(n_1660),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1683),
.A2(n_1711),
.B1(n_1660),
.B2(n_1709),
.C(n_1720),
.Y(n_1791)
);

OA21x2_ASAP7_75t_L g1792 ( 
.A1(n_1680),
.A2(n_1746),
.B(n_1657),
.Y(n_1792)
);

INVx4_ASAP7_75t_L g1793 ( 
.A(n_1734),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1723),
.B(n_1738),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1733),
.B(n_1737),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1727),
.B(n_1731),
.Y(n_1796)
);

OAI211xp5_ASAP7_75t_L g1797 ( 
.A1(n_1671),
.A2(n_1708),
.B(n_1747),
.C(n_1690),
.Y(n_1797)
);

NOR2x1_ASAP7_75t_SL g1798 ( 
.A(n_1761),
.B(n_1663),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1733),
.B(n_1737),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1733),
.B(n_1647),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1647),
.B(n_1651),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1745),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1702),
.B(n_1720),
.Y(n_1803)
);

INVx5_ASAP7_75t_SL g1804 ( 
.A(n_1734),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1675),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1702),
.B(n_1709),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1679),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1753),
.A2(n_1708),
.B(n_1752),
.Y(n_1808)
);

A2O1A1Ixp33_ASAP7_75t_L g1809 ( 
.A1(n_1678),
.A2(n_1690),
.B(n_1747),
.C(n_1753),
.Y(n_1809)
);

NAND2xp33_ASAP7_75t_R g1810 ( 
.A(n_1714),
.B(n_1708),
.Y(n_1810)
);

A2O1A1Ixp33_ASAP7_75t_L g1811 ( 
.A1(n_1678),
.A2(n_1651),
.B(n_1649),
.C(n_1764),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1651),
.B(n_1749),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_SL g1813 ( 
.A(n_1663),
.B(n_1767),
.Y(n_1813)
);

NOR2x1_ASAP7_75t_SL g1814 ( 
.A(n_1761),
.B(n_1663),
.Y(n_1814)
);

AND2x2_ASAP7_75t_SL g1815 ( 
.A(n_1708),
.B(n_1666),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1682),
.B(n_1686),
.Y(n_1816)
);

OAI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1663),
.A2(n_1756),
.B1(n_1734),
.B2(n_1699),
.Y(n_1817)
);

O2A1O1Ixp5_ASAP7_75t_L g1818 ( 
.A1(n_1714),
.A2(n_1736),
.B(n_1677),
.C(n_1684),
.Y(n_1818)
);

NOR2x1_ASAP7_75t_SL g1819 ( 
.A(n_1761),
.B(n_1663),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1709),
.B(n_1756),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1687),
.B(n_1692),
.Y(n_1821)
);

A2O1A1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1736),
.A2(n_1715),
.B(n_1714),
.C(n_1676),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1645),
.Y(n_1823)
);

OAI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1672),
.A2(n_1655),
.B(n_1676),
.Y(n_1824)
);

NOR2x1_ASAP7_75t_SL g1825 ( 
.A(n_1662),
.B(n_1658),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1707),
.B(n_1718),
.Y(n_1826)
);

OR2x6_ASAP7_75t_L g1827 ( 
.A(n_1672),
.B(n_1677),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1645),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1726),
.B(n_1704),
.Y(n_1829)
);

NAND2x1p5_ASAP7_75t_L g1830 ( 
.A(n_1677),
.B(n_1684),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1740),
.B(n_1730),
.Y(n_1831)
);

INVxp67_ASAP7_75t_L g1832 ( 
.A(n_1704),
.Y(n_1832)
);

AO32x1_ASAP7_75t_L g1833 ( 
.A1(n_1661),
.A2(n_1668),
.A3(n_1665),
.B1(n_1657),
.B2(n_1659),
.Y(n_1833)
);

CKINVDCx6p67_ASAP7_75t_R g1834 ( 
.A(n_1670),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1715),
.A2(n_1763),
.B(n_1713),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1744),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1693),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1655),
.B(n_1673),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1768),
.A2(n_1757),
.B1(n_1701),
.B2(n_1670),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1655),
.B(n_1673),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1768),
.A2(n_1670),
.B1(n_1722),
.B2(n_1721),
.Y(n_1841)
);

BUFx2_ASAP7_75t_L g1842 ( 
.A(n_1748),
.Y(n_1842)
);

INVxp67_ASAP7_75t_L g1843 ( 
.A(n_1706),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1648),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1788),
.B(n_1706),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1815),
.B(n_1662),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1815),
.B(n_1662),
.Y(n_1847)
);

OR2x6_ASAP7_75t_L g1848 ( 
.A(n_1827),
.B(n_1672),
.Y(n_1848)
);

INVxp67_ASAP7_75t_L g1849 ( 
.A(n_1820),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1807),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1795),
.B(n_1706),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1788),
.B(n_1706),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1823),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1828),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1844),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1769),
.Y(n_1856)
);

INVx5_ASAP7_75t_L g1857 ( 
.A(n_1827),
.Y(n_1857)
);

CKINVDCx20_ASAP7_75t_R g1858 ( 
.A(n_1805),
.Y(n_1858)
);

NOR2xp67_ASAP7_75t_L g1859 ( 
.A(n_1797),
.B(n_1684),
.Y(n_1859)
);

OAI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1773),
.A2(n_1666),
.B1(n_1673),
.B2(n_1676),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1792),
.B(n_1658),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1820),
.B(n_1654),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1799),
.B(n_1658),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1790),
.A2(n_1666),
.B1(n_1722),
.B2(n_1751),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1792),
.B(n_1648),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1790),
.A2(n_1666),
.B1(n_1751),
.B2(n_1750),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1792),
.B(n_1691),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1772),
.B(n_1767),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1791),
.A2(n_1774),
.B1(n_1796),
.B2(n_1797),
.Y(n_1869)
);

OAI21xp33_ASAP7_75t_L g1870 ( 
.A1(n_1791),
.A2(n_1741),
.B(n_1724),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1806),
.B(n_1725),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1832),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1806),
.B(n_1725),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1802),
.B(n_1832),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1829),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1789),
.B(n_1825),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1843),
.B(n_1652),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1812),
.Y(n_1878)
);

NAND3xp33_ASAP7_75t_L g1879 ( 
.A(n_1775),
.B(n_1729),
.C(n_1728),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1816),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1843),
.B(n_1652),
.Y(n_1881)
);

NAND3xp33_ASAP7_75t_L g1882 ( 
.A(n_1775),
.B(n_1796),
.C(n_1777),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1785),
.B(n_1803),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1826),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1801),
.B(n_1656),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1833),
.Y(n_1886)
);

HB1xp67_ASAP7_75t_L g1887 ( 
.A(n_1802),
.Y(n_1887)
);

BUFx2_ASAP7_75t_SL g1888 ( 
.A(n_1769),
.Y(n_1888)
);

AO21x2_ASAP7_75t_L g1889 ( 
.A1(n_1861),
.A2(n_1808),
.B(n_1809),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1854),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1854),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1851),
.B(n_1883),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1869),
.A2(n_1777),
.B1(n_1770),
.B2(n_1781),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1854),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1845),
.B(n_1779),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1864),
.A2(n_1809),
.B1(n_1811),
.B2(n_1786),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1865),
.Y(n_1897)
);

NAND3xp33_ASAP7_75t_L g1898 ( 
.A(n_1869),
.B(n_1882),
.C(n_1866),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1851),
.B(n_1784),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1855),
.Y(n_1900)
);

OA21x2_ASAP7_75t_L g1901 ( 
.A1(n_1886),
.A2(n_1876),
.B(n_1861),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1882),
.A2(n_1811),
.B1(n_1822),
.B2(n_1778),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1887),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1865),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1845),
.B(n_1794),
.Y(n_1905)
);

NOR3xp33_ASAP7_75t_L g1906 ( 
.A(n_1860),
.B(n_1771),
.C(n_1778),
.Y(n_1906)
);

INVx5_ASAP7_75t_L g1907 ( 
.A(n_1848),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1883),
.B(n_1800),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1852),
.B(n_1787),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1852),
.B(n_1821),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1850),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1850),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1849),
.B(n_1831),
.Y(n_1913)
);

INVxp67_ASAP7_75t_L g1914 ( 
.A(n_1871),
.Y(n_1914)
);

OAI31xp33_ASAP7_75t_SL g1915 ( 
.A1(n_1870),
.A2(n_1817),
.A3(n_1839),
.B(n_1824),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1865),
.Y(n_1916)
);

INVx2_ASAP7_75t_SL g1917 ( 
.A(n_1857),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1867),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1877),
.Y(n_1919)
);

AOI33xp33_ASAP7_75t_L g1920 ( 
.A1(n_1861),
.A2(n_1817),
.A3(n_1837),
.B1(n_1728),
.B2(n_1729),
.B3(n_1780),
.Y(n_1920)
);

BUFx2_ASAP7_75t_L g1921 ( 
.A(n_1848),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1849),
.B(n_1656),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1848),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1878),
.B(n_1798),
.Y(n_1924)
);

INVxp67_ASAP7_75t_SL g1925 ( 
.A(n_1867),
.Y(n_1925)
);

OA21x2_ASAP7_75t_L g1926 ( 
.A1(n_1886),
.A2(n_1818),
.B(n_1822),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1871),
.B(n_1814),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1881),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1873),
.B(n_1842),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1873),
.B(n_1830),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1878),
.B(n_1819),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1863),
.B(n_1818),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1868),
.B(n_1834),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1863),
.B(n_1885),
.Y(n_1934)
);

AOI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1870),
.A2(n_1841),
.B1(n_1835),
.B2(n_1836),
.C(n_1730),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1853),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1859),
.A2(n_1813),
.B1(n_1838),
.B2(n_1840),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_1856),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1936),
.Y(n_1939)
);

NOR2xp67_ASAP7_75t_L g1940 ( 
.A(n_1907),
.B(n_1857),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1936),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1890),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1932),
.B(n_1846),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1890),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1932),
.B(n_1846),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1891),
.Y(n_1946)
);

NAND4xp25_ASAP7_75t_L g1947 ( 
.A(n_1898),
.B(n_1859),
.C(n_1879),
.D(n_1810),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1901),
.B(n_1846),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1901),
.B(n_1847),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1891),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1901),
.B(n_1904),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1921),
.Y(n_1952)
);

NAND3xp33_ASAP7_75t_L g1953 ( 
.A(n_1898),
.B(n_1879),
.C(n_1810),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1894),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1914),
.B(n_1862),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1914),
.B(n_1862),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1903),
.Y(n_1957)
);

HB1xp67_ASAP7_75t_L g1958 ( 
.A(n_1930),
.Y(n_1958)
);

NAND3xp33_ASAP7_75t_L g1959 ( 
.A(n_1915),
.B(n_1847),
.C(n_1876),
.Y(n_1959)
);

INVx3_ASAP7_75t_SL g1960 ( 
.A(n_1907),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1927),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1905),
.B(n_1884),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1905),
.B(n_1884),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1901),
.B(n_1847),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1934),
.B(n_1857),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1904),
.B(n_1876),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1907),
.B(n_1857),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1897),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1897),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1894),
.Y(n_1970)
);

OAI211xp5_ASAP7_75t_SL g1971 ( 
.A1(n_1915),
.A2(n_1874),
.B(n_1872),
.C(n_1886),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1897),
.Y(n_1972)
);

NOR2x1_ASAP7_75t_L g1973 ( 
.A(n_1902),
.B(n_1888),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1916),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1900),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1919),
.B(n_1857),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1919),
.B(n_1928),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1909),
.B(n_1922),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1916),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1919),
.B(n_1857),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1928),
.B(n_1857),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1895),
.B(n_1880),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1909),
.B(n_1872),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1911),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1895),
.B(n_1880),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1910),
.B(n_1887),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1922),
.B(n_1875),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1961),
.B(n_1953),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1961),
.B(n_1920),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1953),
.B(n_1927),
.Y(n_1990)
);

BUFx2_ASAP7_75t_L g1991 ( 
.A(n_1973),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1973),
.B(n_1907),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1939),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1939),
.Y(n_1994)
);

OR3x2_ASAP7_75t_L g1995 ( 
.A(n_1947),
.B(n_1906),
.C(n_1902),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1941),
.Y(n_1996)
);

NAND2xp67_ASAP7_75t_SL g1997 ( 
.A(n_1951),
.B(n_1935),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1984),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1971),
.B(n_1858),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1957),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1984),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1978),
.B(n_1910),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1978),
.B(n_1929),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1941),
.Y(n_2004)
);

NOR2x1_ASAP7_75t_L g2005 ( 
.A(n_1947),
.B(n_1938),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1965),
.B(n_1934),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1958),
.B(n_1930),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1942),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1971),
.B(n_1933),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1955),
.B(n_1908),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1965),
.B(n_1943),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1943),
.B(n_1892),
.Y(n_2012)
);

AND2x4_ASAP7_75t_L g2013 ( 
.A(n_1940),
.B(n_1907),
.Y(n_2013)
);

NOR2xp67_ASAP7_75t_SL g2014 ( 
.A(n_1959),
.B(n_1888),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1943),
.B(n_1945),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1955),
.B(n_1956),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1952),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1945),
.B(n_1892),
.Y(n_2018)
);

INVxp67_ASAP7_75t_SL g2019 ( 
.A(n_1952),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1942),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1959),
.B(n_1935),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1986),
.B(n_1929),
.Y(n_2022)
);

NOR2x1p5_ASAP7_75t_SL g2023 ( 
.A(n_1968),
.B(n_1911),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1945),
.B(n_1921),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1962),
.B(n_1783),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1956),
.B(n_1908),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1962),
.B(n_1899),
.Y(n_2027)
);

NAND2xp67_ASAP7_75t_SL g2028 ( 
.A(n_1951),
.B(n_1981),
.Y(n_2028)
);

AND2x2_ASAP7_75t_SL g2029 ( 
.A(n_1967),
.B(n_1906),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1963),
.B(n_1899),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_1940),
.B(n_1907),
.Y(n_2031)
);

NOR2x1p5_ASAP7_75t_SL g2032 ( 
.A(n_1968),
.B(n_1912),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1944),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_1967),
.B(n_1907),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1944),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_1986),
.B(n_1983),
.Y(n_2036)
);

NOR2xp67_ASAP7_75t_L g2037 ( 
.A(n_1992),
.B(n_1981),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2021),
.B(n_1963),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1999),
.B(n_1783),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1993),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1994),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1996),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2005),
.B(n_1981),
.Y(n_2043)
);

NOR2xp67_ASAP7_75t_SL g2044 ( 
.A(n_1991),
.B(n_1719),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_2011),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2004),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1991),
.B(n_1948),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1992),
.B(n_1948),
.Y(n_2048)
);

INVx1_ASAP7_75t_SL g2049 ( 
.A(n_2029),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2008),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1992),
.B(n_1948),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2021),
.B(n_1989),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_2028),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2020),
.Y(n_2054)
);

AND2x4_ASAP7_75t_L g2055 ( 
.A(n_2019),
.B(n_1967),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_2022),
.B(n_1983),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_2017),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_2000),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_2015),
.B(n_1949),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_2022),
.B(n_1987),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2015),
.B(n_1949),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2011),
.B(n_1949),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2014),
.B(n_2012),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1990),
.B(n_1987),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2012),
.B(n_2018),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_1995),
.A2(n_1896),
.B1(n_1889),
.B2(n_1967),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2009),
.B(n_1893),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2033),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2018),
.B(n_1964),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_2003),
.B(n_1982),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_2003),
.B(n_1982),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2035),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_2013),
.B(n_1967),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2024),
.B(n_1964),
.Y(n_2074)
);

AOI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_1995),
.A2(n_1896),
.B1(n_1889),
.B2(n_1848),
.Y(n_2075)
);

OR2x6_ASAP7_75t_L g2076 ( 
.A(n_1988),
.B(n_1776),
.Y(n_2076)
);

AOI211x1_ASAP7_75t_L g2077 ( 
.A1(n_1997),
.A2(n_1964),
.B(n_1951),
.C(n_1924),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2063),
.B(n_2065),
.Y(n_2078)
);

INVxp67_ASAP7_75t_L g2079 ( 
.A(n_2057),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2063),
.B(n_2029),
.Y(n_2080)
);

AOI221x1_ASAP7_75t_L g2081 ( 
.A1(n_2052),
.A2(n_2067),
.B1(n_2055),
.B2(n_2038),
.C(n_2043),
.Y(n_2081)
);

NOR3xp33_ASAP7_75t_L g2082 ( 
.A(n_2049),
.B(n_2016),
.C(n_2025),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_2075),
.A2(n_1937),
.B1(n_1960),
.B2(n_2026),
.Y(n_2083)
);

AOI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_2066),
.A2(n_1889),
.B1(n_2034),
.B2(n_2007),
.Y(n_2084)
);

NOR2x1_ASAP7_75t_L g2085 ( 
.A(n_2076),
.B(n_2013),
.Y(n_2085)
);

O2A1O1Ixp33_ASAP7_75t_L g2086 ( 
.A1(n_2058),
.A2(n_1960),
.B(n_2036),
.C(n_2013),
.Y(n_2086)
);

INVxp67_ASAP7_75t_L g2087 ( 
.A(n_2043),
.Y(n_2087)
);

O2A1O1Ixp33_ASAP7_75t_SL g2088 ( 
.A1(n_2064),
.A2(n_2039),
.B(n_2077),
.C(n_2042),
.Y(n_2088)
);

O2A1O1Ixp33_ASAP7_75t_L g2089 ( 
.A1(n_2053),
.A2(n_1960),
.B(n_2036),
.C(n_2031),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2065),
.B(n_2024),
.Y(n_2090)
);

OAI21xp5_ASAP7_75t_SL g2091 ( 
.A1(n_2053),
.A2(n_2073),
.B(n_2047),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2042),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2046),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2045),
.B(n_2006),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2046),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2045),
.B(n_2006),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2050),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2050),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2048),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2037),
.A2(n_1889),
.B1(n_2034),
.B2(n_2031),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2055),
.A2(n_2034),
.B1(n_2031),
.B2(n_1848),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_2048),
.Y(n_2102)
);

AOI221xp5_ASAP7_75t_L g2103 ( 
.A1(n_2047),
.A2(n_1925),
.B1(n_2010),
.B2(n_2002),
.C(n_1998),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2055),
.B(n_2027),
.Y(n_2104)
);

O2A1O1Ixp33_ASAP7_75t_L g2105 ( 
.A1(n_2076),
.A2(n_1925),
.B(n_2002),
.C(n_1918),
.Y(n_2105)
);

OAI31xp33_ASAP7_75t_L g2106 ( 
.A1(n_2073),
.A2(n_1917),
.A3(n_1923),
.B(n_1976),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2054),
.Y(n_2107)
);

OAI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_2081),
.A2(n_2076),
.B1(n_2071),
.B2(n_2070),
.Y(n_2108)
);

NOR3xp33_ASAP7_75t_L g2109 ( 
.A(n_2086),
.B(n_2089),
.C(n_2091),
.Y(n_2109)
);

AOI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_2088),
.A2(n_2044),
.B1(n_2073),
.B2(n_2076),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2079),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2079),
.Y(n_2112)
);

O2A1O1Ixp33_ASAP7_75t_SL g2113 ( 
.A1(n_2087),
.A2(n_2054),
.B(n_2068),
.C(n_2072),
.Y(n_2113)
);

OAI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2084),
.A2(n_2071),
.B1(n_2070),
.B2(n_2056),
.Y(n_2114)
);

XOR2x2_ASAP7_75t_L g2115 ( 
.A(n_2080),
.B(n_2051),
.Y(n_2115)
);

O2A1O1Ixp33_ASAP7_75t_L g2116 ( 
.A1(n_2088),
.A2(n_2083),
.B(n_2087),
.C(n_2105),
.Y(n_2116)
);

NOR3xp33_ASAP7_75t_L g2117 ( 
.A(n_2082),
.B(n_2078),
.C(n_2085),
.Y(n_2117)
);

AOI221xp5_ASAP7_75t_SL g2118 ( 
.A1(n_2103),
.A2(n_2051),
.B1(n_2040),
.B2(n_2041),
.C(n_2068),
.Y(n_2118)
);

OAI22xp33_ASAP7_75t_L g2119 ( 
.A1(n_2101),
.A2(n_2060),
.B1(n_2056),
.B2(n_1923),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_L g2120 ( 
.A(n_2082),
.B(n_2060),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2092),
.B(n_2093),
.Y(n_2121)
);

AOI222xp33_ASAP7_75t_L g2122 ( 
.A1(n_2095),
.A2(n_2044),
.B1(n_2023),
.B2(n_2032),
.C1(n_2074),
.C2(n_2062),
.Y(n_2122)
);

OAI21xp33_ASAP7_75t_SL g2123 ( 
.A1(n_2106),
.A2(n_2062),
.B(n_2074),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2097),
.B(n_2098),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_R g2125 ( 
.A(n_2107),
.B(n_1766),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2099),
.B(n_2102),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_SL g2127 ( 
.A(n_2100),
.B(n_1917),
.Y(n_2127)
);

AOI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_2099),
.A2(n_1917),
.B1(n_2061),
.B2(n_2059),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2102),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_2090),
.B(n_2030),
.Y(n_2130)
);

XOR2xp5_ASAP7_75t_L g2131 ( 
.A(n_2115),
.B(n_2094),
.Y(n_2131)
);

AOI221xp5_ASAP7_75t_SL g2132 ( 
.A1(n_2116),
.A2(n_2096),
.B1(n_2104),
.B2(n_2059),
.C(n_2061),
.Y(n_2132)
);

OAI221xp5_ASAP7_75t_L g2133 ( 
.A1(n_2117),
.A2(n_2069),
.B1(n_1938),
.B2(n_2001),
.C(n_1998),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2126),
.B(n_2109),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2120),
.B(n_2069),
.Y(n_2135)
);

BUFx3_ASAP7_75t_L g2136 ( 
.A(n_2111),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2129),
.Y(n_2137)
);

AOI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_2108),
.A2(n_2001),
.B(n_1918),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2112),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2118),
.B(n_1966),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2121),
.Y(n_2141)
);

AOI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_2113),
.A2(n_1984),
.B(n_1950),
.Y(n_2142)
);

AOI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_2110),
.A2(n_1924),
.B1(n_1931),
.B2(n_1976),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2114),
.A2(n_1931),
.B1(n_1976),
.B2(n_1980),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2121),
.Y(n_2145)
);

A2O1A1Ixp33_ASAP7_75t_L g2146 ( 
.A1(n_2123),
.A2(n_2127),
.B(n_2124),
.C(n_2128),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2138),
.A2(n_2119),
.B(n_2124),
.Y(n_2147)
);

AOI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_2131),
.A2(n_2122),
.B(n_2130),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2134),
.B(n_2125),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_2136),
.Y(n_2150)
);

AOI21xp5_ASAP7_75t_L g2151 ( 
.A1(n_2146),
.A2(n_1950),
.B(n_1946),
.Y(n_2151)
);

OAI211xp5_ASAP7_75t_SL g2152 ( 
.A1(n_2133),
.A2(n_1913),
.B(n_1985),
.C(n_1762),
.Y(n_2152)
);

NAND3xp33_ASAP7_75t_L g2153 ( 
.A(n_2132),
.B(n_1755),
.C(n_1758),
.Y(n_2153)
);

NAND4xp25_ASAP7_75t_L g2154 ( 
.A(n_2135),
.B(n_1782),
.C(n_1793),
.D(n_1776),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2135),
.B(n_1980),
.Y(n_2155)
);

OA211x2_ASAP7_75t_L g2156 ( 
.A1(n_2140),
.A2(n_2032),
.B(n_2023),
.C(n_1874),
.Y(n_2156)
);

NAND4xp25_ASAP7_75t_L g2157 ( 
.A(n_2143),
.B(n_1793),
.C(n_1782),
.D(n_1938),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_2144),
.B(n_1856),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2139),
.B(n_1980),
.Y(n_2159)
);

NOR3xp33_ASAP7_75t_L g2160 ( 
.A(n_2150),
.B(n_2137),
.C(n_2141),
.Y(n_2160)
);

O2A1O1Ixp33_ASAP7_75t_L g2161 ( 
.A1(n_2147),
.A2(n_2145),
.B(n_2140),
.C(n_2142),
.Y(n_2161)
);

NAND4xp25_ASAP7_75t_L g2162 ( 
.A(n_2148),
.B(n_1856),
.C(n_1966),
.D(n_1838),
.Y(n_2162)
);

O2A1O1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_2149),
.A2(n_2151),
.B(n_2158),
.C(n_2159),
.Y(n_2163)
);

NAND2xp33_ASAP7_75t_L g2164 ( 
.A(n_2155),
.B(n_1966),
.Y(n_2164)
);

AOI321xp33_ASAP7_75t_L g2165 ( 
.A1(n_2156),
.A2(n_1840),
.A3(n_1977),
.B1(n_1754),
.B2(n_1760),
.C(n_1758),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2157),
.A2(n_1926),
.B1(n_1848),
.B2(n_1804),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_R g2167 ( 
.A(n_2154),
.B(n_1766),
.Y(n_2167)
);

HB1xp67_ASAP7_75t_L g2168 ( 
.A(n_2160),
.Y(n_2168)
);

NAND3xp33_ASAP7_75t_L g2169 ( 
.A(n_2161),
.B(n_2153),
.C(n_2152),
.Y(n_2169)
);

OAI211xp5_ASAP7_75t_L g2170 ( 
.A1(n_2163),
.A2(n_1681),
.B(n_1926),
.C(n_1717),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2164),
.Y(n_2171)
);

NOR3xp33_ASAP7_75t_L g2172 ( 
.A(n_2162),
.B(n_1766),
.C(n_1681),
.Y(n_2172)
);

OAI22x1_ASAP7_75t_L g2173 ( 
.A1(n_2166),
.A2(n_1974),
.B1(n_1968),
.B2(n_1969),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_R g2174 ( 
.A(n_2167),
.B(n_2165),
.Y(n_2174)
);

AOI221xp5_ASAP7_75t_L g2175 ( 
.A1(n_2161),
.A2(n_1954),
.B1(n_1946),
.B2(n_1970),
.C(n_1975),
.Y(n_2175)
);

AOI211xp5_ASAP7_75t_L g2176 ( 
.A1(n_2161),
.A2(n_1760),
.B(n_1759),
.C(n_1977),
.Y(n_2176)
);

XNOR2x1_ASAP7_75t_L g2177 ( 
.A(n_2168),
.B(n_1719),
.Y(n_2177)
);

INVx1_ASAP7_75t_SL g2178 ( 
.A(n_2174),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_2171),
.A2(n_2172),
.B1(n_2169),
.B2(n_2170),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2176),
.Y(n_2180)
);

INVx1_ASAP7_75t_SL g2181 ( 
.A(n_2173),
.Y(n_2181)
);

NAND4xp75_ASAP7_75t_L g2182 ( 
.A(n_2175),
.B(n_1926),
.C(n_1646),
.D(n_1688),
.Y(n_2182)
);

XNOR2x1_ASAP7_75t_L g2183 ( 
.A(n_2168),
.B(n_1926),
.Y(n_2183)
);

NAND3xp33_ASAP7_75t_L g2184 ( 
.A(n_2179),
.B(n_1681),
.C(n_1759),
.Y(n_2184)
);

INVxp67_ASAP7_75t_L g2185 ( 
.A(n_2177),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2178),
.B(n_1954),
.Y(n_2186)
);

HB1xp67_ASAP7_75t_L g2187 ( 
.A(n_2185),
.Y(n_2187)
);

OAI22x1_ASAP7_75t_L g2188 ( 
.A1(n_2187),
.A2(n_2181),
.B1(n_2180),
.B2(n_2184),
.Y(n_2188)
);

OAI22x1_ASAP7_75t_L g2189 ( 
.A1(n_2188),
.A2(n_2186),
.B1(n_2183),
.B2(n_2182),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_2188),
.B(n_1969),
.Y(n_2190)
);

AOI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2189),
.A2(n_2190),
.B1(n_1977),
.B2(n_1979),
.Y(n_2191)
);

XNOR2xp5_ASAP7_75t_L g2192 ( 
.A(n_2189),
.B(n_1646),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2192),
.Y(n_2193)
);

OAI22xp5_ASAP7_75t_SL g2194 ( 
.A1(n_2191),
.A2(n_1713),
.B1(n_1669),
.B2(n_1685),
.Y(n_2194)
);

AOI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_2193),
.A2(n_1972),
.B1(n_1974),
.B2(n_1979),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2195),
.A2(n_2194),
.B1(n_1969),
.B2(n_1972),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2196),
.Y(n_2197)
);

OAI221xp5_ASAP7_75t_R g2198 ( 
.A1(n_2197),
.A2(n_1804),
.B1(n_1979),
.B2(n_1972),
.C(n_1974),
.Y(n_2198)
);

AOI211xp5_ASAP7_75t_L g2199 ( 
.A1(n_2198),
.A2(n_1717),
.B(n_1765),
.C(n_1748),
.Y(n_2199)
);


endmodule