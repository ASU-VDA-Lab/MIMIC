module fake_jpeg_28829_n_176 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_4),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_75),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_59),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_70),
.Y(n_96)
);

CKINVDCx6p67_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_81),
.Y(n_83)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_92),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_59),
.B1(n_69),
.B2(n_61),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_93),
.B1(n_95),
.B2(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_60),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_69),
.B1(n_61),
.B2(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_79),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_61),
.B1(n_70),
.B2(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_2),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_65),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_102),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_82),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_79),
.B(n_57),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_115),
.B(n_116),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_74),
.B1(n_67),
.B2(n_58),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_86),
.B1(n_3),
.B2(n_5),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_107),
.Y(n_124)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_52),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_55),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_9),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_114),
.B(n_87),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_79),
.B(n_71),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_66),
.B(n_64),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_131),
.Y(n_141)
);

NAND2xp67_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_26),
.Y(n_119)
);

NOR4xp25_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_15),
.C(n_16),
.D(n_17),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_136),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_63),
.B(n_86),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_105),
.C(n_31),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_130),
.B1(n_137),
.B2(n_13),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_139),
.B(n_11),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_8),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_134),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_8),
.Y(n_134)
);

OAI32xp33_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_29),
.A3(n_47),
.B1(n_46),
.B2(n_45),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_16),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_104),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_30),
.B(n_43),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_13),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_148),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_149),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_128),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_27),
.C(n_42),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_48),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_14),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_25),
.C(n_38),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_19),
.B(n_23),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_153),
.B(n_154),
.C(n_156),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_15),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_150),
.A2(n_139),
.B(n_119),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_155),
.B1(n_35),
.B2(n_37),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_152),
.B1(n_149),
.B2(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

OAI321xp33_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_135),
.A3(n_145),
.B1(n_142),
.B2(n_122),
.C(n_147),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_168),
.B(n_158),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_165),
.C(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_160),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_170),
.A3(n_163),
.B1(n_161),
.B2(n_41),
.C1(n_32),
.C2(n_129),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_129),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_163),
.C(n_133),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_133),
.Y(n_176)
);


endmodule