module fake_jpeg_14266_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_4),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_14),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_22),
.Y(n_25)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_4),
.B1(n_2),
.B2(n_0),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_19),
.B1(n_20),
.B2(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_21),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_6),
.A2(n_0),
.B1(n_2),
.B2(n_12),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_9),
.B(n_11),
.C(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_26),
.B1(n_19),
.B2(n_20),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_6),
.B1(n_13),
.B2(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_23),
.B1(n_27),
.B2(n_25),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_25),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_26),
.C(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_34),
.A2(n_24),
.B1(n_21),
.B2(n_31),
.Y(n_38)
);

AOI21x1_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_39),
.B(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_16),
.B1(n_22),
.B2(n_35),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_40),
.C(n_37),
.Y(n_43)
);

A2O1A1O1Ixp25_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_36),
.B(n_33),
.C(n_16),
.D(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_42),
.Y(n_46)
);


endmodule