module fake_jpeg_345_n_676 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_676);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_676;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_13),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_62),
.Y(n_154)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_27),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_65),
.B(n_68),
.Y(n_165)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_16),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_70),
.Y(n_198)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_71),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_73),
.B(n_86),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_74),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx12f_ASAP7_75t_SL g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_76),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_81),
.Y(n_190)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_16),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_85),
.B(n_87),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_18),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_88),
.Y(n_188)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_26),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_91),
.B(n_97),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_92),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_58),
.B(n_15),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_98),
.B(n_99),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_21),
.B(n_15),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_100),
.B(n_105),
.Y(n_180)
);

BUFx16f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_101),
.Y(n_212)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_104),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_37),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_30),
.B(n_13),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_108),
.B(n_121),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_33),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_37),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_116),
.B(n_128),
.Y(n_186)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_34),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_22),
.B(n_0),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_123),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_49),
.B(n_2),
.Y(n_121)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_22),
.Y(n_123)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_123),
.Y(n_211)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_34),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_34),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_127),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_37),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_35),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_130),
.Y(n_220)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_59),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_76),
.A2(n_56),
.B1(n_38),
.B2(n_53),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_146),
.B(n_189),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_101),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_147),
.B(n_151),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_64),
.B(n_56),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_81),
.B(n_25),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_160),
.B(n_161),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_94),
.B(n_57),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_106),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_162),
.B(n_166),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_163),
.B(n_104),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_61),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_171),
.B(n_172),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_72),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_95),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_173),
.B(n_187),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_57),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_175),
.B(n_176),
.C(n_183),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_88),
.B(n_53),
.C(n_43),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_82),
.A2(n_21),
.B(n_51),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_109),
.A2(n_24),
.B1(n_51),
.B2(n_50),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_184),
.A2(n_194),
.B1(n_199),
.B2(n_221),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_114),
.A2(n_42),
.B1(n_35),
.B2(n_45),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_89),
.B(n_90),
.C(n_71),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_192),
.B(n_208),
.C(n_107),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_77),
.B(n_59),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_203),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_70),
.A2(n_50),
.B1(n_45),
.B2(n_32),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_213),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_75),
.B(n_32),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_197),
.B(n_207),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_125),
.A2(n_31),
.B1(n_25),
.B2(n_24),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_77),
.B(n_31),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_96),
.B(n_42),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_92),
.B(n_2),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_130),
.B(n_42),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_146),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_110),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_110),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_126),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_92),
.B(n_2),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_104),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_119),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_221)
);

BUFx12_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_224),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_138),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_225),
.Y(n_316)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

INVx11_ASAP7_75t_L g346 ( 
.A(n_227),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_138),
.Y(n_230)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_230),
.Y(n_338)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

NAND3xp33_ASAP7_75t_L g323 ( 
.A(n_234),
.B(n_251),
.C(n_252),
.Y(n_323)
);

CKINVDCx9p33_ASAP7_75t_R g235 ( 
.A(n_132),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_235),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_179),
.A2(n_118),
.B1(n_122),
.B2(n_78),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_238),
.A2(n_259),
.B1(n_260),
.B2(n_280),
.Y(n_337)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_239),
.Y(n_333)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_241),
.Y(n_331)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_134),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_242),
.Y(n_362)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_164),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_243),
.Y(n_343)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_134),
.Y(n_244)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_244),
.Y(n_319)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_174),
.Y(n_245)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_245),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_SL g246 ( 
.A(n_200),
.B(n_83),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_246),
.B(n_295),
.Y(n_349)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_247),
.Y(n_314)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_249),
.Y(n_348)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_250),
.Y(n_336)
);

CKINVDCx12_ASAP7_75t_R g252 ( 
.A(n_154),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_142),
.Y(n_253)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_254),
.B(n_267),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_255),
.B(n_289),
.Y(n_328)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_256),
.Y(n_341)
);

INVx6_ASAP7_75t_SL g258 ( 
.A(n_132),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_258),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_175),
.A2(n_69),
.B1(n_102),
.B2(n_8),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_206),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_159),
.Y(n_261)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_186),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_262),
.B(n_264),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_144),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_180),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_133),
.Y(n_265)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_132),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_191),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_268),
.B(n_293),
.Y(n_356)
);

CKINVDCx12_ASAP7_75t_R g269 ( 
.A(n_154),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_269),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_209),
.B(n_4),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_270),
.B(n_279),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_145),
.B(n_126),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_271),
.B(n_275),
.Y(n_353)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_155),
.Y(n_272)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_141),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_163),
.A2(n_93),
.B1(n_9),
.B2(n_10),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_274),
.A2(n_222),
.B1(n_204),
.B2(n_148),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_181),
.B(n_93),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_153),
.Y(n_276)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_153),
.Y(n_277)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_277),
.Y(n_320)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_185),
.Y(n_278)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_165),
.B(n_7),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_194),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_280)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_144),
.Y(n_281)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_159),
.Y(n_282)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_282),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_215),
.B(n_11),
.C(n_12),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_283),
.B(n_143),
.C(n_201),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_183),
.A2(n_11),
.B1(n_12),
.B2(n_158),
.Y(n_284)
);

AOI22x1_ASAP7_75t_L g310 ( 
.A1(n_284),
.A2(n_201),
.B1(n_198),
.B2(n_141),
.Y(n_310)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_285),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_167),
.Y(n_286)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_286),
.Y(n_327)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_190),
.Y(n_287)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_137),
.A2(n_11),
.B1(n_12),
.B2(n_140),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_288),
.A2(n_218),
.B1(n_202),
.B2(n_168),
.Y(n_347)
);

BUFx12f_ASAP7_75t_L g289 ( 
.A(n_223),
.Y(n_289)
);

INVx13_ASAP7_75t_SL g291 ( 
.A(n_189),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_291),
.A2(n_294),
.B1(n_299),
.B2(n_301),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_139),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g294 ( 
.A(n_223),
.Y(n_294)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_139),
.Y(n_295)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_167),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_296),
.B(n_297),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_211),
.B(n_149),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_150),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_156),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_170),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_149),
.B(n_208),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_300),
.B(n_297),
.Y(n_363)
);

INVx5_ASAP7_75t_SL g301 ( 
.A(n_218),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_135),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_302),
.A2(n_152),
.B1(n_168),
.B2(n_191),
.Y(n_330)
);

OR2x4_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_189),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_309),
.B(n_260),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_310),
.B(n_329),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_228),
.A2(n_157),
.B1(n_158),
.B2(n_170),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_311),
.A2(n_335),
.B1(n_347),
.B2(n_301),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_325),
.B(n_357),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_248),
.B(n_176),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_284),
.B(n_192),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_226),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_228),
.A2(n_202),
.B1(n_174),
.B2(n_198),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_268),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_233),
.A2(n_152),
.B1(n_135),
.B2(n_188),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_354),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_254),
.A2(n_152),
.B1(n_188),
.B2(n_136),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_300),
.B(n_136),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_247),
.C(n_302),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_234),
.A2(n_219),
.B1(n_178),
.B2(n_220),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_360),
.A2(n_312),
.B1(n_357),
.B2(n_309),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_273),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_257),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_364),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_325),
.B(n_292),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_365),
.B(n_372),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_366),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_316),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_367),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_368),
.B(n_380),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_369),
.A2(n_378),
.B1(n_385),
.B2(n_377),
.Y(n_417)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_371),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_340),
.B(n_353),
.Y(n_372)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_326),
.B(n_290),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_374),
.Y(n_416)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_334),
.Y(n_375)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_375),
.Y(n_426)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_332),
.A2(n_232),
.B1(n_229),
.B2(n_288),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_376),
.A2(n_402),
.B1(n_403),
.B2(n_406),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_307),
.A2(n_360),
.B1(n_349),
.B2(n_310),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_308),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_379),
.A2(n_401),
.B1(n_342),
.B2(n_333),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_304),
.B(n_236),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_349),
.A2(n_237),
.B(n_243),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_383),
.A2(n_322),
.B(n_355),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_384),
.B(n_400),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_306),
.Y(n_418)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_314),
.Y(n_386)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_386),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_348),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_387),
.B(n_396),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_389),
.B(n_394),
.Y(n_428)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_334),
.Y(n_390)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_390),
.Y(n_440)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_314),
.Y(n_391)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_323),
.B(n_307),
.Y(n_392)
);

BUFx12_ASAP7_75t_L g431 ( 
.A(n_392),
.Y(n_431)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_393),
.Y(n_448)
);

OR2x2_ASAP7_75t_SL g394 ( 
.A(n_363),
.B(n_287),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_395),
.B(n_397),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_305),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_356),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_399),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_249),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_315),
.B(n_250),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_335),
.A2(n_266),
.B1(n_265),
.B2(n_227),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_310),
.A2(n_282),
.B1(n_261),
.B2(n_299),
.Y(n_402)
);

OAI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_328),
.A2(n_311),
.B1(n_337),
.B2(n_361),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_404),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_307),
.B(n_295),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_407),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_343),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_342),
.B(n_148),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_343),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_409),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_350),
.B(n_244),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_333),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_411),
.Y(n_432)
);

OR2x2_ASAP7_75t_SL g411 ( 
.A(n_351),
.B(n_231),
.Y(n_411)
);

AO21x1_ASAP7_75t_L g465 ( 
.A1(n_417),
.A2(n_394),
.B(n_381),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_418),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_369),
.A2(n_318),
.B1(n_306),
.B2(n_327),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_425),
.A2(n_437),
.B1(n_386),
.B2(n_393),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_427),
.A2(n_436),
.B(n_443),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_377),
.A2(n_318),
.B1(n_245),
.B2(n_281),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_429),
.A2(n_438),
.B1(n_446),
.B2(n_447),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_370),
.A2(n_322),
.B(n_355),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_378),
.A2(n_327),
.B1(n_308),
.B2(n_338),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_384),
.A2(n_296),
.B1(n_225),
.B2(n_286),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_399),
.B(n_388),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_441),
.Y(n_459)
);

OAI32xp33_ASAP7_75t_L g441 ( 
.A1(n_371),
.A2(n_313),
.A3(n_344),
.B1(n_352),
.B2(n_317),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_364),
.B(n_395),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_445),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_370),
.A2(n_362),
.B(n_303),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_389),
.B(n_305),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_366),
.A2(n_411),
.B1(n_405),
.B2(n_383),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_381),
.A2(n_230),
.B1(n_263),
.B2(n_316),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_415),
.B(n_372),
.Y(n_452)
);

NAND3xp33_ASAP7_75t_L g518 ( 
.A(n_452),
.B(n_461),
.C(n_486),
.Y(n_518)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_453),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_398),
.Y(n_454)
);

NOR2x1_ASAP7_75t_L g512 ( 
.A(n_454),
.B(n_476),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_430),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_455),
.B(n_458),
.Y(n_510)
);

INVx13_ASAP7_75t_L g456 ( 
.A(n_420),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_456),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_430),
.Y(n_458)
);

INVx3_ASAP7_75t_SL g460 ( 
.A(n_413),
.Y(n_460)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_460),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_416),
.B(n_365),
.Y(n_461)
);

INVx3_ASAP7_75t_SL g463 ( 
.A(n_450),
.Y(n_463)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_463),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_387),
.Y(n_464)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_464),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_465),
.B(n_469),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_418),
.A2(n_382),
.B(n_404),
.Y(n_466)
);

OA21x2_ASAP7_75t_L g507 ( 
.A1(n_466),
.A2(n_418),
.B(n_436),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_421),
.B(n_324),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_467),
.B(n_472),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_431),
.B(n_392),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_481),
.Y(n_493)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_435),
.Y(n_471)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_471),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_421),
.B(n_320),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_417),
.A2(n_382),
.B1(n_396),
.B2(n_391),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_473),
.A2(n_469),
.B1(n_429),
.B2(n_460),
.Y(n_497)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_448),
.Y(n_475)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_475),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_427),
.B(n_407),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_412),
.B(n_397),
.Y(n_477)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_477),
.Y(n_524)
);

AND2x2_ASAP7_75t_SL g478 ( 
.A(n_428),
.B(n_390),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_478),
.Y(n_504)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_414),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_480),
.Y(n_489)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_414),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_444),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_482),
.B(n_488),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_442),
.B(n_321),
.C(n_336),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_484),
.C(n_445),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_428),
.B(n_341),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_319),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_419),
.B(n_341),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_449),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_434),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_492),
.B(n_498),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_459),
.A2(n_457),
.B1(n_488),
.B2(n_463),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_496),
.A2(n_523),
.B1(n_476),
.B2(n_465),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_497),
.A2(n_522),
.B1(n_474),
.B2(n_466),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_449),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_499),
.B(n_506),
.C(n_513),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_464),
.B(n_434),
.Y(n_501)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_501),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_483),
.B(n_422),
.C(n_432),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_507),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_459),
.B(n_451),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_509),
.B(n_511),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_454),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_462),
.B(n_422),
.C(n_432),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_484),
.B(n_439),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_514),
.B(n_478),
.Y(n_537)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_479),
.Y(n_515)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_515),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_425),
.Y(n_516)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_516),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_487),
.B(n_415),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_517),
.B(n_519),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_454),
.B(n_424),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_453),
.B(n_424),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_521),
.B(n_471),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_457),
.A2(n_437),
.B1(n_438),
.B2(n_443),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_474),
.A2(n_446),
.B1(n_418),
.B2(n_431),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_526),
.A2(n_531),
.B1(n_534),
.B2(n_549),
.Y(n_567)
);

INVxp33_ASAP7_75t_SL g527 ( 
.A(n_493),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_527),
.B(n_544),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_481),
.Y(n_529)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_529),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_502),
.B(n_475),
.Y(n_530)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_530),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_SL g533 ( 
.A(n_523),
.B(n_485),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_533),
.A2(n_542),
.B(n_551),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_496),
.A2(n_470),
.B1(n_473),
.B2(n_418),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_536),
.A2(n_508),
.B1(n_504),
.B2(n_524),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_537),
.B(n_545),
.Y(n_558)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_495),
.Y(n_539)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_539),
.Y(n_568)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_495),
.Y(n_540)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_540),
.Y(n_570)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_501),
.Y(n_541)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_541),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_512),
.A2(n_485),
.B(n_476),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_520),
.B(n_480),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_499),
.B(n_478),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_SL g546 ( 
.A(n_493),
.B(n_468),
.C(n_431),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_546),
.B(n_507),
.C(n_536),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_510),
.B(n_516),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_547),
.B(n_548),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_489),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_503),
.A2(n_470),
.B1(n_482),
.B2(n_456),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_505),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_550),
.B(n_554),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_512),
.A2(n_431),
.B(n_447),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_503),
.A2(n_433),
.B1(n_444),
.B2(n_440),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_553),
.A2(n_494),
.B1(n_515),
.B2(n_426),
.Y(n_577)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_505),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_524),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_555),
.B(n_557),
.Y(n_581)
);

NOR2x1p5_ASAP7_75t_SL g557 ( 
.A(n_508),
.B(n_441),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_549),
.Y(n_559)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_559),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_529),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_560),
.B(n_564),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_561),
.B(n_569),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_532),
.B(n_492),
.C(n_498),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_565),
.A2(n_573),
.B1(n_580),
.B2(n_552),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_532),
.B(n_506),
.C(n_514),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_566),
.B(n_572),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_543),
.B(n_513),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_543),
.B(n_508),
.C(n_507),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_534),
.A2(n_497),
.B1(n_494),
.B2(n_491),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_545),
.B(n_491),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_574),
.B(n_533),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_537),
.B(n_500),
.C(n_490),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_575),
.B(n_582),
.C(n_553),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_577),
.A2(n_552),
.B1(n_551),
.B2(n_542),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_528),
.A2(n_518),
.B1(n_440),
.B2(n_426),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_546),
.B(n_375),
.C(n_319),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_530),
.B(n_379),
.Y(n_584)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_584),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_587),
.B(n_597),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_588),
.A2(n_593),
.B1(n_563),
.B2(n_562),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_589),
.B(n_605),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_566),
.B(n_556),
.C(n_538),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_591),
.B(n_599),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_567),
.A2(n_525),
.B1(n_547),
.B2(n_557),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_584),
.Y(n_594)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_594),
.Y(n_613)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_579),
.Y(n_595)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_595),
.Y(n_615)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_576),
.Y(n_596)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_596),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_578),
.Y(n_598)
);

NOR3xp33_ASAP7_75t_L g612 ( 
.A(n_598),
.B(n_600),
.C(n_602),
.Y(n_612)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_581),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_581),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_SL g601 ( 
.A(n_558),
.B(n_572),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_601),
.B(n_561),
.Y(n_624)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_580),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_565),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_603),
.B(n_568),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_564),
.B(n_535),
.C(n_379),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_605),
.B(n_575),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_583),
.A2(n_535),
.B(n_336),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_606),
.A2(n_585),
.B1(n_587),
.B2(n_592),
.Y(n_625)
);

BUFx12_ASAP7_75t_L g607 ( 
.A(n_558),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_607),
.B(n_582),
.Y(n_623)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_608),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_609),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_591),
.B(n_569),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_610),
.B(n_611),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_590),
.B(n_571),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_586),
.B(n_574),
.C(n_559),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_614),
.B(n_619),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_617),
.A2(n_625),
.B1(n_597),
.B2(n_607),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_618),
.A2(n_593),
.B(n_606),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_586),
.B(n_570),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_589),
.B(n_573),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_621),
.B(n_623),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_624),
.B(n_626),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_604),
.B(n_583),
.C(n_577),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_628),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_609),
.B(n_601),
.C(n_588),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_629),
.B(n_634),
.Y(n_652)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_630),
.Y(n_649)
);

AOI21x1_ASAP7_75t_L g631 ( 
.A1(n_612),
.A2(n_616),
.B(n_626),
.Y(n_631)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_631),
.Y(n_651)
);

CKINVDCx16_ASAP7_75t_R g634 ( 
.A(n_617),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_614),
.B(n_624),
.C(n_623),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_635),
.B(n_642),
.C(n_178),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_615),
.B(n_367),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_639),
.B(n_640),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_620),
.B(n_367),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_613),
.A2(n_607),
.B(n_331),
.Y(n_641)
);

OAI21xp33_ASAP7_75t_L g654 ( 
.A1(n_641),
.A2(n_346),
.B(n_204),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_622),
.B(n_303),
.C(n_362),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_632),
.A2(n_622),
.B1(n_625),
.B2(n_373),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_645),
.B(n_289),
.Y(n_662)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_629),
.B(n_331),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g659 ( 
.A(n_646),
.B(n_650),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_633),
.B(n_220),
.Y(n_647)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_647),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_648),
.Y(n_657)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_636),
.B(n_635),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_SL g653 ( 
.A1(n_628),
.A2(n_293),
.B1(n_339),
.B2(n_227),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_653),
.A2(n_654),
.B1(n_222),
.B2(n_346),
.Y(n_660)
);

XOR2xp5_ASAP7_75t_L g655 ( 
.A(n_650),
.B(n_637),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_655),
.B(n_660),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_643),
.B(n_632),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_658),
.B(n_661),
.Y(n_667)
);

AOI322xp5_ASAP7_75t_L g661 ( 
.A1(n_651),
.A2(n_627),
.A3(n_638),
.B1(n_641),
.B2(n_630),
.C1(n_642),
.C2(n_294),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_662),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_655),
.B(n_652),
.C(n_649),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_663),
.B(n_666),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_657),
.B(n_647),
.C(n_646),
.Y(n_666)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_667),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_SL g672 ( 
.A1(n_669),
.A2(n_670),
.B(n_644),
.Y(n_672)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_664),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g671 ( 
.A(n_668),
.B(n_665),
.C(n_659),
.Y(n_671)
);

AOI322xp5_ASAP7_75t_L g673 ( 
.A1(n_671),
.A2(n_672),
.A3(n_656),
.B1(n_654),
.B2(n_659),
.C1(n_289),
.C2(n_294),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_673),
.A2(n_239),
.B1(n_224),
.B2(n_169),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_674),
.A2(n_224),
.B(n_169),
.Y(n_675)
);

XOR2xp5_ASAP7_75t_L g676 ( 
.A(n_675),
.B(n_219),
.Y(n_676)
);


endmodule