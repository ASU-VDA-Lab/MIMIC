module real_jpeg_8615_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_244;
wire n_213;
wire n_128;
wire n_179;
wire n_167;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx24_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_40),
.B1(n_56),
.B2(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_1),
.A2(n_26),
.B1(n_29),
.B2(n_40),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_2),
.A2(n_26),
.B1(n_29),
.B2(n_46),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_46),
.B1(n_56),
.B2(n_57),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_4),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_4),
.A2(n_53),
.B(n_57),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_4),
.A2(n_51),
.B1(n_59),
.B2(n_147),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_4),
.B(n_63),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_4),
.A2(n_37),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_4),
.B(n_37),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_4),
.A2(n_79),
.B1(n_80),
.B2(n_223),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_37),
.B(n_42),
.C(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_37),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_7),
.A2(n_26),
.B1(n_29),
.B2(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_SL g68 ( 
.A(n_8),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_10),
.A2(n_26),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_10),
.A2(n_34),
.B1(n_51),
.B2(n_59),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_10),
.A2(n_34),
.B1(n_56),
.B2(n_57),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_10),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_11),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_11),
.A2(n_28),
.B1(n_56),
.B2(n_57),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_11),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_11),
.A2(n_28),
.B1(n_51),
.B2(n_59),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_13),
.A2(n_51),
.B1(n_59),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_13),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_13),
.A2(n_56),
.B1(n_57),
.B2(n_143),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_143),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_13),
.A2(n_26),
.B1(n_29),
.B2(n_143),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_14),
.A2(n_51),
.B1(n_59),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_14),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_99),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_14),
.A2(n_26),
.B1(n_29),
.B2(n_99),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_99),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_15),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_15),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_15),
.A2(n_26),
.B1(n_29),
.B2(n_60),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_15),
.A2(n_37),
.B1(n_38),
.B2(n_60),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_126),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_103),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_19),
.B(n_103),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.C(n_87),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_20),
.A2(n_21),
.B1(n_76),
.B2(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_47),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_22),
.B(n_48),
.C(n_75),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_23),
.B(n_35),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_24),
.A2(n_80),
.B(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_25),
.B(n_31),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_26),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_214)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_29),
.B(n_44),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_29),
.B(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_30),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_30),
.A2(n_31),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_31),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_32),
.A2(n_79),
.B(n_207),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_33),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_36),
.A2(n_43),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_38),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_37),
.B(n_67),
.Y(n_251)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_38),
.A2(n_72),
.B1(n_246),
.B2(n_251),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_45),
.B(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_41),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_41),
.A2(n_43),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_41),
.A2(n_43),
.B1(n_213),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_41),
.A2(n_43),
.B1(n_236),
.B2(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_41),
.A2(n_119),
.B(n_244),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_42),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_43),
.B(n_147),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_64),
.B2(n_75),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_58),
.B(n_61),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_55),
.B1(n_58),
.B2(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_50),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_50),
.A2(n_55),
.B1(n_98),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_50),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_54),
.C(n_55),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_51),
.A2(n_52),
.B(n_147),
.C(n_148),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_66),
.B(n_67),
.C(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_67),
.Y(n_72)
);

HAxp5_ASAP7_75t_SL g246 ( 
.A(n_57),
.B(n_147),
.CON(n_246),
.SN(n_246)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_62),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_63),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B(n_70),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_74),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_65),
.A2(n_137),
.B1(n_138),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_65),
.A2(n_137),
.B1(n_168),
.B2(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_65),
.B(n_147),
.Y(n_234)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_71),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_66),
.B(n_101),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_66),
.A2(n_71),
.B1(n_191),
.B2(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_69),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_71),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_76),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_86),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_78),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_82),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B(n_81),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_79),
.A2(n_80),
.B1(n_90),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_79),
.A2(n_80),
.B1(n_205),
.B2(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_79),
.A2(n_81),
.B(n_91),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_80),
.B(n_147),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_84),
.A2(n_95),
.B(n_121),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_96),
.C(n_100),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_89),
.B(n_92),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_103),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_114),
.CI(n_123),
.CON(n_103),
.SN(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_112),
.B2(n_113),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_112),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_118),
.B(n_122),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_154),
.B(n_277),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_151),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_128),
.B(n_151),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_133),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_132),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_133),
.A2(n_134),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.C(n_144),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B(n_139),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_196),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_177),
.B(n_195),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_197),
.C(n_276),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_174),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_174),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.C(n_173),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_167),
.B1(n_173),
.B2(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_173),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_175),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_178),
.B(n_180),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.C(n_186),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_181),
.B(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_184),
.A2(n_186),
.B1(n_187),
.B2(n_274),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_184),
.Y(n_274)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.C(n_193),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_188),
.A2(n_189),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_192),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_270),
.B(n_275),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_255),
.B(n_269),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_239),
.B(n_254),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_230),
.B(n_238),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_219),
.B(n_229),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_203),
.B(n_208),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_218),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_209),
.B(n_218),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_212),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_214),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_224),
.B(n_228),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_222),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_232),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_233),
.B(n_240),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.CI(n_237),
.CON(n_233),
.SN(n_233)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_249),
.B2(n_253),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_245),
.B1(n_247),
.B2(n_248),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_243),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_245),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_248),
.C(n_253),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_249),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_252),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_257),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_263),
.B2(n_264),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_266),
.C(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_265),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_272),
.Y(n_275)
);


endmodule