module fake_jpeg_17545_n_204 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_0),
.B(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_11),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_35),
.B(n_39),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_36),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_15),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_25),
.Y(n_61)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_51),
.B1(n_58),
.B2(n_27),
.Y(n_87)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_28),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_22),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_28),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_17),
.A2(n_9),
.B1(n_24),
.B2(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_33),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_33),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_17),
.A2(n_24),
.B1(n_32),
.B2(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_61),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_62),
.B(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_29),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_70),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_23),
.Y(n_71)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_83),
.Y(n_96)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_23),
.Y(n_78)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_26),
.CI(n_49),
.CON(n_93),
.SN(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_19),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_81),
.B(n_82),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_36),
.B(n_26),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_42),
.B1(n_46),
.B2(n_54),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_89),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_40),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_43),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_99),
.Y(n_120)
);

HAxp5_ASAP7_75t_SL g131 ( 
.A(n_93),
.B(n_85),
.CON(n_131),
.SN(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_114),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_85),
.B1(n_106),
.B2(n_117),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_54),
.A3(n_75),
.B1(n_66),
.B2(n_82),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_103),
.A2(n_105),
.B1(n_115),
.B2(n_116),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_78),
.B1(n_73),
.B2(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_68),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_85),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_63),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_73),
.B(n_63),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_109),
.C(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_67),
.B1(n_65),
.B2(n_89),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_65),
.B1(n_90),
.B2(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_77),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_124),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_77),
.CI(n_76),
.CON(n_124),
.SN(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_74),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_131),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_102),
.B1(n_107),
.B2(n_119),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_141),
.C(n_124),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_85),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_142),
.B(n_120),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_118),
.C(n_114),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_93),
.A2(n_103),
.B(n_116),
.C(n_115),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_113),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_97),
.C(n_119),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_100),
.B1(n_108),
.B2(n_111),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_149),
.B1(n_155),
.B2(n_153),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_151),
.C(n_162),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_95),
.B1(n_104),
.B2(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_142),
.B1(n_132),
.B2(n_133),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_95),
.C(n_139),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_155),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_124),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_SL g168 ( 
.A(n_154),
.B(n_133),
.C(n_125),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_152),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_161),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_121),
.B1(n_126),
.B2(n_129),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_134),
.B1(n_132),
.B2(n_130),
.Y(n_165)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_134),
.C(n_127),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_170),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_160),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_175),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_127),
.C(n_162),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_174),
.C(n_158),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_159),
.C(n_148),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_145),
.B(n_153),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_177),
.A2(n_172),
.B(n_157),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_185),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_161),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_150),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_184),
.A2(n_180),
.B1(n_168),
.B2(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_192),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_164),
.B(n_144),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_190),
.B(n_182),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_175),
.B1(n_154),
.B2(n_164),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_169),
.B(n_173),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_186),
.B(n_181),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_195),
.C(n_188),
.Y(n_201)
);

NAND4xp25_ASAP7_75t_SL g196 ( 
.A(n_192),
.B(n_179),
.C(n_183),
.D(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_190),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

OAI21x1_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_196),
.B(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_189),
.B(n_198),
.C(n_200),
.Y(n_203)
);


endmodule