module fake_jpeg_16893_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_56),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_60),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_0),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_17),
.B(n_32),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_21),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_36),
.B1(n_29),
.B2(n_31),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_72),
.B1(n_41),
.B2(n_27),
.Y(n_92)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_30),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_36),
.B1(n_29),
.B2(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_74),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_85),
.Y(n_128)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_82),
.B(n_106),
.Y(n_118)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_95),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_36),
.B1(n_24),
.B2(n_16),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_104),
.B1(n_109),
.B2(n_64),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_93),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_24),
.B1(n_46),
.B2(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_97),
.B1(n_99),
.B2(n_105),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_41),
.B(n_16),
.C(n_27),
.Y(n_89)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_100),
.B1(n_103),
.B2(n_63),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_17),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_48),
.B1(n_47),
.B2(n_44),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_26),
.B1(n_47),
.B2(n_44),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_26),
.B1(n_35),
.B2(n_34),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_59),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_48),
.B(n_44),
.C(n_43),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_59),
.B(n_32),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_71),
.Y(n_129)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_50),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_32),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_32),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_114),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_71),
.B1(n_53),
.B2(n_50),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_135),
.B1(n_110),
.B2(n_85),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_105),
.B1(n_102),
.B2(n_43),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_96),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_91),
.Y(n_172)
);

CKINVDCx6p67_ASAP7_75t_R g130 ( 
.A(n_75),
.Y(n_130)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_98),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_133),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_98),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_0),
.B(n_1),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_53),
.B1(n_39),
.B2(n_48),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_77),
.B(n_62),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_77),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_93),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_147),
.B1(n_158),
.B2(n_127),
.Y(n_182)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_84),
.B1(n_79),
.B2(n_81),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_76),
.B1(n_105),
.B2(n_80),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_174),
.B1(n_114),
.B2(n_121),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_82),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_79),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_168),
.Y(n_189)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_166),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_117),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_155),
.B(n_161),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_81),
.C(n_111),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_160),
.C(n_163),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_112),
.B(n_89),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_157),
.B(n_165),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_108),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_118),
.B(n_97),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_117),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_40),
.C(n_91),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_113),
.B(n_20),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_101),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_122),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_173),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_172),
.B(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_125),
.A2(n_94),
.B1(n_83),
.B2(n_62),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_183),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_161),
.B1(n_155),
.B2(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_172),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_124),
.A3(n_113),
.B1(n_135),
.B2(n_128),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_151),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_190),
.A2(n_191),
.B1(n_199),
.B2(n_204),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_119),
.B1(n_118),
.B2(n_141),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_192),
.B(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_148),
.A2(n_132),
.B(n_133),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_194),
.A2(n_203),
.B(n_130),
.Y(n_231)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_202),
.B(n_173),
.Y(n_210)
);

NOR2x1_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_128),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_148),
.A2(n_119),
.B1(n_138),
.B2(n_137),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_153),
.B(n_152),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_139),
.B(n_138),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_142),
.A2(n_127),
.B1(n_115),
.B2(n_139),
.Y(n_204)
);

XNOR2x1_ASAP7_75t_SL g205 ( 
.A(n_144),
.B(n_160),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_169),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_147),
.A2(n_127),
.B1(n_39),
.B2(n_43),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_206),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_231),
.B(n_175),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_156),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_212),
.C(n_217),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_163),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_213),
.B(n_221),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_154),
.B(n_168),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_214),
.A2(n_198),
.B(n_177),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_220),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_165),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_235),
.B1(n_237),
.B2(n_195),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_224),
.B(n_230),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_162),
.B(n_130),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_225),
.B(n_203),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_162),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_199),
.A2(n_130),
.B1(n_62),
.B2(n_70),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_228),
.A2(n_190),
.B1(n_208),
.B2(n_201),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_185),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_188),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_234),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_184),
.A2(n_39),
.B1(n_70),
.B2(n_2),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_202),
.B(n_33),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_196),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_247),
.B(n_251),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_239),
.A2(n_228),
.B1(n_226),
.B2(n_13),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_178),
.Y(n_240)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_222),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_212),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_250),
.C(n_258),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_179),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_187),
.C(n_198),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_187),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_210),
.B(n_175),
.C(n_191),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_181),
.B1(n_177),
.B2(n_207),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_237),
.B1(n_234),
.B2(n_209),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_193),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_223),
.Y(n_276)
);

A2O1A1O1Ixp25_ASAP7_75t_L g261 ( 
.A1(n_213),
.A2(n_188),
.B(n_40),
.C(n_176),
.D(n_18),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_261),
.B(n_214),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_40),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_231),
.Y(n_268)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_255),
.B(n_232),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_265),
.B(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_219),
.Y(n_266)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_275),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_241),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_279),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_273),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_229),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_280),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_245),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_253),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_242),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_257),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_238),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_33),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_243),
.C(n_244),
.Y(n_287)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_289),
.C(n_291),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_243),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_290),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_250),
.C(n_252),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_268),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_254),
.C(n_262),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_254),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_251),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_260),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_276),
.B1(n_264),
.B2(n_279),
.Y(n_301)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_301),
.Y(n_320)
);

OAI21x1_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_269),
.B(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_302),
.Y(n_326)
);

OAI321xp33_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_282),
.A3(n_273),
.B1(n_281),
.B2(n_263),
.C(n_276),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_306),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_274),
.C(n_270),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_3),
.Y(n_324)
);

XNOR2x1_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_272),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_3),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_308),
.Y(n_321)
);

AOI221xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_12),
.B1(n_14),
.B2(n_13),
.C(n_11),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_34),
.B1(n_35),
.B2(n_10),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_9),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_290),
.B(n_12),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_285),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_9),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_8),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_317),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_18),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_305),
.A2(n_285),
.B1(n_288),
.B2(n_35),
.Y(n_322)
);

OA21x2_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_324),
.B(n_33),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_307),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g334 ( 
.A1(n_323),
.A2(n_325),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_19),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_326),
.A3(n_306),
.B1(n_319),
.B2(n_322),
.C1(n_313),
.C2(n_314),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_329),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_311),
.B(n_308),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_328),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_321),
.A2(n_303),
.B(n_8),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_34),
.C(n_18),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_331),
.Y(n_339)
);

AOI31xp67_ASAP7_75t_L g336 ( 
.A1(n_332),
.A2(n_334),
.A3(n_3),
.B(n_4),
.Y(n_336)
);

A2O1A1O1Ixp25_ASAP7_75t_L g335 ( 
.A1(n_327),
.A2(n_19),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_335)
);

OAI21x1_ASAP7_75t_SL g341 ( 
.A1(n_335),
.A2(n_336),
.B(n_332),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_333),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_340),
.B(n_341),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_342),
.B(n_337),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_339),
.B(n_5),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_6),
.Y(n_345)
);


endmodule