module fake_jpeg_7822_n_279 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_18),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_19),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_29),
.B1(n_22),
.B2(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_58),
.B1(n_62),
.B2(n_64),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_21),
.B1(n_33),
.B2(n_29),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_50),
.B(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_51),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_21),
.B1(n_33),
.B2(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_22),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_33),
.B1(n_26),
.B2(n_24),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_23),
.C(n_34),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_57),
.C(n_23),
.Y(n_89)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_24),
.B1(n_26),
.B2(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_40),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_24),
.B1(n_26),
.B2(n_17),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_27),
.B1(n_20),
.B2(n_28),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_68),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_82),
.B1(n_66),
.B2(n_56),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_44),
.B1(n_32),
.B2(n_31),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_50),
.B1(n_58),
.B2(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_14),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_86),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_32),
.B1(n_43),
.B2(n_41),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_55),
.B1(n_86),
.B2(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_55),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_1),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_54),
.B(n_52),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_57),
.B(n_53),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_19),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_57),
.Y(n_111)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_46),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_114),
.B(n_90),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_77),
.B1(n_69),
.B2(n_88),
.Y(n_133)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_107),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_117),
.B1(n_89),
.B2(n_84),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_45),
.B1(n_47),
.B2(n_63),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_102),
.B1(n_86),
.B2(n_82),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_47),
.B1(n_66),
.B2(n_63),
.Y(n_102)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_113),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_82),
.B1(n_92),
.B2(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_104),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_66),
.B1(n_61),
.B2(n_56),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_57),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_39),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_88),
.B(n_111),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_119),
.B(n_128),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_75),
.B(n_73),
.C(n_81),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_122),
.B(n_123),
.Y(n_169)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_130),
.B1(n_133),
.B2(n_139),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_138),
.B1(n_106),
.B2(n_95),
.Y(n_159)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_94),
.B(n_118),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_73),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_134),
.B(n_141),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_69),
.B(n_93),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_137),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_104),
.B(n_77),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_100),
.A2(n_61),
.B1(n_53),
.B2(n_67),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_78),
.B1(n_67),
.B2(n_85),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_1),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_19),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_146),
.B(n_148),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_144),
.B1(n_130),
.B2(n_137),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_159),
.B1(n_103),
.B2(n_32),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_153),
.B(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_161),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_97),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_171),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_116),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_167),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_95),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_123),
.A2(n_107),
.B1(n_99),
.B2(n_109),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_92),
.B1(n_103),
.B2(n_141),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_99),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_174),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_127),
.B1(n_131),
.B2(n_120),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_180),
.B1(n_184),
.B2(n_169),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_163),
.B1(n_147),
.B2(n_159),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_131),
.B(n_120),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_188),
.B(n_190),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_142),
.B1(n_119),
.B2(n_103),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_141),
.B1(n_92),
.B2(n_31),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

NAND2x1_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_35),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_32),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_155),
.Y(n_212)
);

NAND2xp33_ASAP7_75t_R g196 ( 
.A(n_150),
.B(n_35),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_164),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_151),
.A2(n_79),
.B(n_2),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_188),
.B1(n_179),
.B2(n_191),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_172),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_206),
.A2(n_208),
.B1(n_209),
.B2(n_212),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_156),
.C(n_184),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_215),
.C(n_203),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_178),
.A2(n_171),
.B1(n_148),
.B2(n_164),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_155),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_217),
.B(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_183),
.B(n_168),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_SL g224 ( 
.A(n_213),
.B(n_181),
.C(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_218),
.B1(n_175),
.B2(n_195),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_43),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_40),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_178),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_225),
.C(n_231),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_224),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_226),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_208),
.C(n_211),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_218),
.B1(n_199),
.B2(n_214),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_229),
.B1(n_198),
.B2(n_201),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_180),
.B1(n_190),
.B2(n_175),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_193),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_176),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_233),
.A2(n_201),
.B1(n_194),
.B2(n_174),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_194),
.A3(n_195),
.B1(n_174),
.B2(n_79),
.C1(n_7),
.C2(n_8),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_234),
.Y(n_240)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_3),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_232),
.B(n_202),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_245),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_248),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_221),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_223),
.C(n_224),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_43),
.C(n_41),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_246),
.C(n_233),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_40),
.C(n_39),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_3),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_4),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_222),
.B(n_4),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_249),
.B(n_256),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_242),
.B(n_40),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_244),
.B(n_242),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_230),
.B(n_227),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_7),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_227),
.B1(n_231),
.B2(n_6),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_6),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_240),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_4),
.B(n_5),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_5),
.B(n_6),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_5),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_264),
.Y(n_271)
);

AOI221xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_266),
.B1(n_10),
.B2(n_12),
.C(n_13),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_262),
.C(n_251),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_265),
.A2(n_253),
.B1(n_252),
.B2(n_13),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_267),
.B(n_268),
.Y(n_273)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_272),
.B(n_14),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_10),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_10),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_23),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_40),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_SL g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_269),
.B(n_271),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_273),
.Y(n_279)
);


endmodule