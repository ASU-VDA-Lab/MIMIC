module fake_netlist_6_1497_n_1434 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_366, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_190, n_262, n_187, n_60, n_361, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1434);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1434;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1382;
wire n_1372;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_1058;
wire n_854;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1109;
wire n_712;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_230),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_345),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_327),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_157),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_84),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_206),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_262),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_61),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_329),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_273),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_186),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_159),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_269),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_228),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_176),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_291),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_42),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_107),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_271),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_235),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_339),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_177),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_80),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_19),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_317),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_201),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_54),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_192),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_95),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_300),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_132),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_250),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_123),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_133),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_264),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_355),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_263),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_180),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_120),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_199),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_87),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_69),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_292),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_119),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_137),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_315),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_5),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_267),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_234),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_312),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_163),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_334),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_13),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_172),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_90),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_216),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_337),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_15),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_217),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_226),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_268),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_111),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_227),
.Y(n_432)
);

BUFx5_ASAP7_75t_L g433 ( 
.A(n_249),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_306),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_81),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_277),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_62),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_168),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_324),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_85),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_242),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_165),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_79),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_310),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_58),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_166),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_354),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_320),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_42),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_104),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_222),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_332),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_49),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_299),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_319),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_330),
.Y(n_456)
);

BUFx10_ASAP7_75t_L g457 ( 
.A(n_215),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_202),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_94),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_130),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_154),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_366),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_239),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_117),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_60),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_335),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_73),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_179),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_279),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_39),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_16),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_96),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_203),
.Y(n_473)
);

BUFx10_ASAP7_75t_L g474 ( 
.A(n_240),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_71),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_48),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_40),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_289),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_350),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_200),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_358),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_189),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_167),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_77),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_255),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_261),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_102),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_333),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_284),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_353),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_25),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_15),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_285),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_128),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_151),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_3),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_357),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_283),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_82),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_149),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_45),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_122),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_270),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_185),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_363),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_280),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_288),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_13),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_218),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_309),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_296),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g512 ( 
.A(n_257),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_139),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_361),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_131),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_118),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_147),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_65),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_34),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_205),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_260),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_31),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_57),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_91),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_77),
.Y(n_525)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_71),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_301),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_27),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_304),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_97),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_243),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_188),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_341),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_244),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_311),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_246),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_316),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_55),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_136),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_148),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_9),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_181),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g543 ( 
.A(n_21),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_340),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_142),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_360),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_433),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_461),
.B(n_0),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_508),
.B(n_0),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_406),
.B(n_1),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_370),
.B(n_1),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_433),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_404),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_367),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_406),
.B(n_2),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_508),
.B(n_2),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_512),
.B(n_3),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_404),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_404),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_392),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_512),
.B(n_4),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_400),
.B(n_417),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_400),
.B(n_4),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_417),
.B(n_5),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_404),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_373),
.B(n_6),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_420),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_416),
.B(n_6),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_392),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_384),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_410),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_422),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_433),
.Y(n_573)
);

BUFx12f_ASAP7_75t_L g574 ( 
.A(n_408),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_445),
.B(n_543),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_418),
.B(n_7),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_465),
.Y(n_577)
);

BUFx12f_ASAP7_75t_L g578 ( 
.A(n_408),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_389),
.B(n_462),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_456),
.B(n_7),
.Y(n_580)
);

BUFx12f_ASAP7_75t_L g581 ( 
.A(n_408),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_418),
.B(n_8),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_419),
.B(n_8),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_429),
.B(n_9),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_369),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_433),
.Y(n_586)
);

BUFx12f_ASAP7_75t_L g587 ( 
.A(n_444),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_419),
.B(n_10),
.Y(n_588)
);

BUFx12f_ASAP7_75t_L g589 ( 
.A(n_444),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_490),
.B(n_10),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_484),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_389),
.B(n_11),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_433),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_433),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_462),
.B(n_472),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_518),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_472),
.B(n_11),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_487),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_487),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_420),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_420),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_420),
.B(n_83),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_490),
.B(n_12),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_475),
.B(n_12),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_368),
.B(n_14),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_371),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_383),
.B(n_14),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_432),
.B(n_16),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_499),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_499),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_464),
.B(n_17),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_395),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_433),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_415),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_507),
.B(n_17),
.Y(n_616)
);

CKINVDCx16_ASAP7_75t_R g617 ( 
.A(n_442),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_499),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_444),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_457),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_505),
.B(n_18),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_521),
.B(n_86),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_375),
.B(n_18),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_427),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_376),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_521),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_521),
.Y(n_627)
);

AND2x6_ASAP7_75t_L g628 ( 
.A(n_521),
.B(n_88),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_437),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_516),
.B(n_19),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_377),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_379),
.B(n_20),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_385),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_546),
.B(n_20),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_386),
.B(n_21),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_388),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_402),
.B(n_22),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_457),
.B(n_22),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_414),
.B(n_23),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_426),
.B(n_23),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_457),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_430),
.B(n_440),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_526),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_443),
.B(n_24),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_474),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_554),
.B(n_447),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_585),
.B(n_460),
.Y(n_647)
);

OAI22xp33_ASAP7_75t_L g648 ( 
.A1(n_623),
.A2(n_612),
.B1(n_619),
.B2(n_591),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_608),
.A2(n_494),
.B1(n_393),
.B2(n_436),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_612),
.A2(n_453),
.B1(n_467),
.B2(n_449),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_558),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_579),
.B(n_474),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_607),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_558),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_613),
.B(n_470),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_558),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_621),
.A2(n_494),
.B1(n_441),
.B2(n_387),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_595),
.B(n_474),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_615),
.B(n_372),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_641),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_559),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_559),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_559),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_624),
.B(n_374),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_SL g665 ( 
.A1(n_548),
.A2(n_491),
.B1(n_501),
.B2(n_471),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_629),
.B(n_575),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_601),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_601),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_598),
.B(n_378),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_SL g670 ( 
.A1(n_551),
.A2(n_542),
.B1(n_510),
.B2(n_477),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_599),
.B(n_380),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_630),
.A2(n_492),
.B1(n_496),
.B2(n_476),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_601),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_641),
.B(n_381),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_641),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_604),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_550),
.A2(n_522),
.B1(n_523),
.B2(n_519),
.Y(n_677)
);

AO22x2_ASAP7_75t_L g678 ( 
.A1(n_592),
.A2(n_597),
.B1(n_638),
.B2(n_555),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_645),
.B(n_525),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_557),
.A2(n_538),
.B1(n_541),
.B2(n_528),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_R g681 ( 
.A1(n_566),
.A2(n_483),
.B1(n_489),
.B2(n_478),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_645),
.B(n_382),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_561),
.A2(n_617),
.B1(n_568),
.B2(n_616),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_604),
.Y(n_684)
);

AO22x2_ASAP7_75t_L g685 ( 
.A1(n_592),
.A2(n_500),
.B1(n_502),
.B2(n_493),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_560),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_625),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_620),
.B(n_503),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_604),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_631),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_609),
.A2(n_391),
.B1(n_394),
.B2(n_390),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_549),
.A2(n_514),
.B1(n_515),
.B2(n_504),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_634),
.A2(n_397),
.B1(n_398),
.B2(n_396),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_618),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_618),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_618),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_626),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_626),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_626),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_627),
.Y(n_700)
);

AO22x2_ASAP7_75t_L g701 ( 
.A1(n_597),
.A2(n_532),
.B1(n_535),
.B2(n_530),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_645),
.B(n_537),
.Y(n_702)
);

OAI22xp33_ASAP7_75t_SL g703 ( 
.A1(n_643),
.A2(n_401),
.B1(n_403),
.B2(n_399),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_580),
.A2(n_407),
.B1(n_409),
.B2(n_405),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_574),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_578),
.B(n_24),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_613),
.B(n_25),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_643),
.A2(n_412),
.B1(n_413),
.B2(n_411),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_L g709 ( 
.A1(n_549),
.A2(n_423),
.B1(n_424),
.B2(n_421),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_581),
.A2(n_428),
.B1(n_431),
.B2(n_425),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_627),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_L g712 ( 
.A1(n_556),
.A2(n_435),
.B1(n_438),
.B2(n_434),
.Y(n_712)
);

OAI22xp33_ASAP7_75t_L g713 ( 
.A1(n_556),
.A2(n_446),
.B1(n_448),
.B2(n_439),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_587),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_589),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_L g716 ( 
.A1(n_605),
.A2(n_451),
.B1(n_452),
.B2(n_450),
.Y(n_716)
);

AO22x2_ASAP7_75t_L g717 ( 
.A1(n_606),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_717)
);

AO22x2_ASAP7_75t_L g718 ( 
.A1(n_606),
.A2(n_29),
.B1(n_26),
.B2(n_28),
.Y(n_718)
);

OAI22xp33_ASAP7_75t_L g719 ( 
.A1(n_605),
.A2(n_455),
.B1(n_458),
.B2(n_454),
.Y(n_719)
);

AO22x2_ASAP7_75t_L g720 ( 
.A1(n_635),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_584),
.A2(n_463),
.B1(n_466),
.B2(n_459),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_588),
.A2(n_469),
.B1(n_473),
.B2(n_468),
.Y(n_722)
);

OAI22xp33_ASAP7_75t_L g723 ( 
.A1(n_632),
.A2(n_639),
.B1(n_640),
.B2(n_637),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_SL g724 ( 
.A1(n_632),
.A2(n_480),
.B1(n_481),
.B2(n_479),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_627),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_SL g726 ( 
.A1(n_645),
.A2(n_485),
.B1(n_486),
.B2(n_482),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_635),
.A2(n_495),
.B1(n_497),
.B2(n_488),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_633),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_569),
.Y(n_729)
);

INVxp33_ASAP7_75t_L g730 ( 
.A(n_666),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_649),
.Y(n_731)
);

XOR2x2_ASAP7_75t_L g732 ( 
.A(n_665),
.B(n_637),
.Y(n_732)
);

AND2x4_ASAP7_75t_SL g733 ( 
.A(n_652),
.B(n_644),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_653),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_687),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_L g736 ( 
.A1(n_723),
.A2(n_642),
.B(n_562),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_690),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_651),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_651),
.Y(n_739)
);

XOR2xp5_ASAP7_75t_L g740 ( 
.A(n_657),
.B(n_498),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_661),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_661),
.Y(n_742)
);

XNOR2x2_ASAP7_75t_L g743 ( 
.A(n_717),
.B(n_563),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_688),
.B(n_644),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_662),
.Y(n_745)
);

XNOR2xp5_ASAP7_75t_L g746 ( 
.A(n_670),
.B(n_639),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_662),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_668),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_668),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_676),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_676),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_675),
.Y(n_752)
);

XOR2xp5_ASAP7_75t_L g753 ( 
.A(n_705),
.B(n_506),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_689),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_689),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_654),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_698),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_658),
.B(n_636),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_698),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_663),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_663),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_684),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_684),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_688),
.B(n_570),
.Y(n_764)
);

XOR2xp5_ASAP7_75t_L g765 ( 
.A(n_715),
.B(n_509),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_669),
.B(n_671),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_696),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_696),
.Y(n_768)
);

XNOR2x2_ASAP7_75t_L g769 ( 
.A(n_717),
.B(n_563),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_686),
.Y(n_770)
);

CKINVDCx16_ASAP7_75t_R g771 ( 
.A(n_710),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_656),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_667),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_673),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_694),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_646),
.B(n_562),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_695),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_697),
.B(n_571),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_659),
.B(n_572),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_699),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_724),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_682),
.B(n_600),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_729),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_700),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_711),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_647),
.B(n_633),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_725),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_725),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_725),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_707),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_664),
.B(n_577),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_660),
.B(n_596),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_728),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_728),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_728),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_678),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_678),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_702),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_685),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_685),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_701),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_701),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_674),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_655),
.B(n_633),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_718),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_718),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_720),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_683),
.B(n_553),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_720),
.Y(n_809)
);

INVxp33_ASAP7_75t_SL g810 ( 
.A(n_691),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_709),
.B(n_564),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_672),
.B(n_693),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_722),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_714),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_679),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_721),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_677),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_727),
.B(n_547),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_680),
.B(n_553),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_704),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_776),
.B(n_712),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_770),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_796),
.B(n_706),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_815),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_776),
.B(n_713),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_758),
.B(n_640),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_786),
.B(n_716),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_783),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_815),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_756),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_783),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_786),
.B(n_719),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_779),
.B(n_564),
.Y(n_833)
);

AND2x2_ASAP7_75t_SL g834 ( 
.A(n_812),
.B(n_576),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_736),
.A2(n_648),
.B(n_692),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_791),
.B(n_576),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_804),
.B(n_582),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_756),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_815),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_811),
.A2(n_708),
.B(n_703),
.Y(n_840)
);

BUFx12f_ASAP7_75t_L g841 ( 
.A(n_814),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_738),
.Y(n_842)
);

NAND2x1p5_ASAP7_75t_L g843 ( 
.A(n_797),
.B(n_815),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_790),
.Y(n_844)
);

INVxp67_ASAP7_75t_SL g845 ( 
.A(n_803),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_733),
.B(n_803),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_798),
.B(n_726),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_730),
.B(n_650),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_733),
.B(n_582),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_SL g850 ( 
.A(n_811),
.B(n_583),
.Y(n_850)
);

AND2x2_ASAP7_75t_SL g851 ( 
.A(n_771),
.B(n_583),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_808),
.B(n_590),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_790),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_778),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_778),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_766),
.B(n_590),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_744),
.B(n_603),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_734),
.B(n_706),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_735),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_752),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_818),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_737),
.Y(n_862)
);

AND2x4_ASAP7_75t_SL g863 ( 
.A(n_818),
.B(n_552),
.Y(n_863)
);

NOR2xp67_ASAP7_75t_L g864 ( 
.A(n_820),
.B(n_511),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_816),
.B(n_513),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_813),
.A2(n_818),
.B(n_819),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_778),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_744),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_744),
.B(n_603),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_799),
.B(n_573),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_739),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_741),
.Y(n_872)
);

BUFx5_ASAP7_75t_L g873 ( 
.A(n_742),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_792),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_745),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_764),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_747),
.B(n_602),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_730),
.B(n_586),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_814),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_800),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_748),
.B(n_602),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_764),
.B(n_593),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_764),
.B(n_594),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_801),
.B(n_602),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_749),
.B(n_602),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_802),
.B(n_614),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_805),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_753),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_750),
.B(n_622),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_806),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_751),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_754),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_772),
.B(n_622),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_765),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_807),
.B(n_517),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_755),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_757),
.B(n_622),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_759),
.B(n_622),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_740),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_773),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_809),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_781),
.B(n_520),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_774),
.B(n_524),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_775),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_777),
.B(n_527),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_732),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_746),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_782),
.B(n_628),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_793),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_794),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_780),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_784),
.Y(n_912)
);

AND2x2_ASAP7_75t_SL g913 ( 
.A(n_769),
.B(n_681),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_785),
.B(n_628),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_810),
.B(n_529),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_760),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_876),
.B(n_761),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_828),
.Y(n_918)
);

NOR2x1_ASAP7_75t_L g919 ( 
.A(n_866),
.B(n_781),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_831),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_852),
.B(n_732),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_902),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_852),
.B(n_731),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_841),
.B(n_769),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_830),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_860),
.B(n_743),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_868),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_837),
.B(n_810),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_833),
.B(n_731),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_837),
.B(n_795),
.Y(n_930)
);

INVx4_ASAP7_75t_L g931 ( 
.A(n_868),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_879),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_841),
.B(n_762),
.Y(n_933)
);

OR2x6_ASAP7_75t_L g934 ( 
.A(n_868),
.B(n_763),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_844),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_868),
.Y(n_936)
);

NAND2x1p5_ASAP7_75t_L g937 ( 
.A(n_824),
.B(n_787),
.Y(n_937)
);

BUFx4f_ASAP7_75t_L g938 ( 
.A(n_868),
.Y(n_938)
);

INVx5_ASAP7_75t_L g939 ( 
.A(n_823),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_853),
.Y(n_940)
);

NAND2x1p5_ASAP7_75t_L g941 ( 
.A(n_824),
.B(n_829),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_856),
.B(n_767),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_856),
.B(n_768),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_909),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_833),
.B(n_836),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_879),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_838),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_861),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_880),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_845),
.B(n_788),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_888),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_829),
.Y(n_952)
);

NOR2x1_ASAP7_75t_L g953 ( 
.A(n_821),
.B(n_789),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_836),
.B(n_628),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_838),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_876),
.B(n_817),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_825),
.B(n_531),
.Y(n_957)
);

AND2x6_ASAP7_75t_L g958 ( 
.A(n_884),
.B(n_628),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_839),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_826),
.B(n_533),
.Y(n_960)
);

NOR2x1_ASAP7_75t_L g961 ( 
.A(n_827),
.B(n_817),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_830),
.Y(n_962)
);

BUFx4f_ASAP7_75t_L g963 ( 
.A(n_843),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_842),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_826),
.B(n_834),
.Y(n_965)
);

INVx5_ASAP7_75t_L g966 ( 
.A(n_823),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_878),
.B(n_534),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_839),
.B(n_822),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_872),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_857),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_842),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_822),
.B(n_846),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_878),
.B(n_536),
.Y(n_973)
);

OR2x6_ASAP7_75t_L g974 ( 
.A(n_843),
.B(n_30),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_857),
.B(n_539),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_909),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_869),
.B(n_540),
.Y(n_977)
);

NAND2x1_ASAP7_75t_SL g978 ( 
.A(n_915),
.B(n_32),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_869),
.B(n_544),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_899),
.B(n_848),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_872),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_846),
.B(n_89),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_887),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_909),
.Y(n_984)
);

INVx6_ASAP7_75t_L g985 ( 
.A(n_858),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_859),
.B(n_92),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_969),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_938),
.B(n_931),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_928),
.B(n_834),
.Y(n_989)
);

CKINVDCx8_ASAP7_75t_R g990 ( 
.A(n_946),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_981),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_920),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_956),
.Y(n_993)
);

BUFx12f_ASAP7_75t_L g994 ( 
.A(n_933),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_938),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_925),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_952),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_931),
.B(n_882),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_947),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_918),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_955),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_932),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_948),
.Y(n_1003)
);

INVxp67_ASAP7_75t_SL g1004 ( 
.A(n_941),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_952),
.Y(n_1005)
);

BUFx12f_ASAP7_75t_L g1006 ( 
.A(n_933),
.Y(n_1006)
);

BUFx8_ASAP7_75t_SL g1007 ( 
.A(n_922),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_952),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_963),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_964),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_971),
.Y(n_1011)
);

BUFx2_ASAP7_75t_SL g1012 ( 
.A(n_935),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_962),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_945),
.B(n_851),
.Y(n_1014)
);

INVx5_ASAP7_75t_L g1015 ( 
.A(n_958),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_968),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_951),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_942),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_972),
.B(n_859),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_968),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_984),
.Y(n_1021)
);

INVx6_ASAP7_75t_SL g1022 ( 
.A(n_974),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_956),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_985),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_970),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_929),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_923),
.B(n_921),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_927),
.Y(n_1028)
);

INVx5_ASAP7_75t_L g1029 ( 
.A(n_958),
.Y(n_1029)
);

INVx5_ASAP7_75t_L g1030 ( 
.A(n_958),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_963),
.B(n_882),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_930),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_980),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_928),
.A2(n_850),
.B1(n_835),
.B2(n_851),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_940),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_944),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_933),
.Y(n_1037)
);

CKINVDCx11_ASAP7_75t_R g1038 ( 
.A(n_924),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_972),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_974),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_970),
.B(n_849),
.Y(n_1041)
);

BUFx12f_ASAP7_75t_L g1042 ( 
.A(n_985),
.Y(n_1042)
);

BUFx24_ASAP7_75t_L g1043 ( 
.A(n_982),
.Y(n_1043)
);

INVx6_ASAP7_75t_L g1044 ( 
.A(n_995),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_996),
.Y(n_1045)
);

CKINVDCx6p67_ASAP7_75t_R g1046 ( 
.A(n_1017),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_992),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1034),
.A2(n_989),
.B1(n_965),
.B2(n_919),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1032),
.A2(n_850),
.B(n_954),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_996),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_989),
.A2(n_965),
.B1(n_919),
.B2(n_961),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_992),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_SL g1053 ( 
.A1(n_1014),
.A2(n_913),
.B1(n_906),
.B2(n_924),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1041),
.B(n_1018),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1027),
.A2(n_913),
.B1(n_961),
.B2(n_1026),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_1009),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_1003),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_999),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1025),
.B(n_960),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_1015),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_1042),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1001),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_987),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_993),
.A2(n_1023),
.B1(n_1019),
.B2(n_924),
.Y(n_1064)
);

OAI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_1033),
.A2(n_926),
.B1(n_907),
.B2(n_974),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_991),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1025),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_995),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1013),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1010),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1016),
.A2(n_1020),
.B1(n_1019),
.B2(n_1031),
.Y(n_1071)
);

INVxp33_ASAP7_75t_L g1072 ( 
.A(n_1035),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1036),
.Y(n_1073)
);

CKINVDCx6p67_ASAP7_75t_R g1074 ( 
.A(n_1017),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_1019),
.A2(n_840),
.B1(n_982),
.B2(n_832),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1031),
.A2(n_957),
.B1(n_977),
.B2(n_843),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_SL g1077 ( 
.A1(n_1040),
.A2(n_894),
.B1(n_986),
.B2(n_979),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1039),
.B(n_975),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1022),
.A2(n_986),
.B1(n_849),
.B2(n_874),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_SL g1080 ( 
.A1(n_1037),
.A2(n_966),
.B1(n_939),
.B2(n_858),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_SL g1081 ( 
.A1(n_1012),
.A2(n_858),
.B1(n_983),
.B2(n_847),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1036),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_1007),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_1015),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_1015),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1022),
.A2(n_874),
.B1(n_949),
.B2(n_953),
.Y(n_1086)
);

CKINVDCx11_ASAP7_75t_R g1087 ( 
.A(n_990),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1011),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_SL g1089 ( 
.A1(n_1037),
.A2(n_939),
.B1(n_966),
.B2(n_959),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1022),
.A2(n_953),
.B1(n_863),
.B2(n_895),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1021),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1021),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1000),
.A2(n_864),
.B1(n_865),
.B2(n_967),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1039),
.A2(n_863),
.B1(n_895),
.B2(n_917),
.Y(n_1094)
);

OAI22x1_ASAP7_75t_L g1095 ( 
.A1(n_1043),
.A2(n_995),
.B1(n_966),
.B2(n_939),
.Y(n_1095)
);

INVxp67_ASAP7_75t_SL g1096 ( 
.A(n_1021),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1039),
.A2(n_917),
.B1(n_855),
.B2(n_867),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1043),
.B(n_886),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1051),
.A2(n_1002),
.B1(n_1038),
.B2(n_973),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_SL g1100 ( 
.A(n_1083),
.B(n_1007),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_SL g1101 ( 
.A1(n_1081),
.A2(n_994),
.B1(n_1006),
.B2(n_1002),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1058),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1068),
.Y(n_1103)
);

CKINVDCx14_ASAP7_75t_R g1104 ( 
.A(n_1083),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1068),
.B(n_1039),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_SL g1106 ( 
.A1(n_1048),
.A2(n_994),
.B1(n_1006),
.B2(n_1038),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1058),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1062),
.Y(n_1108)
);

NAND2xp33_ASAP7_75t_SL g1109 ( 
.A(n_1095),
.B(n_1009),
.Y(n_1109)
);

CKINVDCx6p67_ASAP7_75t_R g1110 ( 
.A(n_1087),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1053),
.A2(n_862),
.B1(n_943),
.B2(n_892),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1075),
.A2(n_990),
.B1(n_1003),
.B2(n_1009),
.Y(n_1112)
);

OAI21xp33_ASAP7_75t_SL g1113 ( 
.A1(n_1079),
.A2(n_978),
.B(n_954),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1062),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1057),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1065),
.A2(n_862),
.B1(n_943),
.B2(n_892),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1068),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1063),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_SL g1119 ( 
.A1(n_1098),
.A2(n_1009),
.B1(n_1042),
.B2(n_1004),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_SL g1120 ( 
.A1(n_1077),
.A2(n_905),
.B(n_903),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_1044),
.Y(n_1121)
);

AND2x4_ASAP7_75t_SL g1122 ( 
.A(n_1046),
.B(n_997),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1055),
.A2(n_871),
.B1(n_891),
.B2(n_875),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_1087),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1063),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1098),
.B(n_890),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1059),
.A2(n_871),
.B1(n_896),
.B2(n_904),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1093),
.A2(n_823),
.B1(n_998),
.B2(n_934),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_1047),
.Y(n_1129)
);

BUFx4f_ASAP7_75t_SL g1130 ( 
.A(n_1046),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1086),
.A2(n_1015),
.B1(n_1030),
.B2(n_1029),
.Y(n_1131)
);

INVx4_ASAP7_75t_L g1132 ( 
.A(n_1044),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1064),
.A2(n_911),
.B1(n_912),
.B2(n_904),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1054),
.B(n_886),
.Y(n_1134)
);

OAI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_1090),
.A2(n_905),
.B(n_903),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_SL g1136 ( 
.A1(n_1080),
.A2(n_998),
.B(n_854),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1067),
.A2(n_911),
.B1(n_912),
.B2(n_900),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1078),
.A2(n_916),
.B1(n_823),
.B2(n_910),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1069),
.A2(n_916),
.B1(n_910),
.B2(n_934),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1069),
.A2(n_1076),
.B1(n_1070),
.B2(n_1088),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1088),
.A2(n_934),
.B1(n_950),
.B2(n_883),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1066),
.A2(n_883),
.B1(n_936),
.B2(n_927),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1072),
.B(n_901),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1072),
.B(n_1024),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1047),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1074),
.A2(n_936),
.B1(n_870),
.B2(n_1024),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1052),
.B(n_1005),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1052),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1094),
.B(n_997),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1045),
.Y(n_1150)
);

BUFx4f_ASAP7_75t_SL g1151 ( 
.A(n_1074),
.Y(n_1151)
);

OAI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1071),
.A2(n_988),
.B1(n_997),
.B2(n_1029),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1089),
.A2(n_1029),
.B1(n_1030),
.B2(n_988),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1049),
.A2(n_870),
.B1(n_1008),
.B2(n_1005),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1045),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1050),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1097),
.A2(n_870),
.B1(n_1008),
.B2(n_1005),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1050),
.A2(n_1008),
.B1(n_1005),
.B2(n_937),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1073),
.B(n_1008),
.Y(n_1159)
);

OAI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_1061),
.A2(n_881),
.B(n_877),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1095),
.A2(n_944),
.B1(n_976),
.B2(n_1028),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1073),
.Y(n_1162)
);

INVx5_ASAP7_75t_L g1163 ( 
.A(n_1044),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1082),
.B(n_884),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1044),
.A2(n_976),
.B1(n_909),
.B2(n_884),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1061),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1082),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_1115),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1120),
.A2(n_1056),
.B1(n_958),
.B2(n_545),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1106),
.A2(n_1056),
.B1(n_1091),
.B2(n_1092),
.Y(n_1170)
);

OAI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1099),
.A2(n_1056),
.B1(n_1096),
.B2(n_1029),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1111),
.A2(n_1056),
.B1(n_1091),
.B2(n_1092),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1134),
.B(n_1056),
.Y(n_1173)
);

OAI221xp5_ASAP7_75t_L g1174 ( 
.A1(n_1135),
.A2(n_908),
.B1(n_889),
.B2(n_897),
.C(n_898),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1108),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1130),
.A2(n_1030),
.B1(n_1084),
.B2(n_1060),
.Y(n_1176)
);

OAI222xp33_ASAP7_75t_L g1177 ( 
.A1(n_1111),
.A2(n_1085),
.B1(n_1084),
.B2(n_1060),
.C1(n_984),
.C2(n_893),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1128),
.A2(n_909),
.B1(n_873),
.B2(n_893),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1112),
.A2(n_1084),
.B1(n_1085),
.B2(n_1060),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1143),
.B(n_1085),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_SL g1181 ( 
.A1(n_1130),
.A2(n_1030),
.B1(n_893),
.B2(n_873),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1101),
.A2(n_1126),
.B1(n_1149),
.B2(n_1138),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_L g1183 ( 
.A(n_1113),
.B(n_914),
.C(n_885),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1147),
.B(n_93),
.Y(n_1184)
);

OAI222xp33_ASAP7_75t_L g1185 ( 
.A1(n_1119),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.C1(n_35),
.C2(n_36),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1138),
.A2(n_873),
.B1(n_600),
.B2(n_567),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1144),
.A2(n_1116),
.B1(n_1151),
.B2(n_1109),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1116),
.B(n_873),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1151),
.A2(n_873),
.B1(n_600),
.B2(n_567),
.Y(n_1189)
);

OAI222xp33_ASAP7_75t_L g1190 ( 
.A1(n_1123),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.C1(n_37),
.C2(n_38),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1163),
.B(n_873),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_L g1192 ( 
.A(n_1123),
.B(n_567),
.C(n_565),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1146),
.A2(n_611),
.B1(n_610),
.B2(n_567),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1127),
.A2(n_873),
.B1(n_38),
.B2(n_39),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1110),
.A2(n_611),
.B1(n_610),
.B2(n_565),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1159),
.B(n_98),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1124),
.A2(n_611),
.B1(n_610),
.B2(n_565),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1114),
.B(n_99),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1102),
.B(n_37),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1146),
.A2(n_611),
.B1(n_610),
.B2(n_565),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1127),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1157),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1136),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1133),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1107),
.B(n_47),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1164),
.B(n_1145),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1100),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1163),
.B(n_100),
.Y(n_1208)
);

AOI222xp33_ASAP7_75t_L g1209 ( 
.A1(n_1133),
.A2(n_1137),
.B1(n_1141),
.B2(n_1129),
.C1(n_1140),
.C2(n_1166),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1118),
.Y(n_1210)
);

AND2x2_ASAP7_75t_SL g1211 ( 
.A(n_1140),
.B(n_50),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1125),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1137),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1141),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1121),
.B(n_101),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1104),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_1216)
);

OAI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_1160),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.C(n_60),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1167),
.B(n_59),
.Y(n_1218)
);

AOI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1142),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.C(n_64),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1121),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1157),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1148),
.B(n_103),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1152),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_1223)
);

OAI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1163),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1139),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1131),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1139),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_SL g1228 ( 
.A1(n_1163),
.A2(n_78),
.B1(n_105),
.B2(n_106),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1153),
.A2(n_78),
.B1(n_108),
.B2(n_109),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_L g1230 ( 
.A(n_1203),
.B(n_1161),
.C(n_1154),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1180),
.B(n_1162),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1168),
.B(n_1155),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1206),
.B(n_1161),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1173),
.B(n_1156),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1210),
.B(n_1150),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1212),
.B(n_1122),
.Y(n_1236)
);

AOI221xp5_ASAP7_75t_L g1237 ( 
.A1(n_1216),
.A2(n_1142),
.B1(n_1154),
.B2(n_1105),
.C(n_1158),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1175),
.B(n_1132),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_1216),
.B(n_1158),
.C(n_1132),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1199),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1211),
.A2(n_1165),
.B1(n_1117),
.B2(n_1103),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1182),
.B(n_1105),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1211),
.B(n_1103),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1177),
.A2(n_1165),
.B(n_1117),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_L g1245 ( 
.A(n_1217),
.B(n_110),
.C(n_112),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1171),
.B(n_113),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_L g1247 ( 
.A(n_1214),
.B(n_114),
.C(n_115),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1187),
.B(n_116),
.Y(n_1248)
);

OAI221xp5_ASAP7_75t_L g1249 ( 
.A1(n_1207),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.C(n_126),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1214),
.A2(n_127),
.B1(n_129),
.B2(n_134),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1219),
.B(n_135),
.C(n_138),
.Y(n_1251)
);

NOR3xp33_ASAP7_75t_L g1252 ( 
.A(n_1185),
.B(n_140),
.C(n_141),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1205),
.B(n_143),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1184),
.B(n_365),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1196),
.B(n_144),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1202),
.A2(n_145),
.B1(n_146),
.B2(n_150),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1170),
.A2(n_152),
.B(n_153),
.Y(n_1257)
);

OAI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_1220),
.A2(n_155),
.B(n_156),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1179),
.B(n_158),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1209),
.B(n_160),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1218),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1170),
.B(n_161),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1172),
.B(n_162),
.Y(n_1263)
);

AOI211xp5_ASAP7_75t_L g1264 ( 
.A1(n_1224),
.A2(n_1190),
.B(n_1221),
.C(n_1223),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1204),
.A2(n_164),
.B1(n_169),
.B2(n_170),
.Y(n_1265)
);

OAI21xp33_ASAP7_75t_L g1266 ( 
.A1(n_1227),
.A2(n_171),
.B(n_173),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1222),
.B(n_364),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1172),
.B(n_174),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1204),
.A2(n_175),
.B1(n_178),
.B2(n_182),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1227),
.B(n_1213),
.C(n_1226),
.Y(n_1270)
);

NAND4xp25_ASAP7_75t_L g1271 ( 
.A(n_1213),
.B(n_183),
.C(n_184),
.D(n_187),
.Y(n_1271)
);

OAI211xp5_ASAP7_75t_L g1272 ( 
.A1(n_1201),
.A2(n_190),
.B(n_191),
.C(n_193),
.Y(n_1272)
);

OAI221xp5_ASAP7_75t_L g1273 ( 
.A1(n_1201),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.C(n_197),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1198),
.B(n_198),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1229),
.A2(n_204),
.B(n_207),
.Y(n_1275)
);

NOR3xp33_ASAP7_75t_L g1276 ( 
.A(n_1228),
.B(n_208),
.C(n_209),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1231),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1252),
.A2(n_1194),
.B1(n_1225),
.B2(n_1188),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1270),
.A2(n_1194),
.B1(n_1169),
.B2(n_1178),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1240),
.B(n_1261),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1236),
.B(n_1215),
.Y(n_1281)
);

NOR2x1_ASAP7_75t_SL g1282 ( 
.A(n_1246),
.B(n_1191),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1232),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1245),
.B(n_1197),
.C(n_1208),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1238),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1234),
.B(n_1233),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1235),
.B(n_1192),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1243),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1242),
.B(n_1181),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1244),
.B(n_1183),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1246),
.B(n_1200),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1252),
.A2(n_1176),
.B1(n_1195),
.B2(n_1193),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1264),
.B(n_1186),
.C(n_1189),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_1253),
.Y(n_1294)
);

NAND4xp25_ASAP7_75t_L g1295 ( 
.A(n_1260),
.B(n_1174),
.C(n_211),
.D(n_212),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1268),
.A2(n_210),
.B(n_213),
.Y(n_1296)
);

NAND4xp75_ASAP7_75t_L g1297 ( 
.A(n_1257),
.B(n_1268),
.C(n_1259),
.D(n_1248),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1244),
.B(n_214),
.Y(n_1298)
);

AOI211xp5_ASAP7_75t_L g1299 ( 
.A1(n_1271),
.A2(n_219),
.B(n_220),
.C(n_221),
.Y(n_1299)
);

AO21x2_ASAP7_75t_L g1300 ( 
.A1(n_1262),
.A2(n_223),
.B(n_224),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1230),
.B(n_225),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1244),
.Y(n_1302)
);

AOI211xp5_ASAP7_75t_L g1303 ( 
.A1(n_1266),
.A2(n_229),
.B(n_231),
.C(n_232),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1241),
.B(n_1237),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1254),
.B(n_362),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1277),
.B(n_1283),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1302),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1280),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1288),
.B(n_1257),
.Y(n_1309)
);

NAND4xp75_ASAP7_75t_SL g1310 ( 
.A(n_1305),
.B(n_1282),
.C(n_1289),
.D(n_1297),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1296),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1286),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1285),
.B(n_1267),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1294),
.B(n_1263),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1290),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1295),
.A2(n_1276),
.B1(n_1275),
.B2(n_1247),
.Y(n_1316)
);

XOR2xp5_ASAP7_75t_L g1317 ( 
.A(n_1304),
.B(n_1255),
.Y(n_1317)
);

NAND4xp75_ASAP7_75t_L g1318 ( 
.A(n_1301),
.B(n_1274),
.C(n_1276),
.D(n_1249),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1287),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1281),
.B(n_1239),
.Y(n_1320)
);

XOR2x2_ASAP7_75t_L g1321 ( 
.A(n_1299),
.B(n_1303),
.Y(n_1321)
);

XOR2x2_ASAP7_75t_L g1322 ( 
.A(n_1299),
.B(n_1251),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1281),
.B(n_1256),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1298),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1300),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1324),
.Y(n_1326)
);

XNOR2xp5_ASAP7_75t_L g1327 ( 
.A(n_1310),
.B(n_1293),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1320),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1307),
.Y(n_1329)
);

XOR2x2_ASAP7_75t_L g1330 ( 
.A(n_1321),
.B(n_1279),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1324),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1316),
.A2(n_1278),
.B1(n_1303),
.B2(n_1292),
.Y(n_1332)
);

XOR2x2_ASAP7_75t_L g1333 ( 
.A(n_1321),
.B(n_1284),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1307),
.Y(n_1334)
);

XNOR2x1_ASAP7_75t_L g1335 ( 
.A(n_1317),
.B(n_1291),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1319),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1315),
.B(n_1300),
.Y(n_1337)
);

XOR2x2_ASAP7_75t_L g1338 ( 
.A(n_1322),
.B(n_1291),
.Y(n_1338)
);

XNOR2x2_ASAP7_75t_L g1339 ( 
.A(n_1322),
.B(n_1273),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1308),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1315),
.B(n_1296),
.Y(n_1341)
);

OA22x2_ASAP7_75t_L g1342 ( 
.A1(n_1327),
.A2(n_1311),
.B1(n_1323),
.B2(n_1313),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1329),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1340),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1329),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1326),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1336),
.Y(n_1347)
);

XNOR2xp5_ASAP7_75t_L g1348 ( 
.A(n_1333),
.B(n_1313),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1334),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1331),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1328),
.Y(n_1351)
);

CKINVDCx8_ASAP7_75t_R g1352 ( 
.A(n_1339),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1332),
.A2(n_1318),
.B1(n_1311),
.B2(n_1314),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1338),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1328),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1341),
.Y(n_1356)
);

OAI322xp33_ASAP7_75t_L g1357 ( 
.A1(n_1354),
.A2(n_1332),
.A3(n_1330),
.B1(n_1335),
.B2(n_1337),
.C1(n_1341),
.C2(n_1311),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1355),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1346),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1346),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1353),
.A2(n_1272),
.B1(n_1258),
.B2(n_1325),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1349),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1344),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1348),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1351),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1365),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1364),
.A2(n_1353),
.B1(n_1342),
.B2(n_1352),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1362),
.Y(n_1368)
);

AOI22x1_ASAP7_75t_L g1369 ( 
.A1(n_1357),
.A2(n_1351),
.B1(n_1349),
.B2(n_1345),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1359),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1358),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1371),
.Y(n_1372)
);

AO22x2_ASAP7_75t_L g1373 ( 
.A1(n_1366),
.A2(n_1363),
.B1(n_1343),
.B2(n_1360),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_SL g1374 ( 
.A1(n_1368),
.A2(n_1361),
.B(n_1356),
.C(n_1357),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1371),
.A2(n_1342),
.B1(n_1361),
.B2(n_1347),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1370),
.Y(n_1376)
);

INVxp33_ASAP7_75t_SL g1377 ( 
.A(n_1367),
.Y(n_1377)
);

OAI221xp5_ASAP7_75t_SL g1378 ( 
.A1(n_1375),
.A2(n_1369),
.B1(n_1337),
.B2(n_1250),
.C(n_1325),
.Y(n_1378)
);

NOR2xp67_ASAP7_75t_L g1379 ( 
.A(n_1372),
.B(n_1350),
.Y(n_1379)
);

AOI221xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1377),
.A2(n_1374),
.B1(n_1376),
.B2(n_1373),
.C(n_1309),
.Y(n_1380)
);

NOR4xp25_ASAP7_75t_L g1381 ( 
.A(n_1376),
.B(n_1250),
.C(n_1269),
.D(n_1265),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1377),
.B(n_1306),
.Y(n_1382)
);

AOI31xp33_ASAP7_75t_L g1383 ( 
.A1(n_1372),
.A2(n_1256),
.A3(n_1312),
.B(n_237),
.Y(n_1383)
);

OA22x2_ASAP7_75t_L g1384 ( 
.A1(n_1375),
.A2(n_233),
.B1(n_236),
.B2(n_238),
.Y(n_1384)
);

NOR2x1_ASAP7_75t_L g1385 ( 
.A(n_1376),
.B(n_241),
.Y(n_1385)
);

NOR2x1_ASAP7_75t_L g1386 ( 
.A(n_1385),
.B(n_245),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1380),
.B(n_1382),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1379),
.Y(n_1388)
);

NOR3xp33_ASAP7_75t_L g1389 ( 
.A(n_1378),
.B(n_247),
.C(n_248),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1384),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1381),
.A2(n_254),
.B1(n_256),
.B2(n_258),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1383),
.Y(n_1392)
);

AND4x1_ASAP7_75t_L g1393 ( 
.A(n_1386),
.B(n_259),
.C(n_265),
.D(n_266),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1388),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1391),
.B(n_356),
.Y(n_1395)
);

OA22x2_ASAP7_75t_L g1396 ( 
.A1(n_1387),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1392),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1389),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1390),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1397),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1393),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1394),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1399),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1393),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1396),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1398),
.A2(n_276),
.B1(n_278),
.B2(n_281),
.Y(n_1406)
);

OA22x2_ASAP7_75t_L g1407 ( 
.A1(n_1395),
.A2(n_282),
.B1(n_286),
.B2(n_287),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1397),
.Y(n_1408)
);

AOI31xp33_ASAP7_75t_L g1409 ( 
.A1(n_1401),
.A2(n_290),
.A3(n_293),
.B(n_294),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1403),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1402),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1404),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_SL g1413 ( 
.A1(n_1400),
.A2(n_302),
.B(n_303),
.C(n_305),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1405),
.A2(n_307),
.B1(n_308),
.B2(n_313),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1408),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1402),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1407),
.A2(n_1406),
.B1(n_318),
.B2(n_321),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1410),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1415),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1411),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1416),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1414),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1422),
.A2(n_1417),
.B1(n_1412),
.B2(n_1413),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1419),
.A2(n_1409),
.B1(n_322),
.B2(n_323),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1418),
.A2(n_314),
.B1(n_325),
.B2(n_326),
.Y(n_1425)
);

AO22x2_ASAP7_75t_L g1426 ( 
.A1(n_1420),
.A2(n_328),
.B1(n_331),
.B2(n_336),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1423),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1426),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1427),
.A2(n_1424),
.B1(n_1428),
.B2(n_1421),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1427),
.A2(n_1425),
.B1(n_343),
.B2(n_344),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1429),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1430),
.Y(n_1432)
);

AOI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1431),
.A2(n_342),
.B1(n_346),
.B2(n_347),
.C(n_348),
.Y(n_1433)
);

AOI211xp5_ASAP7_75t_L g1434 ( 
.A1(n_1433),
.A2(n_1432),
.B(n_349),
.C(n_351),
.Y(n_1434)
);


endmodule