module fake_ibex_1860_n_1507 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_224, n_183, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_68, n_117, n_214, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_228, n_1507);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_224;
input n_183;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;
input n_228;

output n_1507;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_242;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_235;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_234;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_262;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_257;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_252;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1504;
wire n_241;
wire n_1425;
wire n_231;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_236;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_291;
wire n_318;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1495;
wire n_303;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_255;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_270;
wire n_1340;
wire n_259;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_251;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_246;
wire n_922;
wire n_851;
wire n_993;
wire n_253;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1066;
wire n_245;
wire n_648;
wire n_571;
wire n_1169;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_839;
wire n_768;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_1057;
wire n_354;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_248;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_247;
wire n_1411;
wire n_237;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_232;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_249;
wire n_1443;
wire n_478;
wire n_239;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_243;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_244;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_1499;
wire n_1500;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_238;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_233;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_240;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_254;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

BUFx10_ASAP7_75t_L g231 ( 
.A(n_100),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_204),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_123),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_126),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_155),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_72),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_91),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_95),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_169),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_92),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_46),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_165),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_78),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_99),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_172),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_83),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_152),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_27),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_136),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_96),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_140),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_111),
.Y(n_256)
);

BUFx2_ASAP7_75t_SL g257 ( 
.A(n_170),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_132),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_156),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_23),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_90),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_182),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_124),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_112),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_89),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_217),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_159),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_191),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_168),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_30),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_87),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_102),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_121),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_27),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_85),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_230),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_45),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_127),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_37),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_154),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_56),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_207),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_178),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_63),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_26),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_43),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_122),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_29),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_173),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_135),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_66),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_116),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_40),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_138),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_82),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_53),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_23),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_209),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_158),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_143),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_7),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_36),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_221),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_125),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_141),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_113),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_215),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_212),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_29),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_57),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_210),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_32),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_97),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_194),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_119),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_38),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_157),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_105),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_76),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_223),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_183),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_208),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_64),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_37),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_79),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_61),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_216),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_8),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_161),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_190),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_227),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_181),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_188),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_93),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_225),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_206),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_171),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_219),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_68),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_81),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_133),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_192),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_150),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_24),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_86),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_8),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_201),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_16),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_69),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_51),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_197),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_151),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_163),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_106),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_153),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_7),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_52),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_14),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_98),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_88),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_15),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_71),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_146),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_179),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_222),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_94),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_130),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_118),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_25),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_166),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_107),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_50),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_16),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_55),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_35),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_129),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_147),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_202),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_120),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_195),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_13),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_128),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_22),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_164),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_167),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_84),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_175),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_211),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_160),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_43),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_24),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_131),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_47),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_15),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_6),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_20),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_214),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_142),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_114),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_196),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_26),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_203),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_148),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_137),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_117),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_218),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_0),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_34),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_189),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_224),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_186),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_115),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_36),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_30),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_241),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_393),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_265),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_245),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_236),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_240),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_267),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_267),
.Y(n_423)
);

BUFx8_ASAP7_75t_L g424 ( 
.A(n_313),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_231),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_231),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_278),
.B(n_0),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_265),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_245),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_267),
.Y(n_430)
);

INVx5_ASAP7_75t_L g431 ( 
.A(n_231),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_240),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_306),
.B(n_1),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_311),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_247),
.Y(n_436)
);

BUFx12f_ASAP7_75t_L g437 ( 
.A(n_247),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_384),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_278),
.A2(n_357),
.B1(n_294),
.B2(n_349),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_267),
.Y(n_440)
);

AOI22x1_ASAP7_75t_SL g441 ( 
.A1(n_394),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_2),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_296),
.B(n_62),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_333),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_260),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_247),
.B(n_3),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_275),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_302),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_267),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_289),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_251),
.B(n_4),
.Y(n_451)
);

BUFx12f_ASAP7_75t_L g452 ( 
.A(n_251),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g453 ( 
.A(n_252),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_281),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_251),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_296),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_281),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_297),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_330),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_340),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_281),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_351),
.B(n_5),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_330),
.Y(n_463)
);

BUFx8_ASAP7_75t_SL g464 ( 
.A(n_333),
.Y(n_464)
);

BUFx8_ASAP7_75t_SL g465 ( 
.A(n_344),
.Y(n_465)
);

BUFx8_ASAP7_75t_SL g466 ( 
.A(n_344),
.Y(n_466)
);

BUFx12f_ASAP7_75t_L g467 ( 
.A(n_340),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_361),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_267),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_271),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_361),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_359),
.B(n_5),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_373),
.Y(n_473)
);

BUFx8_ASAP7_75t_SL g474 ( 
.A(n_262),
.Y(n_474)
);

OAI22x1_ASAP7_75t_L g475 ( 
.A1(n_415),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_392),
.B(n_9),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_280),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_282),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_336),
.Y(n_479)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_361),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_361),
.Y(n_481)
);

NOR2x1_ASAP7_75t_L g482 ( 
.A(n_395),
.B(n_65),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_347),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_347),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_286),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_396),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_397),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_347),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_287),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_402),
.B(n_12),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_298),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_303),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_347),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_362),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_342),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_362),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_362),
.Y(n_497)
);

OAI22x1_ASAP7_75t_SL g498 ( 
.A1(n_310),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_498)
);

BUFx8_ASAP7_75t_L g499 ( 
.A(n_342),
.Y(n_499)
);

CKINVDCx6p67_ASAP7_75t_R g500 ( 
.A(n_250),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_414),
.B(n_17),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_362),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_234),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_263),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_234),
.Y(n_505)
);

NOR2x1_ASAP7_75t_L g506 ( 
.A(n_233),
.B(n_242),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_350),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_350),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_246),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_372),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_342),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_372),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_317),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_325),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_342),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_256),
.B(n_19),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_295),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_256),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_274),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_327),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_232),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_274),
.Y(n_522)
);

BUFx8_ASAP7_75t_L g523 ( 
.A(n_342),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_342),
.Y(n_524)
);

BUFx12f_ASAP7_75t_L g525 ( 
.A(n_329),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_279),
.A2(n_103),
.B(n_229),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_249),
.Y(n_527)
);

INVx6_ASAP7_75t_L g528 ( 
.A(n_257),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_253),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_279),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_288),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_419),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_507),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_474),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_R g535 ( 
.A(n_500),
.B(n_338),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_528),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_444),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_444),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_R g539 ( 
.A(n_453),
.B(n_446),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_474),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_R g541 ( 
.A(n_437),
.B(n_338),
.Y(n_541)
);

AOI21x1_ASAP7_75t_L g542 ( 
.A1(n_422),
.A2(n_308),
.B(n_288),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_419),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_464),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_464),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_465),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_432),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_477),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_466),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_507),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_466),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_R g552 ( 
.A(n_451),
.B(n_345),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_420),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_425),
.B(n_331),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_504),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_517),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_424),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_447),
.B(n_387),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_R g560 ( 
.A(n_452),
.B(n_467),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_507),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_525),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_470),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_514),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_521),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_521),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_477),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_439),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_478),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g570 ( 
.A(n_478),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_489),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_507),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_508),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_508),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_489),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_490),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_492),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_513),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_490),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_501),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_513),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_520),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_501),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_520),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_499),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_499),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_523),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_523),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_447),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_448),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_429),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_448),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_425),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_425),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_431),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_431),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_431),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_431),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_418),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_427),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_455),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_R g605 ( 
.A(n_436),
.B(n_356),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_441),
.B(n_360),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_455),
.B(n_235),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_426),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_528),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_485),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_R g611 ( 
.A(n_460),
.B(n_366),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_438),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_416),
.Y(n_613)
);

INVxp33_ASAP7_75t_L g614 ( 
.A(n_417),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_498),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_509),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_527),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_435),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_510),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_529),
.Y(n_620)
);

OA21x2_ASAP7_75t_L g621 ( 
.A1(n_422),
.A2(n_316),
.B(n_308),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_421),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_R g623 ( 
.A(n_443),
.B(n_367),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_519),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_510),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_433),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_433),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_519),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_518),
.B(n_266),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_512),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_456),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_R g632 ( 
.A(n_442),
.B(n_358),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_456),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_518),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_459),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_530),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_459),
.Y(n_637)
);

INVxp33_ASAP7_75t_SL g638 ( 
.A(n_434),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_418),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_506),
.B(n_269),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_512),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_463),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_463),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_479),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_512),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_530),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_R g647 ( 
.A(n_443),
.B(n_377),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_445),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_450),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_434),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_462),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_423),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_516),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_458),
.Y(n_654)
);

OA22x2_ASAP7_75t_L g655 ( 
.A1(n_475),
.A2(n_370),
.B1(n_375),
.B2(n_374),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_418),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_473),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_486),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_472),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_487),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_476),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_R g662 ( 
.A(n_443),
.B(n_380),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_449),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_469),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_511),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_502),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_R g667 ( 
.A(n_443),
.B(n_376),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_430),
.B(n_382),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_418),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_440),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_R g671 ( 
.A(n_493),
.B(n_408),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_526),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_428),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_440),
.Y(n_674)
);

NOR2x1p5_ASAP7_75t_L g675 ( 
.A(n_493),
.B(n_409),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_495),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_495),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_515),
.B(n_237),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_515),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_524),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_524),
.B(n_363),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_522),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_522),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_R g684 ( 
.A(n_494),
.B(n_238),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_502),
.B(n_272),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_522),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_483),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_531),
.Y(n_688)
);

CKINVDCx16_ASAP7_75t_R g689 ( 
.A(n_482),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_531),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_531),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_R g692 ( 
.A(n_494),
.B(n_243),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_R g693 ( 
.A(n_531),
.B(n_244),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_480),
.Y(n_694)
);

CKINVDCx16_ASAP7_75t_R g695 ( 
.A(n_484),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_480),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_480),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_484),
.Y(n_698)
);

AND2x2_ASAP7_75t_SL g699 ( 
.A(n_570),
.B(n_273),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_653),
.B(n_276),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_638),
.B(n_239),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_659),
.B(n_283),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_532),
.Y(n_703)
);

INVx8_ASAP7_75t_L g704 ( 
.A(n_622),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_543),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_640),
.B(n_668),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_547),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_675),
.B(n_300),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_536),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_614),
.B(n_277),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_648),
.B(n_305),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_649),
.B(n_307),
.Y(n_712)
);

NOR3xp33_ASAP7_75t_L g713 ( 
.A(n_592),
.B(n_595),
.C(n_593),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_646),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_569),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_559),
.B(n_624),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_661),
.B(n_314),
.C(n_312),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_553),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_565),
.B(n_248),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_628),
.B(n_254),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_635),
.B(n_255),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_646),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_L g723 ( 
.A(n_562),
.B(n_20),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_654),
.B(n_319),
.C(n_315),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_616),
.B(n_258),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_617),
.B(n_259),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_621),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_620),
.B(n_261),
.Y(n_728)
);

NOR2xp67_ASAP7_75t_L g729 ( 
.A(n_563),
.B(n_21),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_566),
.B(n_264),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_657),
.B(n_268),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_658),
.B(n_270),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_660),
.B(n_324),
.C(n_320),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_SL g734 ( 
.A(n_672),
.B(n_284),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_618),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_533),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_L g737 ( 
.A(n_667),
.B(n_285),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_650),
.B(n_337),
.C(n_334),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_631),
.B(n_290),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_SL g740 ( 
.A(n_535),
.B(n_291),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_633),
.B(n_292),
.Y(n_741)
);

BUFx6f_ASAP7_75t_SL g742 ( 
.A(n_558),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_576),
.B(n_582),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_634),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_550),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_583),
.B(n_346),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_561),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_586),
.B(n_348),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_674),
.B(n_352),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_594),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_572),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_573),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_642),
.B(n_293),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_676),
.B(n_354),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_548),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_636),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_629),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_608),
.B(n_299),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_677),
.B(n_365),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_574),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_685),
.Y(n_761)
);

NOR3xp33_ASAP7_75t_L g762 ( 
.A(n_612),
.B(n_578),
.C(n_689),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_679),
.B(n_371),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_567),
.B(n_21),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_609),
.B(n_301),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_663),
.B(n_379),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_552),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_623),
.B(n_304),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_665),
.B(n_643),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_644),
.B(n_309),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_681),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_577),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_L g773 ( 
.A1(n_539),
.A2(n_381),
.B1(n_383),
.B2(n_386),
.Y(n_773)
);

INVxp33_ASAP7_75t_L g774 ( 
.A(n_560),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_581),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_575),
.B(n_25),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_619),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_L g778 ( 
.A(n_632),
.B(n_390),
.C(n_388),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_623),
.B(n_318),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_564),
.B(n_321),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_596),
.B(n_322),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_647),
.B(n_323),
.Y(n_782)
);

NOR2x1p5_ASAP7_75t_L g783 ( 
.A(n_534),
.B(n_326),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_680),
.B(n_405),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_579),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_L g786 ( 
.A(n_580),
.B(n_413),
.C(n_410),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_647),
.B(n_328),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_625),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_630),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_672),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_585),
.B(n_28),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_597),
.B(n_332),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_626),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_598),
.B(n_335),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_599),
.B(n_339),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_600),
.B(n_341),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_641),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_542),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_664),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_687),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_601),
.B(n_343),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_645),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_587),
.B(n_615),
.C(n_556),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_698),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_655),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_651),
.B(n_353),
.Y(n_806)
);

INVxp33_ASAP7_75t_L g807 ( 
.A(n_560),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_682),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_555),
.B(n_355),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_554),
.B(n_28),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_683),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_686),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_688),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_695),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_652),
.B(n_364),
.Y(n_815)
);

BUFx5_ASAP7_75t_L g816 ( 
.A(n_662),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_691),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_670),
.B(n_368),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_678),
.B(n_369),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_690),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_588),
.B(n_378),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_697),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_604),
.B(n_385),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_589),
.B(n_591),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_541),
.B(n_389),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_694),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_666),
.Y(n_827)
);

XOR2xp5_ASAP7_75t_L g828 ( 
.A(n_537),
.B(n_538),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_607),
.B(n_398),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_696),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_671),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_632),
.B(n_400),
.C(n_399),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_627),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_602),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_637),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_692),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_541),
.B(n_401),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_535),
.B(n_404),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_603),
.B(n_406),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_602),
.Y(n_840)
);

NOR3xp33_ASAP7_75t_L g841 ( 
.A(n_557),
.B(n_411),
.C(n_407),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_708),
.B(n_590),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_715),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_750),
.Y(n_844)
);

NOR2x1_ASAP7_75t_L g845 ( 
.A(n_832),
.B(n_571),
.Y(n_845)
);

INVx5_ASAP7_75t_L g846 ( 
.A(n_790),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_704),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_703),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_705),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_707),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_793),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_714),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_755),
.B(n_584),
.Y(n_853)
);

NOR2x1p5_ASAP7_75t_L g854 ( 
.A(n_764),
.B(n_540),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_785),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_713),
.B(n_605),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_708),
.B(n_568),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_706),
.B(n_611),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_804),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_699),
.B(n_611),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_702),
.B(n_412),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_718),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_722),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_798),
.A2(n_639),
.B(n_602),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_833),
.B(n_544),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_704),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_735),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_734),
.B(n_684),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_799),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_756),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_790),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_805),
.A2(n_610),
.B1(n_684),
.B2(n_693),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_822),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_839),
.B(n_546),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_700),
.B(n_31),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_800),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_816),
.B(n_549),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_SL g878 ( 
.A1(n_828),
.A2(n_545),
.B1(n_551),
.B2(n_606),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_744),
.Y(n_879)
);

OR2x6_ASAP7_75t_L g880 ( 
.A(n_704),
.B(n_484),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_826),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_743),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_709),
.B(n_32),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_743),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_716),
.B(n_33),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_814),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_784),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_R g888 ( 
.A(n_740),
.B(n_33),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_SL g889 ( 
.A1(n_776),
.A2(n_488),
.B1(n_496),
.B2(n_497),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_727),
.A2(n_673),
.B(n_669),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_809),
.Y(n_891)
);

AND3x1_ASAP7_75t_L g892 ( 
.A(n_803),
.B(n_39),
.C(n_41),
.Y(n_892)
);

AND2x6_ASAP7_75t_SL g893 ( 
.A(n_742),
.B(n_39),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_736),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_771),
.A2(n_488),
.B1(n_496),
.B2(n_497),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_786),
.A2(n_488),
.B1(n_496),
.B2(n_497),
.Y(n_896)
);

INVxp67_ASAP7_75t_SL g897 ( 
.A(n_820),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_830),
.Y(n_898)
);

INVxp33_ASAP7_75t_L g899 ( 
.A(n_806),
.Y(n_899)
);

AND2x4_ASAP7_75t_SL g900 ( 
.A(n_835),
.B(n_497),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_749),
.B(n_42),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_824),
.Y(n_902)
);

INVx3_ASAP7_75t_SL g903 ( 
.A(n_810),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_710),
.B(n_44),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_711),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_711),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_745),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_712),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_749),
.B(n_45),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_778),
.B(n_67),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_SL g911 ( 
.A1(n_827),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_754),
.B(n_48),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_762),
.B(n_49),
.Y(n_913)
);

HB1xp67_ASAP7_75t_SL g914 ( 
.A(n_742),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_802),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_809),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_791),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_767),
.B(n_49),
.Y(n_918)
);

INVx8_ASAP7_75t_L g919 ( 
.A(n_825),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_746),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_729),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_748),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_816),
.B(n_428),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_757),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_754),
.B(n_759),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_759),
.B(n_51),
.Y(n_926)
);

NOR2x1p5_ASAP7_75t_L g927 ( 
.A(n_769),
.B(n_52),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_780),
.B(n_53),
.Y(n_928)
);

BUFx8_ASAP7_75t_L g929 ( 
.A(n_831),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_761),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_783),
.B(n_54),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_763),
.B(n_55),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_747),
.Y(n_933)
);

BUFx4f_ASAP7_75t_L g934 ( 
.A(n_836),
.Y(n_934)
);

OR2x6_ASAP7_75t_L g935 ( 
.A(n_723),
.B(n_56),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_701),
.B(n_57),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_751),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_773),
.A2(n_471),
.B1(n_454),
.B2(n_457),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_766),
.B(n_58),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_841),
.B(n_58),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_766),
.B(n_59),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_725),
.B(n_59),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_738),
.A2(n_471),
.B1(n_454),
.B2(n_457),
.Y(n_943)
);

OR2x6_ASAP7_75t_L g944 ( 
.A(n_838),
.B(n_837),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_815),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_717),
.B(n_60),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_815),
.Y(n_947)
);

BUFx4f_ASAP7_75t_L g948 ( 
.A(n_808),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_818),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_752),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_811),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_812),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_813),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_R g954 ( 
.A(n_821),
.B(n_61),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_760),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_818),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_819),
.A2(n_733),
.B(n_724),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_772),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_768),
.A2(n_461),
.B1(n_468),
.B2(n_481),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_817),
.Y(n_960)
);

NOR2x1p5_ASAP7_75t_L g961 ( 
.A(n_837),
.B(n_726),
.Y(n_961)
);

INVx8_ASAP7_75t_L g962 ( 
.A(n_774),
.Y(n_962)
);

AND2x6_ASAP7_75t_L g963 ( 
.A(n_721),
.B(n_481),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_775),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_777),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_SL g966 ( 
.A1(n_807),
.A2(n_732),
.B1(n_728),
.B2(n_731),
.Y(n_966)
);

CKINVDCx16_ASAP7_75t_R g967 ( 
.A(n_758),
.Y(n_967)
);

AND2x4_ASAP7_75t_SL g968 ( 
.A(n_765),
.B(n_639),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_788),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_925),
.B(n_882),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_853),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_855),
.Y(n_972)
);

NOR2x1_ASAP7_75t_L g973 ( 
.A(n_931),
.B(n_779),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_884),
.B(n_719),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_SL g975 ( 
.A1(n_942),
.A2(n_730),
.B(n_829),
.C(n_737),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_945),
.A2(n_787),
.B(n_782),
.C(n_720),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_905),
.A2(n_823),
.B1(n_781),
.B2(n_795),
.Y(n_977)
);

AO32x1_ASAP7_75t_L g978 ( 
.A1(n_904),
.A2(n_840),
.A3(n_834),
.B1(n_789),
.B2(n_797),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_844),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_906),
.B(n_792),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_846),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_908),
.B(n_739),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_947),
.A2(n_770),
.B(n_741),
.C(n_753),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_848),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_849),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_850),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_887),
.A2(n_796),
.B1(n_794),
.B2(n_801),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_859),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_851),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_914),
.B(n_70),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_SL g991 ( 
.A(n_954),
.B(n_73),
.C(n_74),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_857),
.B(n_75),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_843),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_883),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_SL g995 ( 
.A(n_967),
.B(n_77),
.C(n_80),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_883),
.B(n_656),
.Y(n_996)
);

INVx5_ASAP7_75t_L g997 ( 
.A(n_880),
.Y(n_997)
);

INVx5_ASAP7_75t_L g998 ( 
.A(n_880),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_920),
.B(n_922),
.Y(n_999)
);

INVx5_ASAP7_75t_L g1000 ( 
.A(n_931),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_901),
.A2(n_912),
.B(n_926),
.C(n_909),
.Y(n_1001)
);

AOI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_899),
.A2(n_858),
.B(n_874),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_862),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_SL g1004 ( 
.A1(n_885),
.A2(n_101),
.B(n_104),
.C(n_108),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_847),
.Y(n_1005)
);

OR2x6_ASAP7_75t_SL g1006 ( 
.A(n_878),
.B(n_109),
.Y(n_1006)
);

NOR2xp67_ASAP7_75t_L g1007 ( 
.A(n_865),
.B(n_110),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_886),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_917),
.B(n_134),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_957),
.A2(n_139),
.B(n_144),
.C(n_145),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_857),
.B(n_149),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_869),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_866),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_879),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_867),
.Y(n_1015)
);

OA21x2_ASAP7_75t_L g1016 ( 
.A1(n_890),
.A2(n_174),
.B(n_176),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_932),
.A2(n_939),
.B(n_941),
.C(n_875),
.Y(n_1017)
);

OAI21xp33_ASAP7_75t_SL g1018 ( 
.A1(n_927),
.A2(n_180),
.B(n_184),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_846),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_SL g1020 ( 
.A(n_902),
.B(n_185),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_SL g1021 ( 
.A(n_967),
.B(n_198),
.C(n_199),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_842),
.B(n_200),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_870),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_842),
.B(n_903),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_846),
.Y(n_1025)
);

AND2x4_ASAP7_75t_SL g1026 ( 
.A(n_935),
.B(n_205),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_888),
.B(n_220),
.Y(n_1027)
);

BUFx10_ASAP7_75t_L g1028 ( 
.A(n_893),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_946),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_860),
.B(n_226),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_891),
.B(n_228),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_876),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_916),
.B(n_966),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_966),
.B(n_919),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_861),
.B(n_961),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_961),
.B(n_936),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_913),
.B(n_856),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_872),
.B(n_928),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_944),
.B(n_881),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_919),
.B(n_871),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_872),
.B(n_940),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_946),
.A2(n_918),
.B(n_897),
.C(n_930),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_871),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_940),
.A2(n_845),
.B1(n_854),
.B2(n_927),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_929),
.Y(n_1045)
);

NOR3xp33_ASAP7_75t_SL g1046 ( 
.A(n_911),
.B(n_924),
.C(n_877),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_910),
.A2(n_938),
.B(n_953),
.C(n_934),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_871),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_852),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_935),
.A2(n_868),
.B(n_921),
.C(n_953),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_952),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_863),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_934),
.A2(n_896),
.B(n_898),
.C(n_881),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_898),
.B(n_960),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_960),
.B(n_944),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_962),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_894),
.A2(n_969),
.B(n_958),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_963),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_873),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_951),
.B(n_873),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_951),
.B(n_952),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_962),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_965),
.A2(n_933),
.B(n_964),
.C(n_937),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_948),
.B(n_854),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_915),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_948),
.B(n_929),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_907),
.A2(n_955),
.B(n_950),
.Y(n_1067)
);

BUFx12f_ASAP7_75t_L g1068 ( 
.A(n_963),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_900),
.Y(n_1069)
);

AO32x1_ASAP7_75t_L g1070 ( 
.A1(n_968),
.A2(n_892),
.A3(n_911),
.B1(n_889),
.B2(n_963),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_943),
.A2(n_959),
.B(n_895),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_895),
.A2(n_947),
.B(n_945),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_851),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_925),
.B(n_882),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_SL g1075 ( 
.A(n_954),
.B(n_540),
.C(n_534),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_853),
.B(n_559),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_869),
.Y(n_1077)
);

AOI21x1_ASAP7_75t_L g1078 ( 
.A1(n_890),
.A2(n_864),
.B(n_923),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_945),
.A2(n_947),
.B(n_956),
.C(n_949),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_925),
.B(n_882),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_853),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_945),
.A2(n_947),
.B(n_956),
.C(n_949),
.Y(n_1082)
);

AO32x2_ASAP7_75t_L g1083 ( 
.A1(n_966),
.A2(n_911),
.A3(n_960),
.B1(n_503),
.B2(n_505),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_853),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_855),
.B(n_755),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_846),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_846),
.Y(n_1087)
);

NOR2x1_ASAP7_75t_R g1088 ( 
.A(n_843),
.B(n_534),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_925),
.B(n_882),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_857),
.B(n_570),
.Y(n_1090)
);

BUFx4f_ASAP7_75t_L g1091 ( 
.A(n_931),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_853),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_SL g1093 ( 
.A1(n_931),
.A2(n_715),
.B1(n_444),
.B2(n_538),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_925),
.B(n_882),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_R g1095 ( 
.A(n_914),
.B(n_715),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_846),
.Y(n_1096)
);

OAI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_925),
.A2(n_593),
.B(n_592),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_945),
.A2(n_947),
.B(n_956),
.C(n_949),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_857),
.B(n_570),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_853),
.B(n_559),
.Y(n_1100)
);

AOI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_925),
.A2(n_439),
.B1(n_614),
.B2(n_773),
.C(n_613),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_853),
.B(n_559),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_SL g1103 ( 
.A(n_888),
.B(n_715),
.C(n_444),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_844),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_945),
.A2(n_947),
.B(n_956),
.C(n_949),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_844),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_847),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_855),
.B(n_755),
.Y(n_1108)
);

BUFx12f_ASAP7_75t_L g1109 ( 
.A(n_1045),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1041),
.A2(n_1091),
.B1(n_1038),
.B2(n_1033),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_997),
.B(n_998),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_SL g1112 ( 
.A1(n_1050),
.A2(n_1074),
.B(n_970),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1080),
.B(n_1089),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1079),
.A2(n_1098),
.B(n_1082),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_979),
.Y(n_1115)
);

NAND2x1_ASAP7_75t_L g1116 ( 
.A(n_981),
.B(n_1019),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1094),
.B(n_1000),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1012),
.Y(n_1118)
);

INVx8_ASAP7_75t_L g1119 ( 
.A(n_997),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1077),
.Y(n_1120)
);

AO21x2_ASAP7_75t_L g1121 ( 
.A1(n_1047),
.A2(n_1078),
.B(n_1071),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_981),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_1093),
.B(n_1064),
.Y(n_1123)
);

BUFx10_ASAP7_75t_L g1124 ( 
.A(n_1026),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_997),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1019),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1076),
.B(n_1100),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_984),
.Y(n_1128)
);

INVxp67_ASAP7_75t_SL g1129 ( 
.A(n_1065),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_1004),
.A2(n_1001),
.B(n_1017),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1000),
.B(n_1105),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1008),
.B(n_972),
.Y(n_1132)
);

AO21x2_ASAP7_75t_L g1133 ( 
.A1(n_1053),
.A2(n_1010),
.B(n_1072),
.Y(n_1133)
);

INVxp67_ASAP7_75t_SL g1134 ( 
.A(n_1065),
.Y(n_1134)
);

AND2x6_ASAP7_75t_L g1135 ( 
.A(n_1019),
.B(n_1025),
.Y(n_1135)
);

NAND2x1_ASAP7_75t_L g1136 ( 
.A(n_1025),
.B(n_1043),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1095),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1025),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1097),
.B(n_1102),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_1043),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_971),
.B(n_1081),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_1065),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1043),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_1048),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_985),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_988),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1000),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_986),
.Y(n_1148)
);

BUFx2_ASAP7_75t_SL g1149 ( 
.A(n_998),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_999),
.A2(n_974),
.B(n_1035),
.Y(n_1150)
);

BUFx4_ASAP7_75t_SL g1151 ( 
.A(n_1107),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1048),
.Y(n_1152)
);

OR2x6_ASAP7_75t_L g1153 ( 
.A(n_1068),
.B(n_989),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1032),
.Y(n_1154)
);

NAND2x1p5_ASAP7_75t_L g1155 ( 
.A(n_998),
.B(n_1086),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_990),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1003),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1086),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_SL g1159 ( 
.A(n_993),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1086),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1101),
.B(n_1014),
.Y(n_1161)
);

BUFx2_ASAP7_75t_SL g1162 ( 
.A(n_1073),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_1084),
.Y(n_1163)
);

CKINVDCx11_ASAP7_75t_R g1164 ( 
.A(n_1006),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1023),
.B(n_1015),
.Y(n_1165)
);

INVxp67_ASAP7_75t_SL g1166 ( 
.A(n_1029),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_1087),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1092),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1087),
.B(n_1096),
.Y(n_1169)
);

BUFx2_ASAP7_75t_R g1170 ( 
.A(n_1085),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1028),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1104),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_1096),
.B(n_1058),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1096),
.Y(n_1174)
);

BUFx2_ASAP7_75t_SL g1175 ( 
.A(n_1056),
.Y(n_1175)
);

NAND2x1p5_ASAP7_75t_L g1176 ( 
.A(n_1058),
.B(n_1069),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_1058),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1106),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_977),
.A2(n_1042),
.B(n_1036),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1049),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_1061),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1052),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1016),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_1062),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_987),
.A2(n_982),
.B(n_976),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1005),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1037),
.B(n_994),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_980),
.A2(n_1067),
.B(n_1057),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1039),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1002),
.B(n_1044),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1034),
.A2(n_1103),
.B1(n_973),
.B2(n_992),
.Y(n_1191)
);

INVxp67_ASAP7_75t_SL g1192 ( 
.A(n_996),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1039),
.B(n_1011),
.Y(n_1193)
);

INVx6_ASAP7_75t_SL g1194 ( 
.A(n_1028),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1051),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1059),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1013),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1060),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1083),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1083),
.Y(n_1200)
);

BUFx2_ASAP7_75t_SL g1201 ( 
.A(n_1108),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1054),
.Y(n_1202)
);

AOI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1007),
.A2(n_1030),
.B(n_1027),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_978),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1055),
.B(n_983),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_1088),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_1063),
.A2(n_995),
.B(n_1021),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1040),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1090),
.B(n_1099),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1083),
.Y(n_1210)
);

INVxp67_ASAP7_75t_SL g1211 ( 
.A(n_1020),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_1075),
.Y(n_1212)
);

BUFx5_ASAP7_75t_L g1213 ( 
.A(n_1009),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1046),
.B(n_1022),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1024),
.B(n_1066),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_991),
.B(n_1031),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1018),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1070),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1070),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_975),
.B(n_1097),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_981),
.Y(n_1221)
);

AO21x1_ASAP7_75t_SL g1222 ( 
.A1(n_1217),
.A2(n_1114),
.B(n_1113),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1115),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1132),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1151),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1129),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1128),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1211),
.A2(n_1110),
.B1(n_1139),
.B2(n_1156),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1145),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1148),
.Y(n_1230)
);

NOR2x1_ASAP7_75t_R g1231 ( 
.A(n_1206),
.B(n_1164),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_1119),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1211),
.A2(n_1110),
.B1(n_1139),
.B2(n_1156),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1157),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_1151),
.Y(n_1235)
);

AOI222xp33_ASAP7_75t_L g1236 ( 
.A1(n_1164),
.A2(n_1127),
.B1(n_1161),
.B2(n_1191),
.C1(n_1179),
.C2(n_1190),
.Y(n_1236)
);

BUFx8_ASAP7_75t_SL g1237 ( 
.A(n_1109),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1131),
.B(n_1178),
.Y(n_1238)
);

CKINVDCx11_ASAP7_75t_R g1239 ( 
.A(n_1124),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1178),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1120),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1172),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1120),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1165),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1165),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1180),
.Y(n_1246)
);

BUFx4f_ASAP7_75t_SL g1247 ( 
.A(n_1194),
.Y(n_1247)
);

INVx8_ASAP7_75t_L g1248 ( 
.A(n_1119),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1119),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1182),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1135),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_1137),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1129),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1118),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1191),
.A2(n_1193),
.B1(n_1117),
.B2(n_1123),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1123),
.A2(n_1216),
.B1(n_1209),
.B2(n_1214),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1154),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1123),
.A2(n_1112),
.B1(n_1117),
.B2(n_1131),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1134),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1134),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1187),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1146),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1196),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1141),
.A2(n_1185),
.B1(n_1215),
.B2(n_1218),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1135),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1159),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1212),
.Y(n_1267)
);

AOI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1183),
.A2(n_1217),
.B(n_1204),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1166),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1141),
.A2(n_1215),
.B1(n_1218),
.B2(n_1205),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1220),
.A2(n_1168),
.B1(n_1163),
.B2(n_1219),
.Y(n_1271)
);

BUFx2_ASAP7_75t_R g1272 ( 
.A(n_1171),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1220),
.A2(n_1219),
.B1(n_1202),
.B2(n_1201),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1166),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1124),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1204),
.A2(n_1210),
.B(n_1200),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1199),
.Y(n_1277)
);

CKINVDCx11_ASAP7_75t_R g1278 ( 
.A(n_1212),
.Y(n_1278)
);

NAND2x1p5_ASAP7_75t_L g1279 ( 
.A(n_1177),
.B(n_1184),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1195),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1142),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1135),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1177),
.B(n_1184),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1197),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1219),
.A2(n_1202),
.B1(n_1150),
.B2(n_1198),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1195),
.Y(n_1286)
);

CKINVDCx16_ASAP7_75t_R g1287 ( 
.A(n_1225),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1284),
.B(n_1197),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1248),
.Y(n_1289)
);

INVx4_ASAP7_75t_SL g1290 ( 
.A(n_1249),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1261),
.B(n_1160),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1224),
.B(n_1181),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1223),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1227),
.B(n_1189),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1240),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1226),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1232),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_R g1298 ( 
.A(n_1247),
.B(n_1159),
.Y(n_1298)
);

CKINVDCx16_ASAP7_75t_R g1299 ( 
.A(n_1235),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1229),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1264),
.A2(n_1188),
.B(n_1192),
.Y(n_1301)
);

NAND2xp33_ASAP7_75t_R g1302 ( 
.A(n_1226),
.B(n_1207),
.Y(n_1302)
);

NOR2xp67_ASAP7_75t_L g1303 ( 
.A(n_1232),
.B(n_1219),
.Y(n_1303)
);

BUFx4f_ASAP7_75t_SL g1304 ( 
.A(n_1232),
.Y(n_1304)
);

CKINVDCx16_ASAP7_75t_R g1305 ( 
.A(n_1252),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1255),
.A2(n_1213),
.B1(n_1149),
.B2(n_1147),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1230),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1234),
.B(n_1189),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1244),
.B(n_1170),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1242),
.B(n_1198),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1249),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1248),
.A2(n_1208),
.B(n_1125),
.C(n_1181),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1253),
.Y(n_1313)
);

NAND2xp33_ASAP7_75t_R g1314 ( 
.A(n_1231),
.B(n_1153),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1245),
.B(n_1125),
.Y(n_1315)
);

INVx4_ASAP7_75t_SL g1316 ( 
.A(n_1249),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1241),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1280),
.B(n_1186),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1241),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1228),
.A2(n_1213),
.B1(n_1207),
.B2(n_1192),
.Y(n_1320)
);

NAND2xp33_ASAP7_75t_R g1321 ( 
.A(n_1253),
.B(n_1207),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1263),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1236),
.B(n_1246),
.Y(n_1323)
);

NAND4xp25_ASAP7_75t_L g1324 ( 
.A(n_1256),
.B(n_1186),
.C(n_1138),
.D(n_1140),
.Y(n_1324)
);

CKINVDCx16_ASAP7_75t_R g1325 ( 
.A(n_1252),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1286),
.B(n_1221),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_R g1327 ( 
.A(n_1248),
.B(n_1239),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1250),
.B(n_1152),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1269),
.B(n_1175),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1274),
.B(n_1152),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_1266),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_R g1332 ( 
.A(n_1248),
.B(n_1239),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1270),
.A2(n_1203),
.B(n_1111),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1254),
.B(n_1138),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1259),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1233),
.A2(n_1213),
.B1(n_1130),
.B2(n_1133),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1262),
.B(n_1249),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_SL g1338 ( 
.A1(n_1258),
.A2(n_1275),
.B(n_1273),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1243),
.Y(n_1339)
);

INVxp67_ASAP7_75t_SL g1340 ( 
.A(n_1259),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1296),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1313),
.B(n_1277),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1313),
.B(n_1222),
.Y(n_1343)
);

INVx5_ASAP7_75t_L g1344 ( 
.A(n_1297),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1335),
.B(n_1222),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1335),
.B(n_1276),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1317),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1323),
.A2(n_1238),
.B1(n_1278),
.B2(n_1130),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1295),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1304),
.Y(n_1350)
);

INVxp33_ASAP7_75t_L g1351 ( 
.A(n_1327),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1293),
.B(n_1300),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1340),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1288),
.B(n_1260),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1319),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1307),
.B(n_1238),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1339),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1322),
.Y(n_1358)
);

INVx5_ASAP7_75t_L g1359 ( 
.A(n_1311),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1301),
.B(n_1276),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1336),
.B(n_1260),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1306),
.B(n_1271),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1336),
.B(n_1281),
.Y(n_1363)
);

OAI222xp33_ASAP7_75t_L g1364 ( 
.A1(n_1306),
.A2(n_1281),
.B1(n_1285),
.B2(n_1283),
.C1(n_1279),
.C2(n_1111),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1304),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1330),
.B(n_1257),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1360),
.B(n_1268),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1358),
.B(n_1292),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1352),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1348),
.B(n_1337),
.C(n_1333),
.Y(n_1370)
);

NAND3xp33_ASAP7_75t_L g1371 ( 
.A(n_1348),
.B(n_1337),
.C(n_1320),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1353),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1354),
.B(n_1310),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1343),
.B(n_1303),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1347),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1352),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1360),
.B(n_1121),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1354),
.B(n_1357),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1353),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1357),
.B(n_1329),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1346),
.B(n_1121),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1355),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1358),
.B(n_1318),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1355),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1349),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1369),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1381),
.B(n_1361),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1376),
.B(n_1342),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1378),
.B(n_1341),
.Y(n_1389)
);

INVxp67_ASAP7_75t_SL g1390 ( 
.A(n_1382),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1381),
.B(n_1361),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1385),
.Y(n_1392)
);

OAI221xp5_ASAP7_75t_L g1393 ( 
.A1(n_1370),
.A2(n_1371),
.B1(n_1314),
.B2(n_1362),
.C(n_1365),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1375),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1384),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1383),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1374),
.B(n_1343),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1378),
.B(n_1341),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1375),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1368),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1372),
.B(n_1342),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1373),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1377),
.B(n_1363),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1377),
.B(n_1363),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1385),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1395),
.B(n_1379),
.Y(n_1406)
);

OA222x2_ASAP7_75t_L g1407 ( 
.A1(n_1389),
.A2(n_1380),
.B1(n_1373),
.B2(n_1289),
.C1(n_1362),
.C2(n_1351),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1390),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1389),
.Y(n_1409)
);

OAI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1393),
.A2(n_1344),
.B1(n_1350),
.B2(n_1365),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1397),
.A2(n_1364),
.B(n_1365),
.Y(n_1411)
);

NAND4xp75_ASAP7_75t_SL g1412 ( 
.A(n_1403),
.B(n_1309),
.C(n_1345),
.D(n_1332),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1402),
.A2(n_1400),
.B1(n_1396),
.B2(n_1397),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1387),
.B(n_1367),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1398),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_SL g1416 ( 
.A(n_1397),
.B(n_1350),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1394),
.B(n_1344),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1398),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1386),
.B(n_1350),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1401),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1403),
.B(n_1367),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1392),
.Y(n_1422)
);

AO22x1_ASAP7_75t_L g1423 ( 
.A1(n_1407),
.A2(n_1350),
.B1(n_1344),
.B2(n_1374),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1416),
.A2(n_1299),
.B1(n_1287),
.B2(n_1344),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1418),
.B(n_1409),
.Y(n_1425)
);

OAI211xp5_ASAP7_75t_L g1426 ( 
.A1(n_1411),
.A2(n_1298),
.B(n_1278),
.C(n_1309),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1415),
.B(n_1404),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1408),
.A2(n_1364),
.B(n_1312),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1422),
.Y(n_1429)
);

AO22x1_ASAP7_75t_L g1430 ( 
.A1(n_1412),
.A2(n_1344),
.B1(n_1374),
.B2(n_1359),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1422),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1413),
.A2(n_1414),
.B(n_1417),
.C(n_1420),
.Y(n_1432)
);

NOR4xp25_ASAP7_75t_SL g1433 ( 
.A(n_1432),
.B(n_1302),
.C(n_1321),
.D(n_1417),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1425),
.B(n_1421),
.Y(n_1434)
);

OAI21xp33_ASAP7_75t_L g1435 ( 
.A1(n_1426),
.A2(n_1406),
.B(n_1419),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1428),
.A2(n_1410),
.B1(n_1419),
.B2(n_1345),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1424),
.A2(n_1331),
.B1(n_1419),
.B2(n_1325),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1429),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1431),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_1414),
.B2(n_1404),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1424),
.A2(n_1320),
.B(n_1275),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1427),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1430),
.Y(n_1443)
);

OAI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1436),
.A2(n_1388),
.B(n_1380),
.Y(n_1444)
);

AOI221x1_ASAP7_75t_L g1445 ( 
.A1(n_1435),
.A2(n_1324),
.B1(n_1338),
.B2(n_1162),
.C(n_1392),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1437),
.A2(n_1272),
.B(n_1237),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1437),
.A2(n_1391),
.B1(n_1387),
.B2(n_1302),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1443),
.B(n_1344),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1441),
.A2(n_1344),
.B(n_1279),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_SL g1450 ( 
.A(n_1442),
.B(n_1305),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1440),
.B(n_1391),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1438),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1434),
.B(n_1237),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1453),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1446),
.B(n_1433),
.C(n_1439),
.Y(n_1455)
);

OA22x2_ASAP7_75t_L g1456 ( 
.A1(n_1446),
.A2(n_1153),
.B1(n_1405),
.B2(n_1194),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1447),
.A2(n_1405),
.B1(n_1267),
.B2(n_1359),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1450),
.A2(n_1267),
.B(n_1153),
.Y(n_1458)
);

OAI211xp5_ASAP7_75t_L g1459 ( 
.A1(n_1445),
.A2(n_1251),
.B(n_1265),
.C(n_1282),
.Y(n_1459)
);

OA211x2_ASAP7_75t_L g1460 ( 
.A1(n_1444),
.A2(n_1315),
.B(n_1316),
.C(n_1290),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1451),
.B(n_1394),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1448),
.A2(n_1449),
.B(n_1452),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_R g1463 ( 
.A(n_1454),
.B(n_1321),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1456),
.B(n_1399),
.Y(n_1464)
);

AOI211xp5_ASAP7_75t_L g1465 ( 
.A1(n_1455),
.A2(n_1315),
.B(n_1265),
.C(n_1282),
.Y(n_1465)
);

AOI221x1_ASAP7_75t_L g1466 ( 
.A1(n_1458),
.A2(n_1167),
.B1(n_1143),
.B2(n_1158),
.C(n_1126),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1461),
.B(n_1462),
.Y(n_1467)
);

AOI21xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1457),
.A2(n_1283),
.B(n_1176),
.Y(n_1468)
);

NOR3xp33_ASAP7_75t_L g1469 ( 
.A(n_1459),
.B(n_1167),
.C(n_1158),
.Y(n_1469)
);

OAI211xp5_ASAP7_75t_L g1470 ( 
.A1(n_1460),
.A2(n_1251),
.B(n_1328),
.C(n_1294),
.Y(n_1470)
);

AOI211xp5_ASAP7_75t_L g1471 ( 
.A1(n_1455),
.A2(n_1326),
.B(n_1291),
.C(n_1308),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1467),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1471),
.A2(n_1356),
.B1(n_1359),
.B2(n_1366),
.Y(n_1473)
);

NOR2xp67_ASAP7_75t_L g1474 ( 
.A(n_1464),
.B(n_1359),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1463),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1466),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1468),
.Y(n_1477)
);

NOR2xp67_ASAP7_75t_SL g1478 ( 
.A(n_1472),
.B(n_1470),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1477),
.Y(n_1479)
);

NAND4xp75_ASAP7_75t_L g1480 ( 
.A(n_1476),
.B(n_1474),
.C(n_1475),
.D(n_1465),
.Y(n_1480)
);

NAND4xp25_ASAP7_75t_L g1481 ( 
.A(n_1473),
.B(n_1469),
.C(n_1174),
.D(n_1144),
.Y(n_1481)
);

NOR2xp67_ASAP7_75t_L g1482 ( 
.A(n_1479),
.B(n_1359),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1478),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1480),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1481),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1479),
.Y(n_1486)
);

XNOR2x2_ASAP7_75t_L g1487 ( 
.A(n_1483),
.B(n_1176),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1486),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1485),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1484),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1490),
.A2(n_1484),
.B1(n_1482),
.B2(n_1135),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1488),
.Y(n_1492)
);

AO22x2_ASAP7_75t_L g1493 ( 
.A1(n_1489),
.A2(n_1290),
.B1(n_1316),
.B2(n_1116),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1487),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1490),
.B(n_1290),
.Y(n_1495)
);

OAI22x1_ASAP7_75t_L g1496 ( 
.A1(n_1494),
.A2(n_1155),
.B1(n_1173),
.B2(n_1169),
.Y(n_1496)
);

XOR2xp5_ASAP7_75t_L g1497 ( 
.A(n_1495),
.B(n_1155),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1492),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1493),
.Y(n_1499)
);

OAI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1498),
.A2(n_1491),
.B1(n_1359),
.B2(n_1173),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1499),
.B(n_1334),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1496),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1502),
.B(n_1497),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1503),
.A2(n_1500),
.B1(n_1501),
.B2(n_1316),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1503),
.A2(n_1174),
.B1(n_1144),
.B2(n_1122),
.Y(n_1505)
);

OR2x6_ASAP7_75t_L g1506 ( 
.A(n_1504),
.B(n_1136),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1506),
.A2(n_1505),
.B1(n_1169),
.B2(n_1122),
.Y(n_1507)
);


endmodule