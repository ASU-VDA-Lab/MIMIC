module fake_ariane_2106_n_188 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_188);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_188;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_178;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVxp33_ASAP7_75t_SL g43 ( 
.A(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVxp67_ASAP7_75t_SL g49 ( 
.A(n_24),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_31),
.A2(n_1),
.B(n_3),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_33),
.B(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_8),
.B1(n_10),
.B2(n_14),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_33),
.B(n_8),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_46),
.B1(n_35),
.B2(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_48),
.B1(n_36),
.B2(n_34),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_42),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_34),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_71),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

OAI221xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_35),
.B1(n_51),
.B2(n_49),
.C(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_56),
.B(n_50),
.Y(n_88)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_15),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_69),
.B(n_64),
.C(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

NAND2x1p5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_60),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_64),
.B(n_60),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_91),
.Y(n_102)
);

O2A1O1Ixp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_79),
.B(n_78),
.C(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_82),
.Y(n_107)
);

NAND2x1p5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_99),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_93),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_105),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_109),
.A2(n_106),
.B(n_84),
.C(n_80),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_97),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_102),
.Y(n_115)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_100),
.B(n_92),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_100),
.B(n_92),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_110),
.B(n_80),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_115),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_87),
.C(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_75),
.B(n_102),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_96),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_126),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_77),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_131),
.Y(n_148)
);

AOI222xp33_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_75),
.B1(n_114),
.B2(n_63),
.C1(n_58),
.C2(n_59),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_122),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_127),
.B(n_114),
.C(n_70),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_143),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_122),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_61),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_149),
.B1(n_75),
.B2(n_114),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_122),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_125),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_154),
.B1(n_158),
.B2(n_131),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_128),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_82),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_128),
.Y(n_169)
);

NAND4xp75_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_60),
.C(n_76),
.D(n_86),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_113),
.B(n_112),
.C(n_114),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_61),
.Y(n_172)
);

NAND4xp75_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_86),
.C(n_76),
.D(n_116),
.Y(n_173)
);

NOR2x1p5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_111),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_166),
.A2(n_108),
.B(n_116),
.Y(n_175)
);

NOR2x1p5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_161),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_175),
.C(n_173),
.Y(n_177)
);

AOI31xp33_ASAP7_75t_SL g178 ( 
.A1(n_168),
.A2(n_160),
.A3(n_161),
.B(n_17),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_111),
.B(n_113),
.C(n_95),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_111),
.B1(n_116),
.B2(n_21),
.Y(n_180)
);

NOR2x1p5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_111),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_16),
.Y(n_183)
);

AOI211xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_177),
.B(n_182),
.C(n_179),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_108),
.B1(n_116),
.B2(n_95),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_184),
.B(n_185),
.C(n_95),
.Y(n_188)
);


endmodule