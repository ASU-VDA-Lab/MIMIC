module fake_jpeg_5150_n_88 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_0),
.Y(n_65)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_60),
.Y(n_66)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_41),
.B1(n_40),
.B2(n_45),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_47),
.B1(n_52),
.B2(n_51),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_44),
.B1(n_49),
.B2(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_1),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_69),
.B1(n_66),
.B2(n_43),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_54),
.B1(n_46),
.B2(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_4),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_67),
.B(n_6),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_3),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_75),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_13),
.C(n_14),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_15),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_81),
.A2(n_77),
.B1(n_18),
.B2(n_25),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_78),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g84 ( 
.A(n_83),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_16),
.C(n_26),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

O2A1O1Ixp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_27),
.B(n_28),
.C(n_30),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_31),
.Y(n_88)
);


endmodule