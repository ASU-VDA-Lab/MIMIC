module fake_jpeg_12281_n_471 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_471);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_471;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_65),
.Y(n_100)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_26),
.B(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_68),
.B(n_71),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx2_ASAP7_75t_SL g123 ( 
.A(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_15),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_15),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_87),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_35),
.Y(n_80)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_37),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_88),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_84),
.Y(n_99)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_86),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_29),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_49),
.Y(n_140)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_28),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_139),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_78),
.A2(n_60),
.B1(n_74),
.B2(n_70),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_115),
.A2(n_60),
.B1(n_74),
.B2(n_86),
.Y(n_166)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_61),
.A2(n_30),
.B1(n_25),
.B2(n_38),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_129),
.A2(n_43),
.B1(n_39),
.B2(n_19),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_77),
.A2(n_30),
.B1(n_48),
.B2(n_49),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_130),
.A2(n_44),
.B1(n_40),
.B2(n_48),
.Y(n_199)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_140),
.Y(n_171)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_53),
.Y(n_149)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_94),
.B(n_38),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_28),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_152),
.B(n_162),
.Y(n_238)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

BUFx24_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_154),
.Y(n_215)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_155),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_80),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_170),
.Y(n_208)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_157),
.Y(n_236)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_158),
.Y(n_244)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_159),
.Y(n_232)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_107),
.B(n_29),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_164),
.B(n_46),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_70),
.B1(n_65),
.B2(n_57),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_123),
.B1(n_115),
.B2(n_143),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_167),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_108),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_169),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_30),
.A3(n_56),
.B1(n_90),
.B2(n_95),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_82),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_98),
.B(n_32),
.C(n_31),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_178),
.Y(n_216)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_101),
.A2(n_83),
.B1(n_69),
.B2(n_64),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_185),
.B1(n_199),
.B2(n_147),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_175),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_31),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_189),
.Y(n_218)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_99),
.B(n_92),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_142),
.A2(n_39),
.B(n_34),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_188),
.Y(n_217)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g234 ( 
.A(n_181),
.Y(n_234)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_109),
.A2(n_63),
.B1(n_62),
.B2(n_36),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_20),
.C(n_32),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_102),
.B(n_34),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_43),
.B1(n_19),
.B2(n_20),
.Y(n_209)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_201),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_106),
.B(n_46),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_193),
.Y(n_222)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_196),
.Y(n_224)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_111),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_198),
.Y(n_225)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_180),
.B1(n_165),
.B2(n_190),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_203),
.A2(n_214),
.B1(n_229),
.B2(n_154),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_211),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_205),
.B(n_223),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_104),
.B1(n_121),
.B2(n_127),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_209),
.A2(n_246),
.B1(n_33),
.B2(n_3),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g286 ( 
.A(n_213),
.B(n_6),
.C(n_7),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_109),
.B1(n_137),
.B2(n_145),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_161),
.A2(n_127),
.B1(n_134),
.B2(n_145),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_220),
.A2(n_155),
.B1(n_163),
.B2(n_45),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_147),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_92),
.Y(n_228)
);

NAND2xp33_ASAP7_75t_SL g269 ( 
.A(n_228),
.B(n_215),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_165),
.A2(n_132),
.B1(n_36),
.B2(n_44),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_156),
.A2(n_166),
.B1(n_184),
.B2(n_177),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_154),
.B(n_157),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_183),
.B(n_100),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_15),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_202),
.A2(n_132),
.B1(n_181),
.B2(n_195),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_187),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_267),
.C(n_279),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_179),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_249),
.B(n_271),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_237),
.A2(n_191),
.B1(n_182),
.B2(n_158),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_250),
.A2(n_261),
.B(n_265),
.Y(n_297)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_252),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_255),
.B1(n_263),
.B2(n_280),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_210),
.A2(n_44),
.B1(n_40),
.B2(n_48),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_257),
.A2(n_277),
.B1(n_215),
.B2(n_228),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_258),
.B(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_217),
.A2(n_87),
.B(n_48),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_262),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_45),
.B1(n_44),
.B2(n_41),
.Y(n_263)
);

NOR3xp33_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_45),
.C(n_41),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_264),
.B(n_272),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_217),
.A2(n_45),
.B1(n_41),
.B2(n_40),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_41),
.C(n_40),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_275),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_269),
.A2(n_270),
.B(n_206),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_230),
.A2(n_1),
.B(n_2),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_238),
.B(n_13),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_218),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_226),
.B(n_13),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_213),
.B(n_12),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_216),
.B(n_1),
.C(n_3),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_211),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_240),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_283),
.Y(n_317)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_245),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_216),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_284),
.A2(n_229),
.B1(n_277),
.B2(n_214),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_225),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_285),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_286),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_208),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_289),
.B(n_295),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_290),
.A2(n_301),
.B1(n_284),
.B2(n_234),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_274),
.B(n_208),
.CI(n_216),
.CON(n_291),
.SN(n_291)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_280),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_208),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_310),
.C(n_315),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_267),
.B(n_222),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_298),
.A2(n_308),
.B1(n_311),
.B2(n_253),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_270),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_256),
.A2(n_209),
.B1(n_204),
.B2(n_246),
.Y(n_301)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_256),
.A2(n_204),
.B1(n_233),
.B2(n_234),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_228),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_256),
.A2(n_204),
.B1(n_234),
.B2(n_241),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_227),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_251),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_318),
.B(n_252),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_279),
.B(n_227),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_294),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_241),
.C(n_242),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_243),
.C(n_245),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_253),
.A2(n_243),
.B(n_244),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_247),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_323),
.A2(n_338),
.B1(n_343),
.B2(n_352),
.Y(n_359)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_324),
.Y(n_354)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_326),
.Y(n_363)
);

AOI21xp33_ASAP7_75t_L g358 ( 
.A1(n_327),
.A2(n_330),
.B(n_350),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_314),
.A2(n_250),
.B(n_265),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_328),
.A2(n_333),
.B(n_342),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_329),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_263),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_331),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_341),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_314),
.A2(n_283),
.B(n_281),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_334),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_207),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_335),
.B(n_344),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_302),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_276),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_346),
.C(n_310),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_311),
.A2(n_266),
.B1(n_262),
.B2(n_259),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_317),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_299),
.A2(n_273),
.B(n_207),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_308),
.A2(n_298),
.B1(n_322),
.B2(n_304),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_306),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_288),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_347),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_303),
.Y(n_348)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_348),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_297),
.A2(n_231),
.B(n_221),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_349),
.B(n_322),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_291),
.A2(n_221),
.B(n_244),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_305),
.Y(n_351)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_351),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_309),
.B(n_231),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_373),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_357),
.B(n_337),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_295),
.C(n_302),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_375),
.C(n_345),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_365),
.A2(n_331),
.B(n_307),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_292),
.Y(n_367)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_343),
.A2(n_301),
.B1(n_287),
.B2(n_291),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_368),
.A2(n_212),
.B1(n_236),
.B2(n_219),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_292),
.Y(n_369)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_315),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_323),
.A2(n_287),
.B1(n_293),
.B2(n_312),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_374),
.A2(n_378),
.B1(n_329),
.B2(n_331),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_319),
.C(n_321),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_316),
.Y(n_377)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_377),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_338),
.A2(n_324),
.B1(n_328),
.B2(n_349),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_296),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_327),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_395),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_388),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_353),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_386),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_350),
.C(n_346),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_390),
.C(n_397),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_361),
.Y(n_384)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

NAND3xp33_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_351),
.C(n_333),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_377),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_391),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_360),
.B(n_327),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_342),
.C(n_334),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_326),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_399),
.B1(n_370),
.B2(n_363),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_236),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_393),
.B(n_364),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_368),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_307),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_396),
.A2(n_365),
.B(n_371),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_320),
.C(n_219),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_376),
.A2(n_354),
.B1(n_371),
.B2(n_372),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_400),
.A2(n_376),
.B1(n_361),
.B2(n_354),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_403),
.A2(n_408),
.B1(n_399),
.B2(n_401),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_355),
.C(n_356),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_404),
.B(n_411),
.Y(n_429)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_400),
.A2(n_398),
.B1(n_372),
.B2(n_401),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_356),
.C(n_359),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_417),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_414),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_379),
.C(n_370),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_415),
.B(n_416),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_363),
.C(n_358),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_383),
.B(n_362),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_388),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_6),
.Y(n_431)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_380),
.C(n_397),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_421),
.B(n_423),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_396),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_391),
.C(n_385),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_424),
.B(n_426),
.C(n_431),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_402),
.B(n_385),
.C(n_395),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g427 ( 
.A(n_411),
.B(n_384),
.CI(n_362),
.CON(n_427),
.SN(n_427)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_428),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_406),
.A2(n_384),
.B(n_212),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_404),
.B(n_7),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g444 ( 
.A(n_432),
.Y(n_444)
);

OAI321xp33_ASAP7_75t_L g434 ( 
.A1(n_433),
.A2(n_419),
.A3(n_409),
.B1(n_416),
.B2(n_413),
.C(n_415),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_434),
.B(n_438),
.Y(n_446)
);

OAI21x1_ASAP7_75t_SL g435 ( 
.A1(n_425),
.A2(n_418),
.B(n_402),
.Y(n_435)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_435),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_424),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_443),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_410),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_422),
.A2(n_410),
.B(n_8),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_442),
.A2(n_431),
.B(n_423),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_429),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_422),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_7),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_448),
.B(n_442),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_421),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_SL g455 ( 
.A(n_449),
.B(n_446),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_439),
.B(n_430),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_453),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_438),
.A2(n_427),
.B(n_430),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_452),
.A2(n_446),
.B(n_437),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_427),
.C(n_9),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_10),
.Y(n_460)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_455),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_437),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_457),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_458),
.A2(n_450),
.B(n_445),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_460),
.B(n_444),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_461),
.B(n_464),
.Y(n_465)
);

AOI21xp33_ASAP7_75t_L g466 ( 
.A1(n_463),
.A2(n_459),
.B(n_456),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_441),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_467),
.A2(n_465),
.B(n_462),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_441),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_10),
.B1(n_11),
.B2(n_443),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_470),
.B(n_10),
.Y(n_471)
);


endmodule