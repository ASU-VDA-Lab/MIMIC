module real_jpeg_17168_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_0),
.A2(n_108),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_0),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_0),
.A2(n_295),
.B1(n_408),
.B2(n_411),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_0),
.A2(n_295),
.B1(n_467),
.B2(n_472),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_1),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_1),
.Y(n_127)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_1),
.Y(n_204)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_3),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_3),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_116),
.B1(n_133),
.B2(n_137),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_3),
.A2(n_116),
.B1(n_208),
.B2(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_3),
.A2(n_116),
.B1(n_387),
.B2(n_390),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_4),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_4),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_4),
.A2(n_320),
.B1(n_422),
.B2(n_424),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_5),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_5),
.A2(n_78),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_5),
.A2(n_78),
.B1(n_218),
.B2(n_222),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_5),
.A2(n_78),
.B1(n_359),
.B2(n_361),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_6),
.Y(n_95)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_6),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_6),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_7),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_7),
.Y(n_239)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_7),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_7),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_8),
.A2(n_253),
.B1(n_257),
.B2(n_258),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_8),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_8),
.A2(n_188),
.B1(n_257),
.B2(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_8),
.A2(n_257),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_9),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_9),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_9),
.A2(n_86),
.B1(n_183),
.B2(n_187),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_9),
.A2(n_86),
.B1(n_366),
.B2(n_369),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_9),
.A2(n_86),
.B1(n_357),
.B2(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_10),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_10),
.Y(n_355)
);

BUFx8_ASAP7_75t_L g389 ( 
.A(n_10),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_11),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_11),
.A2(n_106),
.B1(n_117),
.B2(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_11),
.A2(n_106),
.B1(n_215),
.B2(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_11),
.A2(n_106),
.B1(n_479),
.B2(n_481),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_12),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_12),
.Y(n_340)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_12),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_13),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_13),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_14),
.Y(n_90)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_15),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_15),
.B(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_15),
.B(n_74),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_15),
.A2(n_39),
.B1(n_208),
.B2(n_212),
.Y(n_207)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_15),
.A2(n_227),
.A3(n_231),
.B1(n_235),
.B2(n_240),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_15),
.B(n_283),
.Y(n_282)
);

OAI32xp33_ASAP7_75t_L g321 ( 
.A1(n_15),
.A2(n_322),
.A3(n_326),
.B1(n_331),
.B2(n_334),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_15),
.A2(n_39),
.B1(n_353),
.B2(n_356),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_451),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_376),
.B(n_448),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_304),
.B(n_375),
.Y(n_19)
);

AOI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_263),
.B(n_303),
.Y(n_20)
);

OAI21x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_175),
.B(n_262),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_128),
.B(n_174),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_82),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_24),
.B(n_82),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_48),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_25),
.A2(n_48),
.B1(n_49),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_25),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.A3(n_34),
.B1(n_38),
.B2(n_42),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AO22x2_ASAP7_75t_L g123 ( 
.A1(n_28),
.A2(n_77),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_32),
.Y(n_140)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_39),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_39),
.A2(n_91),
.B1(n_153),
.B2(n_156),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_39),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_39),
.B(n_332),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_41),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_41),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_55),
.B1(n_74),
.B2(n_75),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_55),
.A2(n_74),
.B1(n_75),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_55),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_55),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_55),
.B(n_373),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_67),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_59),
.B1(n_62),
.B2(n_66),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g179 ( 
.A1(n_67),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_67),
.B(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_67),
.A2(n_180),
.B1(n_420),
.B2(n_421),
.Y(n_419)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_68),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_72),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_74),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_74),
.B(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_81),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_81),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_110),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_83),
.B(n_111),
.C(n_122),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_91),
.B(n_96),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_89),
.Y(n_294)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_89),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_90),
.Y(n_261)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_91),
.A2(n_132),
.B1(n_156),
.B2(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_91),
.B(n_252),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_91),
.A2(n_103),
.B(n_144),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_94),
.A2(n_292),
.B(n_296),
.Y(n_291)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_97),
.B(n_296),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_100),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_103),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_122),
.Y(n_110)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_121),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_123),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_123),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_123),
.B(n_439),
.Y(n_438)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_150),
.B(n_173),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_148),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_130),
.B(n_148),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_141),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_141),
.A2(n_292),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_141),
.A2(n_248),
.B(n_316),
.Y(n_404)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_167),
.B(n_172),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_163),
.Y(n_151)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_171),
.Y(n_172)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_176),
.B(n_177),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_225),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_190),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_179),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_180),
.A2(n_273),
.B(n_372),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g460 ( 
.A1(n_180),
.A2(n_372),
.B(n_421),
.Y(n_460)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_182),
.Y(n_271)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_185),
.Y(n_374)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_190),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_207),
.B1(n_217),
.B2(n_224),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_191),
.A2(n_217),
.B1(n_224),
.B2(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_191),
.A2(n_224),
.B1(n_298),
.B2(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_191),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_191),
.A2(n_396),
.B(n_438),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_191),
.A2(n_224),
.B1(n_465),
.B2(n_466),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B1(n_200),
.B2(n_205),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_197),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_199),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_199),
.Y(n_471)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_206),
.Y(n_440)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_211),
.Y(n_333)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

AO22x2_ASAP7_75t_L g283 ( 
.A1(n_220),
.A2(n_284),
.B1(n_286),
.B2(n_289),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_221),
.Y(n_400)
);

INVx3_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_SL g395 ( 
.A(n_224),
.B(n_396),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_265),
.C(n_266),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_246),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_246),
.Y(n_269)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_230),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_230),
.Y(n_442)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_259),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_264),
.B(n_267),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_278),
.B1(n_279),
.B2(n_302),
.Y(n_267)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

XOR2x1_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_270),
.C(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_297),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_290),
.B2(n_291),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_297),
.C(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OR2x6_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_283),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_283),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_283),
.B(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_285),
.Y(n_370)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_288),
.Y(n_289)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_305),
.B(n_306),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_341),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_309),
.B(n_311),
.C(n_341),
.Y(n_445)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_321),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_313),
.B(n_321),
.Y(n_401)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_329),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_329),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_330),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_363),
.Y(n_341)
);

MAJx2_ASAP7_75t_L g402 ( 
.A(n_342),
.B(n_364),
.C(n_371),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_352),
.B1(n_358),
.B2(n_362),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_343),
.Y(n_384)
);

OAI22x1_ASAP7_75t_SL g432 ( 
.A1(n_343),
.A2(n_362),
.B1(n_386),
.B2(n_433),
.Y(n_432)
);

OAI21x1_ASAP7_75t_SL g476 ( 
.A1(n_343),
.A2(n_433),
.B(n_477),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_348),
.B2(n_349),
.Y(n_344)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_346),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_346),
.Y(n_360)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx12f_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_355),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_355),
.Y(n_436)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_371),
.Y(n_363)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_365),
.Y(n_394)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_444),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_414),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_379),
.B(n_414),
.C(n_450),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_402),
.C(n_403),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_380),
.B(n_447),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_401),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_392),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_392),
.C(n_401),
.Y(n_415)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx12f_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_389),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_394),
.B(n_395),
.Y(n_392)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_402),
.B(n_403),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_405),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_413),
.Y(n_405)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_407),
.Y(n_420)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_428),
.C(n_443),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_428),
.B1(n_429),
.B2(n_443),
.Y(n_416)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_418),
.B(n_419),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_430),
.B(n_432),
.C(n_437),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_437),
.Y(n_431)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_445),
.B(n_446),
.Y(n_450)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_486),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_455),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_456),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_455)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_456),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_462),
.Y(n_456)
);

OAI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_460),
.B2(n_461),
.Y(n_457)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_458),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XNOR2x1_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_482),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_476),
.Y(n_463)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_471),
.Y(n_475)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);


endmodule