module fake_jpeg_23845_n_318 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_22),
.B1(n_16),
.B2(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_33),
.B1(n_37),
.B2(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_33),
.B1(n_37),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_25),
.B1(n_19),
.B2(n_27),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_19),
.B1(n_27),
.B2(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_65),
.B(n_79),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_27),
.B1(n_25),
.B2(n_31),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_32),
.B1(n_22),
.B2(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_77),
.Y(n_99)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_23),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_29),
.B(n_38),
.C(n_34),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_31),
.B1(n_32),
.B2(n_44),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_81),
.A2(n_91),
.B1(n_75),
.B2(n_68),
.Y(n_121)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_39),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_94),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_34),
.C(n_38),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_96),
.C(n_98),
.Y(n_106)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_36),
.A3(n_38),
.B1(n_34),
.B2(n_55),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_92),
.B(n_96),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_15),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_38),
.C(n_36),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_98),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_74),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_106),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_108),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_101),
.A2(n_38),
.B(n_55),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_109),
.Y(n_138)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_78),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_76),
.C(n_72),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_95),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_116),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_22),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_56),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_69),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_45),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_119),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_20),
.B(n_15),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_89),
.B(n_94),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_46),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_41),
.B1(n_75),
.B2(n_47),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_72),
.B1(n_95),
.B2(n_62),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_56),
.B1(n_47),
.B2(n_91),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_102),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_126),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_130),
.B(n_143),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_132),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_116),
.B(n_113),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_133),
.B1(n_97),
.B2(n_59),
.Y(n_157)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

OAI22x1_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_18),
.B1(n_22),
.B2(n_58),
.Y(n_133)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_102),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_147),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_124),
.B1(n_111),
.B2(n_119),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_103),
.B(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_148),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_112),
.C(n_114),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_82),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_103),
.B(n_45),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_152),
.Y(n_177)
);

AO21x2_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_80),
.B(n_62),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_59),
.B1(n_74),
.B2(n_73),
.Y(n_165)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_153),
.A2(n_46),
.B1(n_57),
.B2(n_53),
.Y(n_203)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_174),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_157),
.A2(n_164),
.B1(n_19),
.B2(n_14),
.Y(n_204)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_109),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_158),
.A2(n_160),
.B(n_165),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_104),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_173),
.C(n_144),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_106),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_176),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_106),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_171),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_151),
.A2(n_109),
.B1(n_107),
.B2(n_124),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_114),
.B(n_112),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_178),
.B(n_148),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_115),
.C(n_125),
.Y(n_173)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_100),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_15),
.B(n_26),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_128),
.B(n_150),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_90),
.B(n_85),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_28),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_28),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_180),
.A2(n_187),
.B(n_20),
.Y(n_219)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_189),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_73),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_144),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_195),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_192),
.C(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_149),
.C(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_129),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_160),
.B(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_166),
.A2(n_151),
.B1(n_127),
.B2(n_135),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_198),
.A2(n_169),
.B1(n_175),
.B2(n_24),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_151),
.C(n_57),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_200),
.B(n_26),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_151),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_202),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_164),
.B1(n_170),
.B2(n_165),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_153),
.B1(n_165),
.B2(n_166),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_53),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_160),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_207),
.A2(n_218),
.B1(n_204),
.B2(n_198),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_210),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_158),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_169),
.B1(n_174),
.B2(n_165),
.Y(n_213)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_195),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_219),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_225),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_181),
.A2(n_73),
.B1(n_50),
.B2(n_14),
.Y(n_226)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_26),
.C(n_24),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_24),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_205),
.C(n_191),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_184),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_191),
.C(n_196),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_233),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_208),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_196),
.C(n_192),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_242),
.B(n_244),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_199),
.C(n_203),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_17),
.B1(n_23),
.B2(n_13),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_50),
.C(n_17),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_245),
.A2(n_223),
.B1(n_211),
.B2(n_219),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_248),
.B(n_241),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_213),
.B(n_206),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_265),
.C(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

A2O1A1O1Ixp25_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_210),
.B(n_216),
.C(n_209),
.D(n_218),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_251),
.B(n_253),
.Y(n_270)
);

A2O1A1O1Ixp25_ASAP7_75t_L g253 ( 
.A1(n_246),
.A2(n_226),
.B(n_13),
.C(n_12),
.D(n_14),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_13),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_260),
.Y(n_275)
);

AO22x1_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_259)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_17),
.B(n_1),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_238),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_12),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_259),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_274),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_228),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_267),
.B(n_249),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_241),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_269),
.B1(n_254),
.B2(n_252),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_247),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_279),
.B(n_280),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_229),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_0),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_286),
.C(n_287),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_253),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_283),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_275),
.B(n_279),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_289),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_255),
.B1(n_260),
.B2(n_262),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_265),
.C(n_251),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_261),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_270),
.A2(n_12),
.B(n_3),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_293),
.C(n_8),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_0),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_291),
.B(n_292),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_272),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_11),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_295),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_288),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_299),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_6),
.B(n_7),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_303),
.B(n_300),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_293),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_8),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_11),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_309),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_301),
.B1(n_296),
.B2(n_10),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_308),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_8),
.B(n_9),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_304),
.Y(n_313)
);

AO21x1_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_311),
.B(n_306),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_310),
.C(n_10),
.Y(n_316)
);

OAI221xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.C(n_266),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_9),
.Y(n_318)
);


endmodule