module fake_jpeg_29865_n_188 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_44),
.Y(n_49)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_1),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_2),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_17),
.B1(n_31),
.B2(n_29),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_53),
.B1(n_61),
.B2(n_63),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_17),
.C(n_27),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_51),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_3),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_59),
.B1(n_67),
.B2(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_27),
.B1(n_25),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_25),
.B1(n_30),
.B2(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_40),
.Y(n_71)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_35),
.A2(n_23),
.B1(n_25),
.B2(n_22),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_84),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_76),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_65),
.B1(n_51),
.B2(n_69),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_41),
.B1(n_35),
.B2(n_39),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_87),
.B1(n_62),
.B2(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_39),
.B(n_22),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_20),
.C(n_52),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_88),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_36),
.B1(n_16),
.B2(n_39),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_16),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_20),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_13),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_110)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_54),
.B(n_39),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_66),
.A3(n_64),
.B1(n_62),
.B2(n_39),
.Y(n_98)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

AOI221xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_100),
.B1(n_94),
.B2(n_76),
.C(n_79),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_99),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_115),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_77),
.B1(n_83),
.B2(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_113),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_75),
.B1(n_87),
.B2(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_126),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_122),
.B1(n_125),
.B2(n_102),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_124),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_85),
.B1(n_93),
.B2(n_73),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_71),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_107),
.A2(n_76),
.B1(n_92),
.B2(n_60),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_107),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_128),
.B(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_92),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_131),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_76),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_130),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_95),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_101),
.B(n_114),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_103),
.B(n_20),
.C(n_10),
.D(n_11),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_137),
.B1(n_146),
.B2(n_123),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_106),
.B1(n_111),
.B2(n_113),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_144),
.C(n_145),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_103),
.B(n_105),
.C(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_148),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_60),
.C(n_56),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_78),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_57),
.B1(n_8),
.B2(n_9),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_117),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_145),
.B1(n_146),
.B2(n_134),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_133),
.C(n_119),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_156),
.C(n_142),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_118),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_116),
.C(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_129),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_166),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_150),
.A2(n_135),
.B1(n_147),
.B2(n_144),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_157),
.B1(n_154),
.B2(n_9),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_165),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_168),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_136),
.C(n_57),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_20),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_156),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_166),
.B(n_163),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_173),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_157),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_174),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_169),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_165),
.B(n_164),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_177),
.A2(n_179),
.B(n_6),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_11),
.B(n_13),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_183),
.C(n_57),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_181),
.B(n_182),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_171),
.B(n_8),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_184),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_6),
.Y(n_188)
);


endmodule