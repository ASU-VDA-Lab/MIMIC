module fake_netlist_5_1368_n_1774 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1774);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1774;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_60),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_1),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_59),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_113),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_24),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_24),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_47),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_22),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_13),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_50),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_148),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_105),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_73),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_54),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_61),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_74),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_94),
.Y(n_190)
);

BUFx8_ASAP7_75t_SL g191 ( 
.A(n_96),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_26),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_70),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_43),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_84),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_30),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_25),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_68),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_85),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_17),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_23),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_92),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_18),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_102),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_121),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_2),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_57),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_7),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_20),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_72),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_132),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_86),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_29),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_123),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_65),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_64),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_97),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_2),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_89),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_93),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_137),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_48),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_112),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_101),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_62),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_22),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_116),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_131),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_47),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_15),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_35),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_98),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_38),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_51),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_151),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_12),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_45),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_26),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_25),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_8),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_150),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_39),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_18),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_31),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_136),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_39),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_49),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_28),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_1),
.Y(n_257)
);

BUFx2_ASAP7_75t_SL g258 ( 
.A(n_21),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_67),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_56),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_13),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_33),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_10),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_54),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_63),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_134),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_42),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_79),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_122),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_77),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_48),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_56),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_46),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_147),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_125),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_146),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_109),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_29),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_129),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_152),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_155),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_59),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_9),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_42),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_52),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_21),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_117),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_44),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_51),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_138),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_11),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_35),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_6),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_49),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_111),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_45),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_75),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_41),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_57),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_8),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_80),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_36),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_53),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_52),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_78),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_33),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_142),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_55),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_66),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_128),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_55),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_69),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_32),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_3),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_46),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_28),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_225),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_160),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_164),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_184),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_196),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_166),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_184),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_188),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_184),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_184),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_196),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_0),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_195),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_201),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_190),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_198),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_195),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_193),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_199),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_R g337 ( 
.A(n_174),
.B(n_0),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_195),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_241),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_197),
.B(n_3),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_206),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_201),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_241),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_205),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_232),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_192),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_212),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_195),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_203),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_203),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_281),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_203),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_203),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_208),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_308),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_260),
.B(n_4),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_212),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_304),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_300),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_300),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_308),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_204),
.B(n_5),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_204),
.B(n_224),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_281),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_291),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_268),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_291),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_168),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_224),
.B(n_187),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_170),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_165),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_215),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_310),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_216),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_310),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_191),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_316),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_218),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_213),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_223),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_219),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_191),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_226),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_228),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_243),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_247),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_261),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_214),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_192),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_371),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_343),
.B(n_187),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_321),
.B(n_279),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_371),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_321),
.B(n_279),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_324),
.B(n_298),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_371),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_371),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_343),
.B(n_163),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_326),
.B(n_167),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_360),
.Y(n_408)
);

CKINVDCx11_ASAP7_75t_R g409 ( 
.A(n_380),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_326),
.B(n_182),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_169),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_360),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_327),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_327),
.B(n_330),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_334),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_334),
.Y(n_417)
);

NAND2xp33_ASAP7_75t_SL g418 ( 
.A(n_337),
.B(n_202),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_338),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_338),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_348),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_348),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_349),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_349),
.Y(n_424)
);

BUFx8_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_350),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_345),
.B(n_359),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_372),
.B(n_207),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_346),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_352),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_351),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_352),
.B(n_353),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_353),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_354),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_354),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_339),
.B(n_174),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_356),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_356),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_358),
.B(n_189),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_362),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_362),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_367),
.B(n_177),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_363),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_368),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_373),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_373),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_345),
.B(n_192),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_374),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_368),
.B(n_194),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_344),
.B(n_257),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_329),
.B(n_217),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_383),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_365),
.B(n_200),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_322),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_418),
.Y(n_467)
);

BUFx6f_ASAP7_75t_SL g468 ( 
.A(n_449),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_413),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_418),
.A2(n_340),
.B1(n_202),
.B2(n_288),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_396),
.B(n_370),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_414),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_414),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_411),
.B(n_319),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_320),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_432),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_414),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_411),
.B(n_375),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_323),
.Y(n_479)
);

AND3x4_ASAP7_75t_L g480 ( 
.A(n_449),
.B(n_333),
.C(n_307),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_413),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_414),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_413),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_409),
.Y(n_484)
);

BUFx10_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_413),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_429),
.B(n_325),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_417),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_437),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_417),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_395),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_396),
.B(n_370),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_318),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_449),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_461),
.B(n_375),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_409),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_463),
.B(n_332),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_417),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_437),
.B(n_335),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_465),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_449),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_465),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_396),
.B(n_369),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_446),
.B(n_336),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_395),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_425),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_417),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_446),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_420),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_460),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_463),
.B(n_341),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_452),
.B(n_355),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_452),
.B(n_376),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_425),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_403),
.B(n_384),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_403),
.B(n_378),
.Y(n_520)
);

OR2x6_ASAP7_75t_L g521 ( 
.A(n_427),
.B(n_258),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_405),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_427),
.A2(n_392),
.B1(n_388),
.B2(n_387),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_430),
.A2(n_307),
.B1(n_288),
.B2(n_256),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_404),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_430),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_430),
.B(n_382),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_395),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_L g531 ( 
.A(n_403),
.B(n_385),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_425),
.B(n_177),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_420),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_425),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_403),
.B(n_168),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_460),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_425),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_395),
.Y(n_540)
);

BUFx8_ASAP7_75t_SL g541 ( 
.A(n_465),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_415),
.Y(n_542)
);

BUFx6f_ASAP7_75t_SL g543 ( 
.A(n_451),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_404),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_459),
.B(n_328),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_424),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_425),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_424),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_404),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_459),
.B(n_178),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_458),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_400),
.B(n_217),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_395),
.Y(n_553)
);

OAI22xp33_ASAP7_75t_L g554 ( 
.A1(n_400),
.A2(n_254),
.B1(n_229),
.B2(n_211),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_395),
.Y(n_555)
);

INVx5_ASAP7_75t_L g556 ( 
.A(n_404),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_400),
.B(n_178),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_416),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_416),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_416),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_458),
.B(n_389),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_419),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_419),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_419),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_458),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_421),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_404),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_424),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_458),
.B(n_220),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_424),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_445),
.B(n_391),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_445),
.B(n_391),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_421),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_464),
.B(n_180),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_464),
.A2(n_252),
.B1(n_299),
.B2(n_305),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_404),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_421),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_422),
.B(n_248),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_464),
.A2(n_299),
.B1(n_252),
.B2(n_309),
.Y(n_579)
);

AO22x2_ASAP7_75t_L g580 ( 
.A1(n_397),
.A2(n_262),
.B1(n_303),
.B2(n_301),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_464),
.A2(n_297),
.B1(n_289),
.B2(n_278),
.Y(n_581)
);

INVxp33_ASAP7_75t_SL g582 ( 
.A(n_406),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_395),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_395),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_406),
.B(n_389),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_426),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_404),
.B(n_168),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_422),
.B(n_253),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_464),
.A2(n_282),
.B1(n_295),
.B2(n_293),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_464),
.A2(n_267),
.B1(n_272),
.B2(n_186),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_426),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_422),
.B(n_265),
.Y(n_592)
);

NOR3xp33_ASAP7_75t_L g593 ( 
.A(n_406),
.B(n_227),
.C(n_210),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_410),
.B(n_168),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_L g595 ( 
.A(n_410),
.B(n_179),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_L g596 ( 
.A(n_410),
.B(n_179),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_401),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_422),
.B(n_266),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_407),
.B(n_276),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_426),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_401),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_441),
.B(n_390),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_407),
.B(n_412),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_428),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_428),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_441),
.B(n_179),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_445),
.B(n_390),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_407),
.B(n_412),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_407),
.B(n_277),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_451),
.B(n_222),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_451),
.B(n_230),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_454),
.B(n_180),
.Y(n_612)
);

AND3x1_ASAP7_75t_L g613 ( 
.A(n_454),
.B(n_457),
.C(n_455),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_401),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_401),
.Y(n_615)
);

NOR2xp67_ASAP7_75t_SL g616 ( 
.A(n_509),
.B(n_179),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_500),
.B(n_404),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_492),
.B(n_186),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_492),
.B(n_404),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_467),
.B(n_231),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_466),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_511),
.B(n_582),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_516),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_565),
.B(n_462),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_487),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_537),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_549),
.A2(n_399),
.B(n_397),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_511),
.B(n_485),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_537),
.B(n_173),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_514),
.B(n_408),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_466),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_472),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_504),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_479),
.B(n_408),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_565),
.B(n_408),
.Y(n_635)
);

INVxp33_ASAP7_75t_L g636 ( 
.A(n_541),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_474),
.B(n_489),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_504),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_569),
.A2(n_472),
.B1(n_477),
.B2(n_473),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_473),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_497),
.B(n_408),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_485),
.B(n_186),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_485),
.B(n_186),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_477),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_471),
.B(n_454),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_485),
.B(n_331),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_551),
.B(n_482),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_497),
.B(n_408),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_471),
.B(n_455),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_482),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_488),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_490),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_551),
.B(n_234),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_SL g654 ( 
.A1(n_524),
.A2(n_377),
.B1(n_342),
.B2(n_357),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_478),
.B(n_364),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_488),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_475),
.A2(n_379),
.B1(n_311),
.B2(n_306),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_571),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_522),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_571),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_467),
.A2(n_296),
.B1(n_287),
.B2(n_185),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_572),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_613),
.B(n_234),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_521),
.A2(n_181),
.B1(n_183),
.B2(n_185),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_490),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_572),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_607),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_521),
.A2(n_181),
.B1(n_183),
.B2(n_280),
.Y(n_668)
);

NOR3xp33_ASAP7_75t_L g669 ( 
.A(n_545),
.B(n_457),
.C(n_455),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_506),
.B(n_408),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_607),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_522),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_495),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_506),
.B(n_408),
.Y(n_674)
);

OAI22xp33_ASAP7_75t_L g675 ( 
.A1(n_521),
.A2(n_238),
.B1(n_233),
.B2(n_242),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_498),
.B(n_386),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_521),
.A2(n_613),
.B1(n_496),
.B2(n_507),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_476),
.Y(n_678)
);

BUFx12f_ASAP7_75t_SL g679 ( 
.A(n_521),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_496),
.B(n_561),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_487),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_561),
.B(n_408),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_495),
.B(n_408),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_569),
.B(n_407),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_569),
.B(n_407),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_527),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_527),
.Y(n_687)
);

OR2x6_ASAP7_75t_L g688 ( 
.A(n_552),
.B(n_259),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_538),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_538),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_519),
.B(n_457),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_502),
.A2(n_269),
.B1(n_290),
.B2(n_275),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_542),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_542),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_558),
.Y(n_695)
);

AOI221xp5_ASAP7_75t_L g696 ( 
.A1(n_554),
.A2(n_175),
.B1(n_176),
.B2(n_312),
.C(n_314),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_558),
.Y(n_697)
);

O2A1O1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_585),
.A2(n_441),
.B(n_397),
.C(n_399),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_503),
.B(n_312),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_476),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_519),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_585),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_520),
.B(n_161),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_529),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_569),
.B(n_412),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_552),
.A2(n_274),
.B1(n_212),
.B2(n_302),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_559),
.B(n_412),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_529),
.B(n_162),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_559),
.B(n_412),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_523),
.B(n_171),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_560),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_560),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_552),
.A2(n_212),
.B1(n_221),
.B2(n_270),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_562),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_562),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_563),
.Y(n_716)
);

INVxp33_ASAP7_75t_L g717 ( 
.A(n_480),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_563),
.B(n_564),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_602),
.B(n_234),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_SL g720 ( 
.A(n_547),
.B(n_257),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_564),
.B(n_412),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_552),
.A2(n_302),
.B1(n_221),
.B2(n_270),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_566),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_566),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_552),
.A2(n_302),
.B1(n_221),
.B2(n_270),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_573),
.B(n_428),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_487),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_573),
.B(n_577),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_577),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_586),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_599),
.A2(n_399),
.B(n_433),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_586),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_550),
.B(n_462),
.C(n_285),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_591),
.B(n_438),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_591),
.B(n_438),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_600),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_600),
.B(n_438),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_604),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_604),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_605),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_605),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_602),
.B(n_440),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_513),
.Y(n_743)
);

CKINVDCx6p67_ASAP7_75t_R g744 ( 
.A(n_543),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_610),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_487),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_469),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_578),
.B(n_440),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_531),
.A2(n_462),
.B1(n_456),
.B2(n_453),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_593),
.B(n_234),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_515),
.B(n_172),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_547),
.B(n_212),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_588),
.B(n_440),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_610),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_517),
.B(n_209),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_513),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_611),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_611),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_469),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_557),
.A2(n_456),
.B(n_453),
.C(n_450),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_470),
.B(n_286),
.C(n_235),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_513),
.B(n_236),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_592),
.B(n_436),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_481),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_598),
.B(n_436),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_481),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_609),
.B(n_212),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_580),
.A2(n_212),
.B1(n_221),
.B2(n_270),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_513),
.B(n_543),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_483),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_508),
.B(n_436),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_543),
.B(n_237),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_508),
.B(n_436),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_483),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_590),
.A2(n_456),
.B1(n_453),
.B2(n_450),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_580),
.B(n_470),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_580),
.A2(n_302),
.B1(n_270),
.B2(n_221),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_484),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_505),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_486),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_580),
.A2(n_302),
.B1(n_270),
.B2(n_221),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_505),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_508),
.B(n_530),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_486),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_637),
.B(n_509),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_633),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_702),
.A2(n_574),
.B(n_612),
.C(n_532),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_701),
.B(n_518),
.Y(n_788)
);

BUFx8_ASAP7_75t_L g789 ( 
.A(n_756),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_670),
.A2(n_576),
.B(n_525),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_633),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_674),
.A2(n_576),
.B(n_525),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_617),
.A2(n_576),
.B(n_525),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_702),
.B(n_494),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_680),
.B(n_494),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_623),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_715),
.B(n_494),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_715),
.B(n_758),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_634),
.A2(n_576),
.B(n_525),
.Y(n_799)
);

OAI321xp33_ASAP7_75t_L g800 ( 
.A1(n_710),
.A2(n_526),
.A3(n_524),
.B1(n_579),
.B2(n_575),
.C(n_589),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_758),
.B(n_494),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_701),
.B(n_540),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_677),
.A2(n_480),
.B1(n_468),
.B2(n_536),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_633),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_622),
.B(n_518),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_647),
.A2(n_480),
.B1(n_468),
.B2(n_536),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_665),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_630),
.A2(n_608),
.B(n_603),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_779),
.B(n_526),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_678),
.B(n_535),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_639),
.A2(n_535),
.B1(n_539),
.B2(n_468),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_625),
.A2(n_487),
.B(n_539),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_678),
.B(n_581),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_624),
.B(n_530),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_686),
.B(n_540),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_624),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_731),
.A2(n_553),
.B(n_530),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_624),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_782),
.Y(n_819)
);

CKINVDCx10_ASAP7_75t_R g820 ( 
.A(n_756),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_703),
.A2(n_615),
.B(n_614),
.C(n_540),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_647),
.A2(n_594),
.B(n_606),
.C(n_595),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_645),
.B(n_553),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_625),
.A2(n_556),
.B(n_567),
.Y(n_824)
);

AND2x6_ASAP7_75t_L g825 ( 
.A(n_776),
.B(n_615),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_625),
.A2(n_556),
.B(n_567),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_628),
.B(n_484),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_751),
.A2(n_615),
.B(n_614),
.C(n_601),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_687),
.B(n_693),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_683),
.A2(n_556),
.B(n_567),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_694),
.B(n_540),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_711),
.B(n_555),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_635),
.A2(n_556),
.B(n_567),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_628),
.B(n_499),
.Y(n_834)
);

CKINVDCx10_ASAP7_75t_R g835 ( 
.A(n_756),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_681),
.A2(n_556),
.B(n_567),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_712),
.B(n_555),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_700),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_621),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_626),
.B(n_499),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_714),
.B(n_555),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_682),
.A2(n_556),
.B(n_567),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_L g843 ( 
.A1(n_708),
.A2(n_314),
.B(n_315),
.Y(n_843)
);

OAI21xp33_ASAP7_75t_L g844 ( 
.A1(n_755),
.A2(n_315),
.B(n_239),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_645),
.B(n_553),
.Y(n_845)
);

OAI21xp33_ASAP7_75t_L g846 ( 
.A1(n_696),
.A2(n_251),
.B(n_244),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_704),
.B(n_652),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_724),
.B(n_555),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_700),
.B(n_240),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_627),
.A2(n_615),
.B(n_614),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_619),
.A2(n_491),
.B(n_501),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_743),
.B(n_745),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_684),
.A2(n_544),
.B(n_601),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_778),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_631),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_691),
.B(n_450),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_717),
.B(n_245),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_685),
.A2(n_544),
.B(n_601),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_705),
.A2(n_544),
.B(n_601),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_763),
.A2(n_765),
.B(n_783),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_649),
.B(n_583),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_649),
.B(n_583),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_754),
.B(n_583),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_757),
.B(n_583),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_632),
.A2(n_614),
.B(n_597),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_748),
.A2(n_544),
.B(n_597),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_633),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_633),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_640),
.A2(n_597),
.B(n_584),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_644),
.A2(n_597),
.B(n_584),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_691),
.B(n_450),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_650),
.A2(n_584),
.B1(n_491),
.B2(n_570),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_651),
.A2(n_584),
.B(n_501),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_654),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_656),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_691),
.B(n_536),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_742),
.B(n_536),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_753),
.A2(n_544),
.B(n_596),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_638),
.A2(n_544),
.B(n_401),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_658),
.B(n_536),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_669),
.A2(n_536),
.B1(n_587),
.B2(n_453),
.Y(n_881)
);

AND3x2_ASAP7_75t_L g882 ( 
.A(n_720),
.B(n_257),
.C(n_456),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_698),
.A2(n_528),
.B(n_570),
.C(n_568),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_641),
.A2(n_401),
.B(n_568),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_717),
.B(n_246),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_653),
.A2(n_433),
.B(n_548),
.C(n_546),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_673),
.A2(n_536),
.B1(n_587),
.B2(n_546),
.Y(n_887)
);

INVx11_ASAP7_75t_L g888 ( 
.A(n_744),
.Y(n_888)
);

AOI21xp33_ASAP7_75t_L g889 ( 
.A1(n_660),
.A2(n_433),
.B(n_512),
.Y(n_889)
);

BUFx4f_ASAP7_75t_L g890 ( 
.A(n_744),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_659),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_679),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_648),
.A2(n_401),
.B(n_548),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_730),
.B(n_493),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_762),
.B(n_249),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_718),
.A2(n_401),
.B(n_534),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_778),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_662),
.A2(n_493),
.B1(n_534),
.B2(n_533),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_646),
.B(n_250),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_666),
.A2(n_510),
.B(n_533),
.C(n_528),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_728),
.A2(n_401),
.B(n_512),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_771),
.A2(n_510),
.B(n_398),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_667),
.B(n_255),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_671),
.A2(n_221),
.B1(n_270),
.B2(n_302),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_655),
.B(n_263),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_699),
.B(n_264),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_653),
.A2(n_436),
.B(n_443),
.C(n_434),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_732),
.B(n_436),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_743),
.B(n_302),
.Y(n_909)
);

INVxp67_ASAP7_75t_SL g910 ( 
.A(n_727),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_672),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_736),
.B(n_443),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_738),
.B(n_740),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_773),
.A2(n_398),
.B(n_402),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_672),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_668),
.A2(n_443),
.B(n_448),
.C(n_447),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_629),
.B(n_271),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_663),
.A2(n_643),
.B(n_642),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_719),
.A2(n_443),
.B(n_439),
.C(n_435),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_629),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_719),
.B(n_443),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_661),
.B(n_273),
.C(n_283),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_769),
.B(n_444),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_620),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_620),
.Y(n_925)
);

BUFx4f_ASAP7_75t_L g926 ( 
.A(n_620),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_689),
.B(n_443),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_664),
.B(n_444),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_760),
.A2(n_448),
.B(n_447),
.C(n_444),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_776),
.A2(n_772),
.B(n_733),
.C(n_692),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_663),
.A2(n_587),
.B(n_402),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_657),
.B(n_284),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_689),
.B(n_444),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_727),
.B(n_447),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_690),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_727),
.A2(n_398),
.B(n_402),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_690),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_642),
.A2(n_587),
.B(n_402),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_643),
.A2(n_434),
.B(n_439),
.C(n_435),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_707),
.A2(n_587),
.B(n_394),
.Y(n_940)
);

AO21x1_ASAP7_75t_L g941 ( 
.A1(n_750),
.A2(n_394),
.B(n_398),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_746),
.A2(n_394),
.B(n_439),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_676),
.B(n_292),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_675),
.B(n_448),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_618),
.A2(n_434),
.B(n_435),
.C(n_439),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_746),
.A2(n_394),
.B(n_435),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_695),
.A2(n_448),
.B(n_447),
.C(n_294),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_679),
.B(n_6),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_620),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_618),
.A2(n_434),
.B(n_9),
.C(n_10),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_697),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_697),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_716),
.B(n_587),
.Y(n_953)
);

NOR3xp33_ASAP7_75t_L g954 ( 
.A(n_761),
.B(n_7),
.C(n_11),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_709),
.A2(n_587),
.B(n_442),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_716),
.B(n_723),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_688),
.B(n_12),
.Y(n_957)
);

AO22x1_ASAP7_75t_L g958 ( 
.A1(n_636),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_723),
.B(n_442),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_721),
.A2(n_442),
.B(n_431),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_729),
.A2(n_442),
.B1(n_431),
.B2(n_423),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_688),
.B(n_14),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_729),
.A2(n_442),
.B(n_431),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_739),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_688),
.B(n_16),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_739),
.B(n_442),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_741),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_SL g968 ( 
.A1(n_874),
.A2(n_809),
.B1(n_897),
.B2(n_949),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_860),
.A2(n_767),
.B(n_741),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_943),
.A2(n_688),
.B1(n_752),
.B2(n_750),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_926),
.B(n_749),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_798),
.A2(n_746),
.B1(n_706),
.B2(n_726),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_905),
.A2(n_767),
.B(n_752),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_906),
.B(n_636),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_786),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_786),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_847),
.B(n_734),
.Y(n_977)
);

NOR2x1_ASAP7_75t_L g978 ( 
.A(n_854),
.B(n_735),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_799),
.A2(n_737),
.B(n_784),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_817),
.A2(n_784),
.B(n_775),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_786),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_932),
.A2(n_713),
.B(n_722),
.C(n_725),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_911),
.Y(n_983)
);

INVxp33_ASAP7_75t_L g984 ( 
.A(n_840),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_911),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_917),
.B(n_781),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_926),
.B(n_764),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_795),
.B(n_764),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_798),
.A2(n_780),
.B1(n_774),
.B2(n_777),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_920),
.B(n_768),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_829),
.A2(n_770),
.B1(n_766),
.B2(n_759),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_787),
.A2(n_770),
.B(n_766),
.C(n_759),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_795),
.B(n_747),
.Y(n_993)
);

NAND2x1p5_ASAP7_75t_L g994 ( 
.A(n_868),
.B(n_791),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_816),
.B(n_747),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_915),
.Y(n_996)
);

INVxp67_ASAP7_75t_L g997 ( 
.A(n_807),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_829),
.B(n_616),
.Y(n_998)
);

BUFx2_ASAP7_75t_SL g999 ( 
.A(n_838),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_819),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_899),
.B(n_616),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_861),
.B(n_442),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_793),
.A2(n_442),
.B(n_431),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_895),
.A2(n_857),
.B1(n_885),
.B2(n_825),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_924),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_850),
.A2(n_442),
.B(n_431),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_808),
.A2(n_431),
.B(n_423),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_862),
.B(n_431),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_903),
.B(n_17),
.Y(n_1009)
);

BUFx12f_ASAP7_75t_L g1010 ( 
.A(n_789),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_800),
.B(n_431),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_891),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_843),
.B(n_19),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_935),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_930),
.A2(n_19),
.B(n_23),
.C(n_27),
.Y(n_1015)
);

OR2x6_ASAP7_75t_SL g1016 ( 
.A(n_922),
.B(n_27),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_844),
.A2(n_431),
.B(n_423),
.C(n_34),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_791),
.Y(n_1018)
);

INVx5_ASAP7_75t_L g1019 ( 
.A(n_825),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_791),
.Y(n_1020)
);

AND2x2_ASAP7_75t_SL g1021 ( 
.A(n_890),
.B(n_31),
.Y(n_1021)
);

BUFx8_ASAP7_75t_L g1022 ( 
.A(n_892),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_804),
.Y(n_1023)
);

O2A1O1Ixp5_ASAP7_75t_L g1024 ( 
.A1(n_918),
.A2(n_785),
.B(n_909),
.C(n_923),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_954),
.A2(n_32),
.B(n_34),
.C(n_36),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_823),
.B(n_423),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_845),
.B(n_423),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_818),
.A2(n_423),
.B1(n_95),
.B2(n_99),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_796),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_790),
.A2(n_423),
.B(n_90),
.Y(n_1030)
);

AO22x1_ASAP7_75t_L g1031 ( 
.A1(n_957),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_951),
.B(n_423),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_804),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_SL g1034 ( 
.A1(n_827),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_SL g1035 ( 
.A(n_846),
.B(n_43),
.C(n_44),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_813),
.A2(n_50),
.B(n_53),
.C(n_58),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_913),
.A2(n_58),
.B(n_71),
.C(n_76),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_937),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_825),
.A2(n_423),
.B1(n_82),
.B2(n_87),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_792),
.A2(n_81),
.B(n_88),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_839),
.B(n_100),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_865),
.A2(n_103),
.B(n_104),
.Y(n_1042)
);

INVx6_ASAP7_75t_L g1043 ( 
.A(n_789),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_925),
.B(n_106),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_855),
.B(n_875),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_856),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_804),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_867),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_964),
.B(n_114),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_849),
.B(n_118),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_834),
.B(n_119),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_805),
.A2(n_127),
.B(n_130),
.C(n_133),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_869),
.A2(n_135),
.B(n_140),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_825),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_967),
.B(n_158),
.Y(n_1055)
);

INVx4_ASAP7_75t_L g1056 ( 
.A(n_867),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_877),
.A2(n_821),
.B(n_828),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_951),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_863),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_825),
.A2(n_803),
.B1(n_856),
.B2(n_871),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_871),
.B(n_794),
.Y(n_1061)
);

INVx3_ASAP7_75t_SL g1062 ( 
.A(n_888),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_867),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_951),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_952),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_952),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_794),
.B(n_952),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_950),
.A2(n_928),
.B(n_965),
.C(n_962),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_801),
.B(n_802),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_801),
.B(n_802),
.Y(n_1070)
);

NOR2x1_ASAP7_75t_SL g1071 ( 
.A(n_868),
.B(n_811),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_948),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_788),
.B(n_806),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_852),
.B(n_864),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_870),
.A2(n_873),
.B(n_960),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_894),
.B(n_797),
.Y(n_1076)
);

OR2x6_ASAP7_75t_L g1077 ( 
.A(n_788),
.B(n_876),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_958),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_933),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_894),
.B(n_797),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_882),
.B(n_814),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_890),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_933),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_956),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_822),
.A2(n_901),
.B(n_896),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_966),
.A2(n_866),
.B(n_940),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_934),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_815),
.B(n_848),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_934),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_SL g1090 ( 
.A1(n_955),
.A2(n_938),
.B(n_878),
.C(n_931),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_963),
.A2(n_853),
.B(n_858),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_815),
.B(n_848),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_880),
.B(n_810),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_889),
.B(n_841),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_908),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_820),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_831),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_831),
.B(n_841),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_883),
.A2(n_953),
.B(n_900),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_889),
.B(n_837),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_947),
.B(n_904),
.C(n_881),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_832),
.Y(n_1102)
);

AOI21x1_ASAP7_75t_L g1103 ( 
.A1(n_851),
.A2(n_959),
.B(n_837),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_908),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_832),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_SL g1106 ( 
.A1(n_886),
.A2(n_812),
.B(n_939),
.C(n_907),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_912),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_910),
.Y(n_1108)
);

BUFx8_ASAP7_75t_SL g1109 ( 
.A(n_835),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_927),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1003),
.A2(n_893),
.B(n_884),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1045),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1003),
.A2(n_859),
.B(n_902),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_SL g1114 ( 
.A(n_1019),
.B(n_1010),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1072),
.B(n_944),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_977),
.B(n_986),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_1065),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_969),
.A2(n_842),
.B(n_830),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_984),
.B(n_941),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_969),
.A2(n_833),
.B(n_836),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1102),
.B(n_921),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1075),
.A2(n_872),
.B(n_826),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1004),
.B(n_953),
.Y(n_1123)
);

AOI31xp67_ASAP7_75t_L g1124 ( 
.A1(n_970),
.A2(n_887),
.A3(n_929),
.B(n_916),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_SL g1125 ( 
.A(n_1019),
.B(n_879),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1012),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1007),
.A2(n_914),
.B(n_936),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1014),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1075),
.A2(n_824),
.B(n_898),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1097),
.B(n_942),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_1109),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1038),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_990),
.B(n_946),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1076),
.A2(n_961),
.B(n_919),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_1000),
.B(n_945),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1076),
.A2(n_1080),
.B(n_1085),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1096),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_973),
.A2(n_1085),
.A3(n_1091),
.B(n_1071),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_997),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1080),
.A2(n_980),
.B(n_1092),
.Y(n_1140)
);

OAI21xp33_ASAP7_75t_L g1141 ( 
.A1(n_1013),
.A2(n_1051),
.B(n_1035),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1095),
.B(n_1104),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_SL g1143 ( 
.A1(n_982),
.A2(n_1050),
.B(n_1088),
.Y(n_1143)
);

O2A1O1Ixp5_ASAP7_75t_L g1144 ( 
.A1(n_1001),
.A2(n_971),
.B(n_1057),
.C(n_1091),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1079),
.B(n_1083),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1061),
.B(n_1059),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_980),
.A2(n_1098),
.B(n_979),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1029),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_974),
.B(n_1078),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1007),
.A2(n_979),
.B(n_1006),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1009),
.B(n_1094),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1094),
.B(n_1100),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1100),
.B(n_1069),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1062),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1060),
.A2(n_1019),
.B1(n_1054),
.B2(n_1073),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1034),
.A2(n_1081),
.B1(n_968),
.B2(n_1031),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1015),
.A2(n_1025),
.B(n_1068),
.C(n_1017),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1006),
.A2(n_1099),
.B(n_1103),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1086),
.A2(n_1026),
.B(n_1027),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_976),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1086),
.A2(n_1090),
.B(n_1070),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1046),
.B(n_1021),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1069),
.B(n_1070),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1036),
.A2(n_1037),
.B(n_987),
.C(n_1041),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_1065),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_1030),
.A2(n_992),
.A3(n_1053),
.B(n_989),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_SL g1167 ( 
.A1(n_1041),
.A2(n_1049),
.B(n_1093),
.C(n_1106),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1024),
.A2(n_1101),
.B(n_972),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1005),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1019),
.A2(n_1108),
.B1(n_998),
.B2(n_1074),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1026),
.A2(n_1027),
.B(n_1008),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_976),
.Y(n_1172)
);

AO32x2_ASAP7_75t_L g1173 ( 
.A1(n_991),
.A2(n_1028),
.A3(n_1056),
.B1(n_975),
.B2(n_1033),
.Y(n_1173)
);

OA21x2_ASAP7_75t_L g1174 ( 
.A1(n_1030),
.A2(n_1053),
.B(n_998),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_978),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_1042),
.A2(n_1040),
.A3(n_1049),
.B(n_988),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1082),
.B(n_1016),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1084),
.A2(n_1110),
.B1(n_1077),
.B2(n_995),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_SL g1179 ( 
.A(n_1039),
.B(n_1052),
.C(n_1040),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_1011),
.A2(n_1008),
.B(n_1002),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_988),
.A2(n_993),
.A3(n_1055),
.B(n_1002),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_999),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1043),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_SL g1184 ( 
.A1(n_1055),
.A2(n_1067),
.B(n_993),
.C(n_1032),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1067),
.A2(n_1105),
.B(n_1077),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1044),
.A2(n_1077),
.B(n_996),
.C(n_985),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_1065),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_R g1188 ( 
.A(n_1043),
.B(n_975),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1044),
.A2(n_983),
.B(n_1064),
.C(n_1058),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1107),
.A2(n_1089),
.B(n_994),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1066),
.B(n_1087),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1018),
.A2(n_1047),
.B(n_1056),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1107),
.A2(n_1047),
.B(n_1018),
.C(n_1089),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1020),
.A2(n_1033),
.A3(n_1107),
.B(n_1089),
.Y(n_1194)
);

AO21x2_ASAP7_75t_L g1195 ( 
.A1(n_976),
.A2(n_981),
.B(n_1023),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1020),
.A2(n_981),
.B(n_1023),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1023),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_SL g1198 ( 
.A1(n_1048),
.A2(n_1063),
.B(n_1044),
.C(n_1043),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1048),
.A2(n_637),
.B(n_982),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1063),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_SL g1201 ( 
.A1(n_1015),
.A2(n_1025),
.B1(n_1013),
.B2(n_675),
.C(n_1036),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1022),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_SL g1203 ( 
.A1(n_982),
.A2(n_518),
.B(n_509),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1003),
.A2(n_851),
.B(n_1007),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1013),
.A2(n_809),
.B1(n_986),
.B2(n_905),
.Y(n_1205)
);

O2A1O1Ixp5_ASAP7_75t_L g1206 ( 
.A1(n_1001),
.A2(n_943),
.B(n_905),
.C(n_1050),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1109),
.Y(n_1207)
);

AOI221xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1015),
.A2(n_1025),
.B1(n_1013),
.B2(n_675),
.C(n_1036),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1013),
.A2(n_809),
.B1(n_986),
.B2(n_905),
.Y(n_1209)
);

OAI22x1_ASAP7_75t_L g1210 ( 
.A1(n_1078),
.A2(n_524),
.B1(n_480),
.B2(n_470),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1050),
.A2(n_637),
.B(n_905),
.C(n_982),
.Y(n_1211)
);

AO21x2_ASAP7_75t_L g1212 ( 
.A1(n_1085),
.A2(n_1057),
.B(n_1091),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_973),
.A2(n_918),
.A3(n_1085),
.B(n_941),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1003),
.A2(n_851),
.B(n_1007),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1003),
.A2(n_851),
.B(n_1007),
.Y(n_1215)
);

AO32x2_ASAP7_75t_L g1216 ( 
.A1(n_1034),
.A2(n_989),
.A3(n_972),
.B1(n_991),
.B2(n_1028),
.Y(n_1216)
);

BUFx5_ASAP7_75t_L g1217 ( 
.A(n_1095),
.Y(n_1217)
);

NOR2xp67_ASAP7_75t_L g1218 ( 
.A(n_1019),
.B(n_1004),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_973),
.A2(n_918),
.A3(n_1085),
.B(n_941),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1013),
.A2(n_809),
.B1(n_986),
.B2(n_905),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1003),
.A2(n_851),
.B(n_1007),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_969),
.A2(n_617),
.B(n_860),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1000),
.B(n_622),
.Y(n_1223)
);

OAI221xp5_ASAP7_75t_L g1224 ( 
.A1(n_1013),
.A2(n_545),
.B1(n_905),
.B2(n_943),
.C(n_655),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_969),
.A2(n_617),
.B(n_860),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1022),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_977),
.B(n_322),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1003),
.A2(n_851),
.B(n_1007),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_969),
.A2(n_617),
.B(n_860),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_973),
.A2(n_918),
.A3(n_1085),
.B(n_941),
.Y(n_1230)
);

OAI22x1_ASAP7_75t_L g1231 ( 
.A1(n_1078),
.A2(n_524),
.B1(n_480),
.B2(n_470),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1000),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1003),
.A2(n_851),
.B(n_1007),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_973),
.A2(n_918),
.A3(n_1085),
.B(n_941),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_973),
.A2(n_918),
.A3(n_1085),
.B(n_941),
.Y(n_1235)
);

BUFx4_ASAP7_75t_SL g1236 ( 
.A(n_1096),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1006),
.A2(n_980),
.B(n_969),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_980),
.A2(n_1057),
.B(n_1075),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_977),
.B(n_637),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_977),
.B(n_637),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_969),
.A2(n_617),
.B(n_860),
.Y(n_1241)
);

CKINVDCx9p33_ASAP7_75t_R g1242 ( 
.A(n_977),
.Y(n_1242)
);

BUFx12f_ASAP7_75t_L g1243 ( 
.A(n_1010),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_973),
.A2(n_918),
.A3(n_1085),
.B(n_941),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_977),
.B(n_322),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1013),
.A2(n_710),
.B1(n_905),
.B2(n_943),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_997),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_977),
.B(n_322),
.Y(n_1248)
);

NAND2x1p5_ASAP7_75t_L g1249 ( 
.A(n_1114),
.B(n_1182),
.Y(n_1249)
);

BUFx4f_ASAP7_75t_SL g1250 ( 
.A(n_1131),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1224),
.A2(n_1248),
.B1(n_1245),
.B2(n_1227),
.Y(n_1251)
);

BUFx10_ASAP7_75t_L g1252 ( 
.A(n_1154),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1160),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1246),
.A2(n_1205),
.B1(n_1209),
.B2(n_1220),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1207),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1116),
.B(n_1205),
.Y(n_1257)
);

BUFx4_ASAP7_75t_SL g1258 ( 
.A(n_1202),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1209),
.A2(n_1220),
.B1(n_1141),
.B2(n_1210),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1141),
.A2(n_1211),
.B1(n_1156),
.B2(n_1143),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1126),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1183),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1139),
.Y(n_1263)
);

OAI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1156),
.A2(n_1151),
.B1(n_1231),
.B2(n_1112),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1132),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1238),
.A2(n_1168),
.B1(n_1179),
.B2(n_1149),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1148),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1162),
.B(n_1115),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1242),
.A2(n_1177),
.B1(n_1175),
.B2(n_1155),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1223),
.A2(n_1163),
.B1(n_1178),
.B2(n_1182),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1247),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1178),
.A2(n_1142),
.B1(n_1153),
.B2(n_1232),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1146),
.B(n_1152),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1194),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1169),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1145),
.B(n_1121),
.Y(n_1276)
);

CKINVDCx11_ASAP7_75t_R g1277 ( 
.A(n_1243),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1135),
.A2(n_1218),
.B1(n_1199),
.B2(n_1189),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1188),
.Y(n_1279)
);

INVx5_ASAP7_75t_L g1280 ( 
.A(n_1172),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1191),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1238),
.A2(n_1212),
.B1(n_1140),
.B2(n_1147),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1212),
.A2(n_1119),
.B1(n_1218),
.B2(n_1133),
.Y(n_1283)
);

OAI22x1_ASAP7_75t_L g1284 ( 
.A1(n_1206),
.A2(n_1191),
.B1(n_1174),
.B2(n_1197),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_1137),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1170),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1186),
.A2(n_1157),
.B1(n_1193),
.B2(n_1123),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1185),
.A2(n_1208),
.B1(n_1201),
.B2(n_1130),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1136),
.A2(n_1174),
.B1(n_1161),
.B2(n_1217),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1217),
.B(n_1208),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1226),
.A2(n_1190),
.B1(n_1134),
.B2(n_1201),
.Y(n_1291)
);

CKINVDCx11_ASAP7_75t_R g1292 ( 
.A(n_1236),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1217),
.A2(n_1216),
.B1(n_1192),
.B2(n_1198),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1180),
.A2(n_1158),
.B1(n_1171),
.B2(n_1159),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1222),
.A2(n_1225),
.B(n_1241),
.Y(n_1295)
);

BUFx4f_ASAP7_75t_SL g1296 ( 
.A(n_1172),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1200),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1216),
.A2(n_1180),
.B1(n_1165),
.B2(n_1117),
.Y(n_1298)
);

BUFx4_ASAP7_75t_R g1299 ( 
.A(n_1188),
.Y(n_1299)
);

INVx3_ASAP7_75t_SL g1300 ( 
.A(n_1172),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1195),
.Y(n_1301)
);

BUFx12f_ASAP7_75t_L g1302 ( 
.A(n_1117),
.Y(n_1302)
);

OAI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1216),
.A2(n_1187),
.B1(n_1165),
.B2(n_1237),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1195),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1150),
.A2(n_1125),
.B1(n_1129),
.B2(n_1229),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1181),
.B(n_1167),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1144),
.A2(n_1187),
.B1(n_1203),
.B2(n_1164),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1122),
.A2(n_1204),
.B1(n_1214),
.B2(n_1221),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1196),
.A2(n_1118),
.B1(n_1120),
.B2(n_1173),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1173),
.A2(n_1184),
.B1(n_1124),
.B2(n_1166),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1113),
.A2(n_1127),
.B1(n_1228),
.B2(n_1215),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1233),
.A2(n_1111),
.B1(n_1166),
.B2(n_1176),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1166),
.A2(n_1173),
.B1(n_1176),
.B2(n_1138),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1176),
.A2(n_1138),
.B1(n_1181),
.B2(n_1213),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1213),
.B(n_1219),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1219),
.A2(n_1230),
.B1(n_1234),
.B2(n_1235),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1230),
.A2(n_1234),
.B1(n_1235),
.B2(n_1244),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1234),
.A2(n_1224),
.B1(n_328),
.B2(n_331),
.Y(n_1318)
);

BUFx8_ASAP7_75t_L g1319 ( 
.A(n_1235),
.Y(n_1319)
);

AOI21xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1244),
.A2(n_1245),
.B(n_1227),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1236),
.Y(n_1321)
);

INVx11_ASAP7_75t_L g1322 ( 
.A(n_1243),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1246),
.A2(n_1205),
.B1(n_1220),
.B2(n_1209),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1223),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1131),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1224),
.A2(n_1246),
.B1(n_1205),
.B2(n_1220),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1205),
.A2(n_1209),
.B1(n_1220),
.B2(n_1239),
.Y(n_1328)
);

BUFx10_ASAP7_75t_L g1329 ( 
.A(n_1154),
.Y(n_1329)
);

INVx8_ASAP7_75t_L g1330 ( 
.A(n_1160),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1194),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1205),
.A2(n_1209),
.B1(n_1220),
.B2(n_1239),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1162),
.B(n_467),
.Y(n_1333)
);

INVx11_ASAP7_75t_L g1334 ( 
.A(n_1243),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1183),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1160),
.Y(n_1336)
);

CKINVDCx6p67_ASAP7_75t_R g1337 ( 
.A(n_1243),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_1243),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1224),
.A2(n_1246),
.B1(n_1205),
.B2(n_1220),
.Y(n_1339)
);

CKINVDCx11_ASAP7_75t_R g1340 ( 
.A(n_1131),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1224),
.A2(n_328),
.B1(n_331),
.B2(n_322),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1205),
.A2(n_1209),
.B1(n_1220),
.B2(n_1239),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1246),
.B(n_1205),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1160),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1131),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1224),
.A2(n_1205),
.B1(n_1220),
.B2(n_1209),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1139),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1139),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1128),
.Y(n_1352)
);

CKINVDCx11_ASAP7_75t_R g1353 ( 
.A(n_1131),
.Y(n_1353)
);

CKINVDCx11_ASAP7_75t_R g1354 ( 
.A(n_1131),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1224),
.A2(n_1246),
.B1(n_1205),
.B2(n_1220),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1224),
.A2(n_1246),
.B1(n_1205),
.B2(n_1220),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1246),
.A2(n_1205),
.B1(n_1220),
.B2(n_1209),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1139),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1128),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1162),
.B(n_467),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1224),
.A2(n_1246),
.B1(n_1205),
.B2(n_1220),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1224),
.A2(n_1246),
.B1(n_1205),
.B2(n_1220),
.Y(n_1362)
);

INVxp67_ASAP7_75t_SL g1363 ( 
.A(n_1272),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1292),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1295),
.A2(n_1306),
.B(n_1309),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1301),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1304),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1315),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1340),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1266),
.B(n_1268),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1319),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1319),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1273),
.B(n_1328),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1290),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1308),
.A2(n_1289),
.B(n_1305),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1275),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1270),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1297),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1249),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1274),
.B(n_1331),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1255),
.B(n_1327),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1308),
.A2(n_1289),
.B(n_1305),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1278),
.B(n_1284),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1266),
.B(n_1259),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1312),
.A2(n_1294),
.B(n_1311),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1312),
.A2(n_1294),
.B(n_1282),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1261),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1265),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1310),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1324),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1326),
.A2(n_1362),
.B(n_1361),
.C(n_1339),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1316),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1286),
.B(n_1257),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1359),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1249),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1259),
.B(n_1283),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1344),
.A2(n_1282),
.B(n_1332),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1286),
.B(n_1316),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1267),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1283),
.B(n_1254),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1317),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1280),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1298),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1313),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1314),
.A2(n_1287),
.B(n_1260),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1280),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1254),
.B(n_1333),
.Y(n_1407)
);

INVxp67_ASAP7_75t_L g1408 ( 
.A(n_1263),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1344),
.A2(n_1342),
.B(n_1332),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1251),
.B(n_1360),
.Y(n_1410)
);

OR2x6_ASAP7_75t_L g1411 ( 
.A(n_1323),
.B(n_1357),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1288),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1314),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1349),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1303),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1326),
.A2(n_1362),
.B(n_1361),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_SL g1417 ( 
.A(n_1343),
.B(n_1345),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1358),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1328),
.B(n_1342),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1280),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1351),
.B(n_1348),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1350),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1281),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1271),
.B(n_1341),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1352),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_1347),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1276),
.Y(n_1427)
);

CKINVDCx8_ASAP7_75t_R g1428 ( 
.A(n_1321),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1291),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1339),
.B(n_1355),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1280),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1355),
.A2(n_1356),
.B(n_1307),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1291),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1293),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1264),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1264),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1427),
.B(n_1356),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1404),
.B(n_1320),
.Y(n_1438)
);

OR2x6_ASAP7_75t_L g1439 ( 
.A(n_1383),
.B(n_1279),
.Y(n_1439)
);

A2O1A1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1409),
.A2(n_1318),
.B(n_1269),
.C(n_1335),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1404),
.B(n_1392),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1392),
.B(n_1401),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1394),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1390),
.Y(n_1444)
);

BUFx12f_ASAP7_75t_L g1445 ( 
.A(n_1364),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1379),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1391),
.A2(n_1419),
.B(n_1421),
.C(n_1411),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1397),
.A2(n_1299),
.B(n_1300),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1414),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1398),
.B(n_1262),
.Y(n_1450)
);

A2O1A1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1432),
.A2(n_1410),
.B(n_1419),
.C(n_1405),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1387),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1388),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1411),
.A2(n_1330),
.B(n_1336),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1388),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_SL g1456 ( 
.A1(n_1421),
.A2(n_1325),
.B(n_1256),
.C(n_1285),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1388),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1381),
.B(n_1373),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1411),
.A2(n_1250),
.B1(n_1337),
.B2(n_1296),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1398),
.B(n_1300),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1413),
.B(n_1374),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1399),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1374),
.B(n_1346),
.Y(n_1463)
);

O2A1O1Ixp33_ASAP7_75t_SL g1464 ( 
.A1(n_1371),
.A2(n_1258),
.B(n_1354),
.C(n_1353),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1383),
.B(n_1330),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1411),
.A2(n_1338),
.B1(n_1302),
.B2(n_1277),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1376),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1378),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1386),
.A2(n_1346),
.B(n_1330),
.Y(n_1469)
);

A2O1A1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1432),
.A2(n_1346),
.B(n_1296),
.C(n_1252),
.Y(n_1470)
);

NOR2x1_ASAP7_75t_SL g1471 ( 
.A(n_1383),
.B(n_1253),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1368),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1424),
.B(n_1250),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1411),
.A2(n_1252),
.B(n_1329),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1366),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1405),
.A2(n_1329),
.B(n_1322),
.C(n_1334),
.Y(n_1476)
);

CKINVDCx8_ASAP7_75t_R g1477 ( 
.A(n_1369),
.Y(n_1477)
);

AO21x2_ASAP7_75t_L g1478 ( 
.A1(n_1365),
.A2(n_1375),
.B(n_1382),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1363),
.A2(n_1430),
.B(n_1384),
.Y(n_1479)
);

INVxp33_ASAP7_75t_L g1480 ( 
.A(n_1417),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1373),
.B(n_1417),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1430),
.A2(n_1377),
.B1(n_1416),
.B2(n_1384),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1403),
.B(n_1415),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1371),
.B(n_1372),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1403),
.B(n_1415),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1416),
.A2(n_1400),
.B(n_1435),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1478),
.B(n_1386),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1475),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1453),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1478),
.B(n_1385),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1477),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1475),
.Y(n_1492)
);

OAI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1440),
.A2(n_1436),
.B1(n_1435),
.B2(n_1383),
.C(n_1412),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1455),
.B(n_1457),
.Y(n_1494)
);

CKINVDCx11_ASAP7_75t_R g1495 ( 
.A(n_1445),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1462),
.B(n_1380),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1462),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1461),
.B(n_1412),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1441),
.B(n_1429),
.Y(n_1499)
);

AND2x2_ASAP7_75t_SL g1500 ( 
.A(n_1438),
.B(n_1396),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1468),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1481),
.B(n_1436),
.Y(n_1502)
);

AND2x4_ASAP7_75t_SL g1503 ( 
.A(n_1446),
.B(n_1383),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1478),
.B(n_1385),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1442),
.B(n_1389),
.Y(n_1505)
);

NOR2x1_ASAP7_75t_L g1506 ( 
.A(n_1448),
.B(n_1379),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1449),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1442),
.B(n_1389),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_1477),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1437),
.A2(n_1416),
.B1(n_1400),
.B2(n_1396),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1469),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1452),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1443),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1447),
.B(n_1416),
.C(n_1433),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1472),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1493),
.A2(n_1439),
.B1(n_1448),
.B2(n_1480),
.Y(n_1516)
);

AOI221xp5_ASAP7_75t_L g1517 ( 
.A1(n_1493),
.A2(n_1502),
.B1(n_1451),
.B2(n_1514),
.C(n_1458),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1502),
.B(n_1467),
.Y(n_1518)
);

OAI21xp33_ASAP7_75t_L g1519 ( 
.A1(n_1500),
.A2(n_1480),
.B(n_1438),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1512),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1512),
.Y(n_1521)
);

OAI321xp33_ASAP7_75t_L g1522 ( 
.A1(n_1514),
.A2(n_1486),
.A3(n_1482),
.B1(n_1439),
.B2(n_1465),
.C(n_1479),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1500),
.B(n_1439),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1515),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1488),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1500),
.A2(n_1448),
.B1(n_1439),
.B2(n_1459),
.Y(n_1526)
);

NOR2x1_ASAP7_75t_L g1527 ( 
.A(n_1506),
.B(n_1474),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1489),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1500),
.B(n_1496),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1496),
.B(n_1465),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1496),
.B(n_1465),
.Y(n_1531)
);

OAI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1510),
.A2(n_1466),
.B1(n_1476),
.B2(n_1470),
.C(n_1456),
.Y(n_1532)
);

NAND3xp33_ASAP7_75t_SL g1533 ( 
.A(n_1510),
.B(n_1473),
.C(n_1450),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1496),
.B(n_1483),
.Y(n_1534)
);

OAI21xp33_ASAP7_75t_L g1535 ( 
.A1(n_1506),
.A2(n_1485),
.B(n_1450),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1488),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1503),
.A2(n_1372),
.B1(n_1434),
.B2(n_1484),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1513),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1507),
.B(n_1485),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1511),
.B(n_1471),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1492),
.Y(n_1541)
);

INVx5_ASAP7_75t_L g1542 ( 
.A(n_1511),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1501),
.B(n_1444),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1507),
.B(n_1484),
.Y(n_1544)
);

NAND3xp33_ASAP7_75t_L g1545 ( 
.A(n_1487),
.B(n_1460),
.C(n_1393),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1501),
.A2(n_1498),
.B1(n_1487),
.B2(n_1376),
.C(n_1490),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1492),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1494),
.Y(n_1548)
);

INVx5_ASAP7_75t_L g1549 ( 
.A(n_1511),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1490),
.A2(n_1471),
.B(n_1367),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1497),
.Y(n_1551)
);

NOR2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1498),
.B(n_1445),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1499),
.B(n_1463),
.Y(n_1553)
);

NOR3xp33_ASAP7_75t_L g1554 ( 
.A(n_1495),
.B(n_1454),
.C(n_1395),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1495),
.Y(n_1555)
);

NOR3xp33_ASAP7_75t_SL g1556 ( 
.A(n_1499),
.B(n_1434),
.C(n_1425),
.Y(n_1556)
);

NOR3xp33_ASAP7_75t_L g1557 ( 
.A(n_1490),
.B(n_1395),
.C(n_1393),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1505),
.B(n_1484),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1505),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1525),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1525),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1520),
.B(n_1505),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1528),
.Y(n_1563)
);

INVx6_ASAP7_75t_L g1564 ( 
.A(n_1542),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1548),
.B(n_1511),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1536),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1536),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1517),
.B(n_1446),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1540),
.B(n_1513),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1541),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1533),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1521),
.B(n_1508),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1548),
.B(n_1487),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1551),
.B(n_1515),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1556),
.A2(n_1532),
.B1(n_1516),
.B2(n_1526),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1548),
.B(n_1504),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1528),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1529),
.B(n_1504),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1541),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1529),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1547),
.Y(n_1581)
);

NOR2x1_ASAP7_75t_L g1582 ( 
.A(n_1527),
.B(n_1491),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1538),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1534),
.B(n_1538),
.Y(n_1584)
);

BUFx8_ASAP7_75t_SL g1585 ( 
.A(n_1555),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1542),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1540),
.B(n_1513),
.Y(n_1587)
);

NOR2x1_ASAP7_75t_L g1588 ( 
.A(n_1527),
.B(n_1509),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1551),
.B(n_1489),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1521),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1546),
.B(n_1539),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1547),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1542),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1534),
.B(n_1544),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1542),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1539),
.B(n_1524),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1585),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1564),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1560),
.Y(n_1599)
);

NAND2x1p5_ASAP7_75t_L g1600 ( 
.A(n_1582),
.B(n_1523),
.Y(n_1600)
);

AOI211xp5_ASAP7_75t_L g1601 ( 
.A1(n_1575),
.A2(n_1571),
.B(n_1522),
.C(n_1568),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1582),
.B(n_1552),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_1588),
.Y(n_1603)
);

AOI32xp33_ASAP7_75t_L g1604 ( 
.A1(n_1588),
.A2(n_1519),
.A3(n_1535),
.B1(n_1554),
.B2(n_1523),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1583),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1580),
.B(n_1550),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1571),
.A2(n_1407),
.B1(n_1552),
.B2(n_1370),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1560),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1591),
.B(n_1545),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1561),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1580),
.B(n_1594),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1591),
.B(n_1553),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1564),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1590),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1561),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1596),
.Y(n_1616)
);

OAI21xp33_ASAP7_75t_L g1617 ( 
.A1(n_1575),
.A2(n_1557),
.B(n_1504),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1596),
.B(n_1518),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1594),
.B(n_1544),
.Y(n_1619)
);

NOR2xp67_ASAP7_75t_SL g1620 ( 
.A(n_1564),
.B(n_1428),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1566),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1590),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1594),
.B(n_1543),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1566),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1559),
.B(n_1562),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1578),
.B(n_1530),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1567),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1564),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1559),
.B(n_1558),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1584),
.B(n_1530),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1567),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1583),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1564),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1578),
.B(n_1531),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1570),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1570),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1586),
.B(n_1550),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1579),
.Y(n_1638)
);

NAND2xp33_ASAP7_75t_SL g1639 ( 
.A(n_1584),
.B(n_1426),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1617),
.A2(n_1503),
.B1(n_1540),
.B2(n_1407),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1601),
.B(n_1584),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1603),
.Y(n_1642)
);

CKINVDCx16_ASAP7_75t_R g1643 ( 
.A(n_1639),
.Y(n_1643)
);

NOR2xp67_ASAP7_75t_SL g1644 ( 
.A(n_1609),
.B(n_1428),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1611),
.B(n_1603),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1616),
.B(n_1562),
.Y(n_1646)
);

AOI211xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1622),
.A2(n_1464),
.B(n_1593),
.C(n_1595),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1600),
.B(n_1578),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1600),
.B(n_1569),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1614),
.Y(n_1650)
);

OAI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1602),
.A2(n_1537),
.B1(n_1572),
.B2(n_1595),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1586),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1597),
.B(n_1408),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1623),
.B(n_1558),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1639),
.B(n_1540),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1612),
.B(n_1572),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1623),
.B(n_1579),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1614),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1602),
.B(n_1569),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1602),
.B(n_1569),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1611),
.Y(n_1661)
);

NAND4xp25_ASAP7_75t_L g1662 ( 
.A(n_1604),
.B(n_1607),
.C(n_1633),
.D(n_1618),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1607),
.B(n_1581),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1599),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1606),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1619),
.B(n_1581),
.Y(n_1666)
);

INVxp33_ASAP7_75t_L g1667 ( 
.A(n_1620),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1598),
.B(n_1418),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1619),
.B(n_1592),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1630),
.B(n_1569),
.Y(n_1670)
);

INVxp33_ASAP7_75t_L g1671 ( 
.A(n_1630),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1608),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1629),
.B(n_1592),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1598),
.A2(n_1503),
.B1(n_1550),
.B2(n_1370),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1613),
.B(n_1422),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1643),
.B(n_1648),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1647),
.A2(n_1628),
.B(n_1613),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1650),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1643),
.A2(n_1628),
.B1(n_1605),
.B2(n_1632),
.Y(n_1679)
);

OAI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1641),
.A2(n_1625),
.B1(n_1595),
.B2(n_1593),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1645),
.Y(n_1681)
);

NOR2xp67_ASAP7_75t_SL g1682 ( 
.A(n_1655),
.B(n_1395),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1650),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1656),
.B(n_1605),
.Y(n_1684)
);

AOI222xp33_ASAP7_75t_L g1685 ( 
.A1(n_1642),
.A2(n_1606),
.B1(n_1610),
.B2(n_1636),
.C1(n_1635),
.C2(n_1638),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1644),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1645),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1640),
.A2(n_1634),
.B1(n_1626),
.B2(n_1606),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1645),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1658),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1658),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1664),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1668),
.B(n_1632),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1648),
.B(n_1569),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1664),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1645),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1644),
.B(n_1414),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1661),
.Y(n_1698)
);

AOI21xp33_ASAP7_75t_L g1699 ( 
.A1(n_1667),
.A2(n_1586),
.B(n_1593),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1661),
.B(n_1587),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1675),
.Y(n_1701)
);

NAND2x1p5_ASAP7_75t_L g1702 ( 
.A(n_1687),
.B(n_1659),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1676),
.A2(n_1662),
.B1(n_1651),
.B2(n_1660),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1681),
.B(n_1671),
.Y(n_1704)
);

OAI21xp33_ASAP7_75t_L g1705 ( 
.A1(n_1679),
.A2(n_1663),
.B(n_1660),
.Y(n_1705)
);

OAI321xp33_ASAP7_75t_L g1706 ( 
.A1(n_1680),
.A2(n_1659),
.A3(n_1649),
.B1(n_1665),
.B2(n_1674),
.C(n_1657),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1676),
.A2(n_1649),
.B1(n_1652),
.B2(n_1653),
.Y(n_1707)
);

OAI31xp33_ASAP7_75t_L g1708 ( 
.A1(n_1686),
.A2(n_1646),
.A3(n_1652),
.B(n_1672),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1701),
.A2(n_1654),
.B1(n_1656),
.B2(n_1646),
.Y(n_1709)
);

NAND2x1_ASAP7_75t_L g1710 ( 
.A(n_1687),
.B(n_1652),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_SL g1711 ( 
.A1(n_1688),
.A2(n_1652),
.B(n_1670),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1698),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1699),
.A2(n_1665),
.B(n_1672),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1677),
.A2(n_1673),
.B(n_1669),
.Y(n_1714)
);

AOI31xp33_ASAP7_75t_L g1715 ( 
.A1(n_1697),
.A2(n_1670),
.A3(n_1666),
.B(n_1615),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1681),
.B(n_1621),
.Y(n_1716)
);

NAND2x1_ASAP7_75t_L g1717 ( 
.A(n_1687),
.B(n_1637),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1681),
.B(n_1624),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1698),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1689),
.B(n_1627),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1706),
.A2(n_1683),
.B1(n_1690),
.B2(n_1691),
.C(n_1678),
.Y(n_1721)
);

NAND2x1_ASAP7_75t_L g1722 ( 
.A(n_1707),
.B(n_1687),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1712),
.Y(n_1723)
);

NOR3x1_ASAP7_75t_L g1724 ( 
.A(n_1704),
.B(n_1714),
.C(n_1710),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1703),
.A2(n_1693),
.B1(n_1689),
.B2(n_1696),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1719),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1705),
.A2(n_1690),
.B1(n_1683),
.B2(n_1678),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1709),
.B(n_1689),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1702),
.B(n_1696),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1716),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1718),
.Y(n_1731)
);

XOR2x2_ASAP7_75t_L g1732 ( 
.A(n_1713),
.B(n_1691),
.Y(n_1732)
);

NAND3xp33_ASAP7_75t_L g1733 ( 
.A(n_1721),
.B(n_1708),
.C(n_1696),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1728),
.B(n_1708),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1725),
.B(n_1698),
.Y(n_1735)
);

NOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1722),
.B(n_1692),
.Y(n_1736)
);

NAND3xp33_ASAP7_75t_L g1737 ( 
.A(n_1727),
.B(n_1685),
.C(n_1711),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1729),
.B(n_1715),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1730),
.B(n_1682),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1723),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1731),
.B(n_1682),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1724),
.B(n_1694),
.Y(n_1742)
);

AND3x1_ASAP7_75t_L g1743 ( 
.A(n_1736),
.B(n_1727),
.C(n_1726),
.Y(n_1743)
);

OAI211xp5_ASAP7_75t_L g1744 ( 
.A1(n_1733),
.A2(n_1717),
.B(n_1732),
.C(n_1720),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1735),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1742),
.Y(n_1746)
);

AOI222xp33_ASAP7_75t_L g1747 ( 
.A1(n_1737),
.A2(n_1695),
.B1(n_1692),
.B2(n_1700),
.C1(n_1637),
.C2(n_1694),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1743),
.A2(n_1734),
.B1(n_1739),
.B2(n_1741),
.Y(n_1748)
);

OAI31xp33_ASAP7_75t_L g1749 ( 
.A1(n_1744),
.A2(n_1738),
.A3(n_1740),
.B(n_1695),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1745),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1746),
.A2(n_1700),
.B1(n_1684),
.B2(n_1637),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1745),
.A2(n_1684),
.B1(n_1631),
.B2(n_1583),
.C(n_1565),
.Y(n_1752)
);

OAI22xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1747),
.A2(n_1549),
.B1(n_1542),
.B2(n_1574),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1750),
.Y(n_1754)
);

NOR2x1_ASAP7_75t_SL g1755 ( 
.A(n_1753),
.B(n_1542),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1748),
.B(n_1574),
.Y(n_1756)
);

NAND4xp75_ASAP7_75t_L g1757 ( 
.A(n_1749),
.B(n_1565),
.C(n_1576),
.D(n_1573),
.Y(n_1757)
);

NAND2x1p5_ASAP7_75t_L g1758 ( 
.A(n_1751),
.B(n_1402),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1757),
.A2(n_1752),
.B1(n_1574),
.B2(n_1549),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1754),
.Y(n_1760)
);

NOR2xp67_ASAP7_75t_SL g1761 ( 
.A(n_1756),
.B(n_1423),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1760),
.A2(n_1755),
.B(n_1758),
.Y(n_1762)
);

OAI22x1_ASAP7_75t_L g1763 ( 
.A1(n_1762),
.A2(n_1761),
.B1(n_1759),
.B2(n_1549),
.Y(n_1763)
);

AOI22x1_ASAP7_75t_L g1764 ( 
.A1(n_1763),
.A2(n_1563),
.B1(n_1577),
.B2(n_1565),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1763),
.A2(n_1573),
.B1(n_1576),
.B2(n_1587),
.Y(n_1765)
);

AOI22x1_ASAP7_75t_L g1766 ( 
.A1(n_1764),
.A2(n_1765),
.B1(n_1563),
.B2(n_1577),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1764),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1767),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1766),
.A2(n_1573),
.B(n_1563),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1768),
.B(n_1576),
.Y(n_1770)
);

AO21x2_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1769),
.B(n_1577),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1771),
.Y(n_1772)
);

AOI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1587),
.B1(n_1549),
.B2(n_1589),
.C(n_1423),
.Y(n_1773)
);

AOI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1406),
.B(n_1420),
.C(n_1431),
.Y(n_1774)
);


endmodule