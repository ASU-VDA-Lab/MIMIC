module fake_jpeg_24330_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_31),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_30),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_65),
.B1(n_37),
.B2(n_35),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_55),
.A2(n_21),
.B1(n_25),
.B2(n_38),
.Y(n_104)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_62),
.Y(n_103)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_39),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_64),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_29),
.B1(n_20),
.B2(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_22),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_68),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_74),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_22),
.Y(n_72)
);

OR2x4_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_23),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_33),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_33),
.Y(n_90)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_43),
.B(n_23),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_83),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_0),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_45),
.B1(n_40),
.B2(n_50),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_88),
.A2(n_96),
.B1(n_78),
.B2(n_76),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_71),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_29),
.B1(n_20),
.B2(n_37),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_107),
.B1(n_58),
.B2(n_28),
.Y(n_133)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_114),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_37),
.B1(n_35),
.B2(n_26),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_104),
.B1(n_116),
.B2(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_123),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_45),
.B(n_40),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_21),
.B1(n_38),
.B2(n_25),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_70),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_45),
.B1(n_28),
.B2(n_14),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_28),
.B1(n_16),
.B2(n_13),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_50),
.B1(n_30),
.B2(n_27),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_57),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_54),
.A2(n_28),
.B1(n_30),
.B2(n_18),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_42),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_71),
.B(n_54),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_146),
.C(n_9),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_126),
.B(n_6),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_60),
.C(n_62),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_139),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_18),
.B(n_30),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_130),
.A2(n_132),
.B(n_6),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_61),
.B1(n_58),
.B2(n_67),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_90),
.B(n_108),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_133),
.A2(n_119),
.B1(n_100),
.B2(n_112),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_85),
.B(n_56),
.C(n_42),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_149),
.B1(n_115),
.B2(n_92),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_82),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_57),
.B1(n_85),
.B2(n_56),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_0),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_157),
.B(n_159),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_18),
.B(n_19),
.C(n_27),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_104),
.B(n_27),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_0),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_1),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_148),
.B(n_156),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_94),
.A2(n_27),
.B1(n_19),
.B2(n_10),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_102),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_153),
.B1(n_114),
.B2(n_87),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_19),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_120),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_99),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_113),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_158),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_97),
.B(n_5),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_93),
.B(n_5),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_163),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_164),
.A2(n_166),
.B1(n_179),
.B2(n_154),
.Y(n_209)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_169),
.Y(n_200)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_92),
.B(n_93),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_177),
.B(n_192),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_172),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_113),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_184),
.B1(n_164),
.B2(n_188),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_133),
.A2(n_151),
.B1(n_125),
.B2(n_146),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_175),
.B(n_187),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_115),
.B1(n_95),
.B2(n_89),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_176),
.A2(n_191),
.B1(n_128),
.B2(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_183),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_119),
.B1(n_100),
.B2(n_105),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_119),
.B(n_89),
.C(n_87),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_190),
.B1(n_137),
.B2(n_124),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_126),
.B(n_95),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_156),
.Y(n_222)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_112),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_148),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_126),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_131),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_142),
.B(n_159),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_209),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_196),
.A2(n_198),
.B1(n_223),
.B2(n_168),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_174),
.B1(n_189),
.B2(n_187),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_190),
.A2(n_146),
.B1(n_129),
.B2(n_128),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_199),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_206),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_132),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_221),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_170),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_160),
.B(n_161),
.Y(n_229)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_126),
.A3(n_153),
.B1(n_147),
.B2(n_142),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_185),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_210),
.B(n_212),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_185),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_215),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_175),
.B(n_162),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_171),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_150),
.B1(n_158),
.B2(n_124),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_165),
.A2(n_135),
.B1(n_154),
.B2(n_142),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_135),
.B1(n_159),
.B2(n_127),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_159),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_181),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_161),
.A2(n_127),
.B1(n_8),
.B2(n_6),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_225),
.B(n_234),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_167),
.C(n_172),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_235),
.C(n_247),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_193),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_233),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_229),
.A2(n_240),
.B(n_194),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_160),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_177),
.C(n_163),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_212),
.Y(n_250)
);

BUFx4f_ASAP7_75t_SL g238 ( 
.A(n_221),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_238),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_183),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_239),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_242),
.B1(n_195),
.B2(n_219),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_162),
.B(n_169),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_176),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_199),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_200),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_202),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_166),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_246),
.B(n_210),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_181),
.C(n_191),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_254),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_260),
.B1(n_226),
.B2(n_205),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_244),
.A2(n_216),
.B1(n_201),
.B2(n_213),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_253),
.A2(n_263),
.B(n_229),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_257),
.Y(n_282)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_224),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_232),
.A2(n_207),
.B1(n_194),
.B2(n_215),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_220),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_267),
.Y(n_283)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_223),
.Y(n_284)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_196),
.B1(n_201),
.B2(n_205),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_241),
.B1(n_247),
.B2(n_243),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_202),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_206),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_227),
.C(n_232),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_278),
.C(n_257),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_244),
.B(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_271),
.B(n_273),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_267),
.B1(n_260),
.B2(n_270),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_274),
.A2(n_279),
.B1(n_284),
.B2(n_265),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_261),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_250),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_256),
.B(n_235),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_277),
.B(n_285),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_224),
.C(n_222),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_233),
.B1(n_228),
.B2(n_217),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_214),
.Y(n_285)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_269),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_272),
.B1(n_284),
.B2(n_274),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_282),
.C(n_286),
.Y(n_303)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_248),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_297),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_254),
.B1(n_253),
.B2(n_248),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_259),
.Y(n_297)
);

FAx1_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_9),
.CI(n_11),
.CON(n_298),
.SN(n_298)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_16),
.C(n_11),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_285),
.C(n_276),
.Y(n_301)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_309),
.C(n_299),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_307),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_295),
.B1(n_288),
.B2(n_294),
.Y(n_307)
);

AOI221xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_297),
.B1(n_293),
.B2(n_280),
.C(n_271),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_281),
.C(n_280),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_289),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_300),
.B(n_268),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_314),
.Y(n_319)
);

INVx11_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_291),
.C(n_281),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_318),
.A2(n_314),
.B1(n_296),
.B2(n_313),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_320),
.B(n_298),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_323),
.A2(n_321),
.B(n_318),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_311),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_316),
.C(n_319),
.Y(n_328)
);

OAI321xp33_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_326),
.A3(n_315),
.B1(n_325),
.B2(n_317),
.C(n_313),
.Y(n_329)
);

AOI21xp33_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_306),
.B(n_287),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_306),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_13),
.B1(n_16),
.B2(n_322),
.Y(n_332)
);


endmodule