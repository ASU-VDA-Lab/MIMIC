module real_jpeg_28717_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_334, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_334;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx5_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_2),
.A2(n_27),
.B1(n_35),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_2),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_2),
.A2(n_31),
.B1(n_33),
.B2(n_184),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_184),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_2),
.A2(n_63),
.B1(n_65),
.B2(n_184),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_4),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_4),
.B(n_30),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_4),
.B(n_33),
.Y(n_221)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_4),
.A2(n_33),
.B(n_221),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_182),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_4),
.A2(n_60),
.B(n_63),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_4),
.B(n_88),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_4),
.A2(n_111),
.B1(n_129),
.B2(n_269),
.Y(n_271)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_6),
.A2(n_31),
.B1(n_33),
.B2(n_38),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_6),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_6),
.A2(n_38),
.B1(n_63),
.B2(n_65),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_7),
.A2(n_27),
.B1(n_35),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_7),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_7),
.A2(n_31),
.B1(n_33),
.B2(n_150),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_150),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_7),
.A2(n_63),
.B1(n_65),
.B2(n_150),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_8),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_8),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_8),
.A2(n_36),
.B1(n_63),
.B2(n_65),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_9),
.A2(n_31),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_9),
.A2(n_27),
.B1(n_35),
.B2(n_53),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_9),
.A2(n_53),
.B1(n_63),
.B2(n_65),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_134)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_31),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_11),
.A2(n_50),
.B1(n_63),
.B2(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_11),
.A2(n_27),
.B1(n_35),
.B2(n_50),
.Y(n_125)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_13),
.A2(n_31),
.B1(n_33),
.B2(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_14),
.A2(n_27),
.B1(n_35),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_14),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_14),
.A2(n_31),
.B1(n_33),
.B2(n_123),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_123),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_14),
.A2(n_63),
.B1(n_65),
.B2(n_123),
.Y(n_256)
);

INVx11_ASAP7_75t_SL g64 ( 
.A(n_15),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_95),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_80),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_74),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_40),
.B1(n_41),
.B2(n_69),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_23),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_23),
.A2(n_39),
.B1(n_122),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_23),
.A2(n_39),
.B1(n_149),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_24),
.B(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_24),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_24),
.A2(n_85),
.B(n_125),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_24),
.A2(n_30),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_25),
.B(n_33),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g181 ( 
.A(n_27),
.B(n_182),
.CON(n_181),
.SN(n_181)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_29),
.A2(n_31),
.B1(n_181),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_30),
.B(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_31),
.A2(n_46),
.A3(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_34),
.A2(n_39),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_39),
.B(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_57),
.B2(n_68),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_43),
.B(n_57),
.C(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_51),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_44),
.A2(n_76),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_45),
.A2(n_54),
.B1(n_78),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_45),
.A2(n_54),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_45),
.A2(n_54),
.B1(n_178),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_45),
.A2(n_54),
.B1(n_206),
.B2(n_225),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g222 ( 
.A(n_47),
.B(n_220),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_47),
.A2(n_61),
.B(n_182),
.C(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_51),
.A2(n_88),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_56),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_57),
.A2(n_68),
.B1(n_75),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_66),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_58),
.A2(n_62),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_115),
.B(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_58),
.A2(n_66),
.B(n_133),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_58),
.A2(n_62),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_58),
.A2(n_156),
.B(n_229),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_58),
.A2(n_62),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_58),
.A2(n_62),
.B1(n_228),
.B2(n_246),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_62),
.A2(n_114),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_62),
.B(n_182),
.Y(n_267)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_65),
.B(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_67),
.B(n_135),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.C(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_70),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_70),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_74),
.B(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_75),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_79),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_76),
.A2(n_79),
.B(n_89),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI321xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_313),
.A3(n_325),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_167),
.B(n_312),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_151),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_98),
.B(n_151),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_126),
.C(n_137),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_99),
.A2(n_100),
.B1(n_126),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_116),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_101),
.B(n_118),
.C(n_120),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_102),
.B(n_113),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_103),
.A2(n_130),
.B(n_197),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_104),
.A2(n_112),
.B(n_142),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_104),
.A2(n_110),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_111),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_109),
.A2(n_129),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_111),
.A2(n_129),
.B1(n_261),
.B2(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_111),
.B(n_182),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_126),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_136),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_128),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_132),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_128),
.A2(n_161),
.B(n_164),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_129),
.A2(n_130),
.B1(n_140),
.B2(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_134),
.B(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_137),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_146),
.C(n_147),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_138),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_143),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_146),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_165),
.B2(n_166),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_154),
.B(n_160),
.C(n_166),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B(n_159),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_157),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_159),
.B(n_315),
.C(n_321),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_159),
.A2(n_315),
.B1(n_316),
.B2(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_159),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_165),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_306),
.B(n_311),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_210),
.B(n_292),
.C(n_305),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_198),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_170),
.B(n_198),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_185),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_172),
.B(n_173),
.C(n_185),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_180),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_187),
.B(n_191),
.C(n_193),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_196),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.C(n_204),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_199),
.A2(n_200),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_204),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.C(n_209),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_291),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_284),
.B(n_290),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_239),
.B(n_283),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_230),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_214),
.B(n_230),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.C(n_226),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_215),
.A2(n_216),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_218),
.Y(n_237)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_231),
.B(n_237),
.C(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_277),
.B(n_282),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_257),
.B(n_276),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_242),
.B(n_249),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_255),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_256),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_265),
.B(n_275),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_263),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_270),
.B(n_274),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_285),
.B(n_286),
.Y(n_290)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_294),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_303),
.B2(n_304),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_300),
.C(n_304),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_323),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_321),
.A2(n_322),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);


endmodule