module fake_aes_1505_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_16;
wire n_25;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_8), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_4), .Y(n_13) );
INVxp67_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
OA21x2_ASAP7_75t_L g15 ( .A1(n_1), .A2(n_2), .B(n_9), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_16), .B(n_1), .Y(n_19) );
NAND3xp33_ASAP7_75t_L g20 ( .A(n_12), .B(n_7), .C(n_3), .Y(n_20) );
OR2x6_ASAP7_75t_L g21 ( .A(n_12), .B(n_2), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_18), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_14), .B(n_3), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_17), .Y(n_24) );
INVx2_ASAP7_75t_SL g25 ( .A(n_24), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_22), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_21), .A2(n_11), .B1(n_13), .B2(n_15), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_21), .B(n_15), .Y(n_28) );
AOI22xp33_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_23), .B1(n_19), .B2(n_15), .Y(n_29) );
BUFx3_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
OAI21x1_ASAP7_75t_L g31 ( .A1(n_27), .A2(n_16), .B(n_20), .Y(n_31) );
INVx1_ASAP7_75t_SL g32 ( .A(n_30), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_32), .B(n_25), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_33), .B(n_30), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_26), .B1(n_27), .B2(n_25), .Y(n_37) );
AND2x2_ASAP7_75t_L g38 ( .A(n_35), .B(n_31), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_37), .B(n_36), .Y(n_39) );
CKINVDCx5p33_ASAP7_75t_R g40 ( .A(n_38), .Y(n_40) );
CKINVDCx20_ASAP7_75t_R g41 ( .A(n_40), .Y(n_41) );
OAI221xp5_ASAP7_75t_R g42 ( .A1(n_41), .A2(n_29), .B1(n_5), .B2(n_4), .C(n_39), .Y(n_42) );
endmodule