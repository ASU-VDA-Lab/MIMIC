module fake_jpeg_26999_n_170 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx11_ASAP7_75t_SL g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_3),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx24_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_72),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_92),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_79),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_55),
.B1(n_50),
.B2(n_60),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_62),
.B1(n_67),
.B2(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_97),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_92),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_59),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_67),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_48),
.B1(n_58),
.B2(n_71),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_49),
.B1(n_53),
.B2(n_65),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_49),
.B1(n_61),
.B2(n_63),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_108),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_80),
.B1(n_82),
.B2(n_94),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_113),
.B1(n_116),
.B2(n_95),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_48),
.B(n_64),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_68),
.B(n_47),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_101),
.B1(n_58),
.B2(n_87),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_68),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_0),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_126),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_27),
.C(n_39),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_112),
.B(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_1),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_126),
.B(n_119),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_139),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_137),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_143),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_26),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_145),
.B1(n_4),
.B2(n_5),
.Y(n_155)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_70),
.B1(n_56),
.B2(n_51),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_148),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_21),
.B1(n_37),
.B2(n_36),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_152),
.A2(n_154),
.B(n_155),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_142),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_153),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_140),
.B(n_141),
.C(n_143),
.D(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_160),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_150),
.B1(n_155),
.B2(n_146),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_158),
.C(n_149),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_146),
.B(n_25),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_18),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_28),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_17),
.C(n_38),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_15),
.A3(n_35),
.B1(n_34),
.B2(n_32),
.C1(n_31),
.C2(n_30),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_151),
.C(n_29),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_11),
.B(n_7),
.Y(n_170)
);


endmodule