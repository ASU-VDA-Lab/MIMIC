module fake_ariane_453_n_1699 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1699);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1699;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_19),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_72),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_88),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_21),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_37),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_44),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_43),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_56),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_63),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_41),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_9),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_82),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_98),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_83),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_116),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_28),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_62),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_8),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_139),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_96),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_94),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_108),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_64),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_92),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_104),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_24),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_42),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_11),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_54),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_77),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_44),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_20),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_15),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_17),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_15),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_67),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_133),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_70),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_68),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_43),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_132),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_127),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_36),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_23),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_36),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_18),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_100),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_71),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_2),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_142),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_39),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_49),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_144),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_134),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_0),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_90),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_33),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_95),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_6),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_85),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_35),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_23),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_145),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_117),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_111),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_3),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_5),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_14),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_54),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_1),
.Y(n_235)
);

BUFx2_ASAP7_75t_SL g236 ( 
.A(n_1),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_17),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_7),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_32),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_26),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_124),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_143),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_107),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_66),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_91),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_69),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_32),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_103),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_4),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_51),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_58),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_76),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_118),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_136),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_47),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_89),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_138),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_49),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_61),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_125),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_81),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_135),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_53),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_87),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_20),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_12),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_78),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_86),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_120),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_73),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_84),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_130),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_101),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_39),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_146),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_37),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_105),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_55),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_137),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_3),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_75),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_112),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_121),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_80),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_31),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_33),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_25),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_115),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_24),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_148),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_11),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_110),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_126),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_97),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_123),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_45),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_2),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_119),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_12),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_0),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_93),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_150),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_141),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_52),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_122),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_51),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_13),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_57),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_79),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_55),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_46),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_27),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_60),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_46),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_129),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_38),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_310),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_158),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_166),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_218),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_166),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_196),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_158),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_271),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_162),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_168),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_5),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_185),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_168),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_155),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_177),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_234),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_299),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_170),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_239),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_159),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_170),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_299),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_161),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_183),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_183),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_192),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_163),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_291),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_175),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_222),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_177),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_191),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_186),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_247),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_192),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_193),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_191),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_193),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_206),
.B(n_6),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_191),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_177),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_194),
.B(n_202),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_187),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_194),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_190),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_202),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_177),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_198),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_205),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_209),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_210),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_215),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_205),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_216),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_211),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_219),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_223),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_225),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_177),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_164),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_226),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_229),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_208),
.B(n_7),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_208),
.B(n_251),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_211),
.B(n_9),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_232),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_235),
.Y(n_384)
);

BUFx6f_ASAP7_75t_SL g385 ( 
.A(n_242),
.Y(n_385)
);

INVxp33_ASAP7_75t_SL g386 ( 
.A(n_236),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_220),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_220),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_236),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_230),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_213),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_230),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_237),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_241),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_241),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_243),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_251),
.B(n_10),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_243),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_238),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_249),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_245),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_245),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_255),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_263),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_252),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_297),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_325),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_348),
.B(n_252),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_254),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_351),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_364),
.B(n_254),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_297),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g417 ( 
.A1(n_318),
.A2(n_264),
.B(n_260),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_404),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_320),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_318),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_381),
.B(n_300),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_323),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_360),
.Y(n_424)
);

NAND2xp33_ASAP7_75t_R g425 ( 
.A(n_317),
.B(n_274),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_323),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_324),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_390),
.B(n_300),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_359),
.B(n_260),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_R g431 ( 
.A(n_331),
.B(n_156),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_326),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_337),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_329),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_358),
.B(n_213),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_335),
.B(n_338),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_335),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_338),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_341),
.B(n_164),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_341),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_358),
.B(n_264),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_342),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_342),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_321),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_343),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_343),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_352),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_352),
.B(n_268),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_319),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_355),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_349),
.B(n_224),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_362),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_340),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_361),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_361),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_344),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_319),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_363),
.B(n_169),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_382),
.A2(n_366),
.B(n_363),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_366),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_346),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_370),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_328),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_350),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_330),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_372),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_372),
.B(n_268),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_367),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_333),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g477 ( 
.A(n_356),
.B(n_213),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_392),
.B(n_169),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_365),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_394),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_270),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g482 ( 
.A(n_436),
.B(n_356),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_436),
.B(n_270),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_418),
.B(n_334),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_275),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_429),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_411),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_439),
.B(n_275),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_414),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_429),
.B(n_349),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_421),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_413),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_432),
.Y(n_493)
);

AO21x2_ASAP7_75t_L g494 ( 
.A1(n_435),
.A2(n_248),
.B(n_298),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_418),
.B(n_339),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_452),
.A2(n_327),
.B1(n_386),
.B2(n_354),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_413),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_409),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_430),
.A2(n_389),
.B1(n_330),
.B2(n_285),
.Y(n_499)
);

BUFx8_ASAP7_75t_SL g500 ( 
.A(n_424),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_443),
.Y(n_501)
);

CKINVDCx6p67_ASAP7_75t_R g502 ( 
.A(n_409),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_421),
.Y(n_503)
);

BUFx10_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_432),
.Y(n_505)
);

INVxp33_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_426),
.B(n_369),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_467),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_426),
.B(n_371),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_432),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_442),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_446),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_435),
.B(n_395),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_476),
.B(n_336),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_L g516 ( 
.A(n_426),
.B(n_213),
.Y(n_516)
);

BUFx6f_ASAP7_75t_SL g517 ( 
.A(n_428),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_442),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_426),
.B(n_373),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_430),
.B(n_385),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_439),
.B(n_298),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_426),
.B(n_374),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_445),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_443),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_476),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_416),
.B(n_406),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_416),
.B(n_406),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_451),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_451),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_443),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_426),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_426),
.B(n_375),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_448),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_426),
.B(n_378),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_450),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_457),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_450),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_457),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_417),
.A2(n_401),
.B1(n_405),
.B2(n_396),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_452),
.A2(n_385),
.B1(n_383),
.B2(n_403),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_457),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_432),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_410),
.B(n_415),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_450),
.B(n_384),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_450),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_450),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_446),
.B(n_395),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_449),
.B(n_393),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_459),
.B(n_399),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_453),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_417),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_456),
.Y(n_553)
);

OR2x2_ASAP7_75t_SL g554 ( 
.A(n_465),
.B(n_368),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_450),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_414),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_458),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_416),
.B(n_422),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_462),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_415),
.B(n_400),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_447),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_467),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_463),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_449),
.A2(n_306),
.B1(n_278),
.B2(n_289),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_424),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_471),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_447),
.B(n_396),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_450),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_417),
.A2(n_405),
.B1(n_402),
.B2(n_401),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_471),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_470),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_447),
.B(n_398),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_470),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_414),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_464),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_444),
.B(n_377),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_474),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_417),
.A2(n_402),
.B1(n_398),
.B2(n_397),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_474),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_475),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_466),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_471),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_L g583 ( 
.A(n_464),
.B(n_301),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_444),
.B(n_250),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_479),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_447),
.B(n_347),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_475),
.Y(n_587)
);

AND2x6_ASAP7_75t_L g588 ( 
.A(n_439),
.B(n_301),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_480),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_468),
.B(n_302),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_480),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_420),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_468),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_464),
.B(n_302),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_448),
.A2(n_380),
.B1(n_287),
.B2(n_286),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_468),
.B(n_303),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_480),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_468),
.B(n_357),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_464),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_460),
.B(n_303),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_417),
.A2(n_434),
.B1(n_423),
.B2(n_437),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_434),
.B(n_437),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_464),
.B(n_305),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_477),
.A2(n_425),
.B1(n_422),
.B2(n_379),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_578),
.B(n_417),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_487),
.B(n_427),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_492),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_491),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_489),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_497),
.B(n_322),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_484),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_543),
.B(n_422),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_484),
.B(n_465),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_503),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_489),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_574),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_574),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_543),
.B(n_533),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_560),
.B(n_440),
.Y(n_620)
);

NAND3xp33_ASAP7_75t_L g621 ( 
.A(n_560),
.B(n_425),
.C(n_464),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_540),
.B(n_431),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_505),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_549),
.B(n_424),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_482),
.A2(n_485),
.B1(n_483),
.B2(n_488),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_598),
.B(n_586),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_483),
.A2(n_485),
.B1(n_521),
.B2(n_488),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_482),
.A2(n_460),
.B1(n_478),
.B2(n_473),
.Y(n_628)
);

BUFx5_ASAP7_75t_L g629 ( 
.A(n_561),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_496),
.B(n_454),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_562),
.B(n_454),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_483),
.A2(n_440),
.B1(n_473),
.B2(n_428),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_505),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_592),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_486),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_520),
.B(n_473),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_604),
.B(n_472),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_512),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_490),
.B(n_481),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_542),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_585),
.B(n_472),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_495),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_567),
.B(n_572),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_506),
.B(n_576),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_506),
.B(n_472),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_508),
.B(n_345),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_567),
.B(n_478),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_518),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_572),
.A2(n_461),
.B(n_481),
.C(n_469),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_550),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_526),
.B(n_428),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_498),
.Y(n_653)
);

BUFx5_ASAP7_75t_L g654 ( 
.A(n_561),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_523),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_514),
.B(n_461),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_565),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_488),
.B(n_521),
.Y(n_658)
);

INVxp33_ASAP7_75t_L g659 ( 
.A(n_515),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_488),
.B(n_461),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_526),
.B(n_428),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_493),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_548),
.A2(n_287),
.B(n_240),
.C(n_233),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_528),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_563),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_488),
.B(n_428),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_521),
.B(n_464),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_529),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_527),
.Y(n_669)
);

INVx8_ASAP7_75t_L g670 ( 
.A(n_482),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_493),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_504),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_504),
.B(n_296),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_588),
.B(n_408),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_558),
.B(n_312),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_588),
.B(n_412),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_551),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_547),
.B(n_314),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_511),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_588),
.B(n_419),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_SL g681 ( 
.A1(n_482),
.A2(n_221),
.B1(n_266),
.B2(n_265),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_558),
.B(n_188),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_511),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_588),
.B(n_412),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_517),
.B(n_316),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_547),
.B(n_581),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_517),
.B(n_188),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_581),
.B(n_157),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_527),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_486),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_588),
.B(n_315),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_600),
.B(n_195),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_553),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_525),
.Y(n_694)
);

BUFx12f_ASAP7_75t_SL g695 ( 
.A(n_500),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_600),
.B(n_195),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_578),
.A2(n_221),
.B1(n_313),
.B2(n_203),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_552),
.Y(n_698)
);

OR2x6_ASAP7_75t_L g699 ( 
.A(n_584),
.B(n_197),
.Y(n_699)
);

NOR3xp33_ASAP7_75t_L g700 ( 
.A(n_499),
.B(n_203),
.C(n_197),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_SL g701 ( 
.A1(n_482),
.A2(n_231),
.B1(n_276),
.B2(n_313),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_502),
.B(n_231),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_600),
.B(n_233),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_600),
.Y(n_704)
);

INVx8_ASAP7_75t_L g705 ( 
.A(n_600),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_559),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_483),
.A2(n_276),
.B1(n_265),
.B2(n_311),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_485),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_525),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_571),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_595),
.A2(n_280),
.B1(n_311),
.B2(n_286),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_513),
.B(n_258),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_500),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_593),
.B(n_304),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_593),
.B(n_304),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_539),
.B(n_160),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_501),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_564),
.B(n_539),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_590),
.A2(n_307),
.B(n_308),
.C(n_309),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_573),
.B(n_307),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_507),
.B(n_510),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_554),
.Y(n_722)
);

NOR3xp33_ASAP7_75t_L g723 ( 
.A(n_595),
.B(n_308),
.C(n_309),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_577),
.B(n_165),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_579),
.B(n_171),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_580),
.B(n_172),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_590),
.A2(n_244),
.B(n_207),
.C(n_182),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_569),
.B(n_407),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_587),
.B(n_10),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_507),
.B(n_14),
.Y(n_730)
);

INVx8_ASAP7_75t_L g731 ( 
.A(n_535),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_524),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_510),
.B(n_16),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_602),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_519),
.B(n_522),
.Y(n_735)
);

NOR2xp67_ASAP7_75t_SL g736 ( 
.A(n_634),
.B(n_665),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_635),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_613),
.B(n_569),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_657),
.Y(n_739)
);

NOR2x1p5_ASAP7_75t_SL g740 ( 
.A(n_629),
.B(n_530),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_619),
.A2(n_522),
.B(n_519),
.Y(n_741)
);

OAI21xp5_ASAP7_75t_L g742 ( 
.A1(n_660),
.A2(n_601),
.B(n_596),
.Y(n_742)
);

O2A1O1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_606),
.A2(n_596),
.B(n_532),
.C(n_534),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_608),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_640),
.B(n_494),
.Y(n_745)
);

NAND3xp33_ASAP7_75t_L g746 ( 
.A(n_631),
.B(n_534),
.C(n_532),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_627),
.A2(n_601),
.B1(n_589),
.B2(n_541),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_650),
.A2(n_566),
.B(n_536),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_644),
.A2(n_544),
.B(n_599),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_653),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_689),
.B(n_494),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_689),
.B(n_538),
.Y(n_752)
);

CKINVDCx8_ASAP7_75t_R g753 ( 
.A(n_694),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_730),
.A2(n_733),
.B(n_620),
.C(n_640),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_627),
.A2(n_591),
.B1(n_570),
.B2(n_597),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_L g756 ( 
.A(n_629),
.B(n_535),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_637),
.A2(n_544),
.B(n_599),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_626),
.B(n_582),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_645),
.B(n_594),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_656),
.A2(n_546),
.B(n_537),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_730),
.A2(n_603),
.B(n_594),
.C(n_583),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_625),
.A2(n_603),
.B1(n_575),
.B2(n_568),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_670),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_700),
.A2(n_648),
.B(n_711),
.C(n_712),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_718),
.A2(n_701),
.B1(n_681),
.B2(n_733),
.Y(n_765)
);

OA21x2_ASAP7_75t_L g766 ( 
.A1(n_727),
.A2(n_167),
.B(n_182),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_635),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_735),
.A2(n_531),
.B(n_516),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_735),
.A2(n_555),
.B(n_546),
.C(n_545),
.Y(n_769)
);

AOI33xp33_ASAP7_75t_L g770 ( 
.A1(n_682),
.A2(n_167),
.A3(n_207),
.B1(n_244),
.B2(n_414),
.B3(n_407),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_628),
.A2(n_734),
.B(n_721),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_662),
.A2(n_531),
.B(n_174),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_671),
.A2(n_173),
.B(n_295),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_614),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_609),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_635),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_635),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_667),
.A2(n_293),
.B(n_292),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_605),
.A2(n_290),
.B(n_288),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_681),
.A2(n_284),
.B1(n_283),
.B2(n_282),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_657),
.B(n_176),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_605),
.A2(n_281),
.B(n_279),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_669),
.B(n_16),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_714),
.B(n_178),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_670),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_714),
.B(n_179),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_700),
.A2(n_711),
.B(n_719),
.C(n_675),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_670),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_731),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_679),
.A2(n_277),
.B(n_273),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_715),
.B(n_180),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_701),
.B(n_181),
.Y(n_792)
);

BUFx4f_ASAP7_75t_L g793 ( 
.A(n_709),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_621),
.A2(n_272),
.B(n_269),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_R g795 ( 
.A(n_695),
.B(n_184),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_611),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_652),
.B(n_18),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_651),
.B(n_708),
.Y(n_798)
);

OAI21xp33_ASAP7_75t_L g799 ( 
.A1(n_715),
.A2(n_267),
.B(n_262),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_661),
.B(n_19),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_615),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_731),
.Y(n_802)
);

O2A1O1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_675),
.A2(n_21),
.B(n_22),
.C(n_25),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_683),
.A2(n_261),
.B(n_259),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_611),
.B(n_22),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_658),
.A2(n_257),
.B(n_256),
.Y(n_806)
);

OAI22xp33_ASAP7_75t_L g807 ( 
.A1(n_699),
.A2(n_253),
.B1(n_246),
.B2(n_228),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_SL g808 ( 
.A(n_610),
.B(n_227),
.Y(n_808)
);

NAND2x1_ASAP7_75t_L g809 ( 
.A(n_690),
.B(n_698),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_707),
.A2(n_217),
.B1(n_214),
.B2(n_212),
.Y(n_810)
);

AO21x1_ASAP7_75t_L g811 ( 
.A1(n_723),
.A2(n_74),
.B(n_154),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_724),
.A2(n_204),
.B(n_201),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_725),
.A2(n_200),
.B(n_199),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_616),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_731),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_708),
.B(n_189),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_643),
.B(n_26),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_636),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_698),
.B(n_151),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_639),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_617),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_704),
.B(n_632),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_726),
.A2(n_147),
.B(n_140),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_649),
.B(n_27),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_704),
.B(n_28),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_705),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_707),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_655),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_618),
.Y(n_829)
);

OAI21xp33_ASAP7_75t_L g830 ( 
.A1(n_729),
.A2(n_29),
.B(n_30),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_705),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_SL g832 ( 
.A1(n_622),
.A2(n_34),
.B(n_35),
.C(n_38),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_607),
.B(n_699),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_664),
.B(n_668),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_632),
.B(n_40),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_698),
.Y(n_836)
);

BUFx12f_ASAP7_75t_L g837 ( 
.A(n_672),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_729),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_677),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_717),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_713),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_693),
.A2(n_47),
.B(n_48),
.C(n_50),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_702),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_647),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_697),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_607),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_706),
.B(n_58),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_710),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_687),
.B(n_128),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_723),
.A2(n_692),
.B(n_696),
.C(n_703),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_720),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_674),
.A2(n_680),
.B(n_684),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_705),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_713),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_732),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_676),
.A2(n_623),
.B(n_633),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_682),
.B(n_699),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_646),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_641),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_663),
.A2(n_624),
.B(n_678),
.C(n_673),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_666),
.B(n_685),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_716),
.A2(n_691),
.B(n_728),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_722),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_629),
.B(n_654),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_688),
.A2(n_686),
.B(n_630),
.C(n_642),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_638),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_654),
.B(n_659),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_654),
.A2(n_660),
.B(n_656),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_619),
.A2(n_644),
.B(n_637),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_619),
.A2(n_644),
.B(n_637),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_660),
.A2(n_552),
.B(n_650),
.Y(n_871)
);

AND2x4_ASAP7_75t_SL g872 ( 
.A(n_713),
.B(n_504),
.Y(n_872)
);

NOR2xp67_ASAP7_75t_L g873 ( 
.A(n_657),
.B(n_492),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_619),
.B(n_606),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_606),
.B(n_418),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_635),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_606),
.B(n_418),
.Y(n_877)
);

CKINVDCx8_ASAP7_75t_R g878 ( 
.A(n_694),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_619),
.B(n_606),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_619),
.A2(n_627),
.B1(n_644),
.B2(n_612),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_670),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_754),
.A2(n_877),
.B(n_875),
.C(n_764),
.Y(n_882)
);

HB1xp67_ASAP7_75t_SL g883 ( 
.A(n_753),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_796),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_744),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_874),
.B(n_879),
.Y(n_886)
);

OAI21x1_ASAP7_75t_L g887 ( 
.A1(n_871),
.A2(n_748),
.B(n_760),
.Y(n_887)
);

BUFx12f_ASAP7_75t_L g888 ( 
.A(n_837),
.Y(n_888)
);

AO31x2_ASAP7_75t_L g889 ( 
.A1(n_769),
.A2(n_880),
.A3(n_747),
.B(n_757),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_801),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_808),
.A2(n_844),
.B1(n_765),
.B2(n_858),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_802),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_833),
.B(n_738),
.Y(n_893)
);

OAI21x1_ASAP7_75t_L g894 ( 
.A1(n_748),
.A2(n_871),
.B(n_864),
.Y(n_894)
);

AO31x2_ASAP7_75t_L g895 ( 
.A1(n_747),
.A2(n_749),
.A3(n_811),
.B(n_850),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_750),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_771),
.B(n_743),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_756),
.A2(n_742),
.B(n_758),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_793),
.Y(n_899)
);

AO31x2_ASAP7_75t_L g900 ( 
.A1(n_755),
.A2(n_762),
.A3(n_852),
.B(n_761),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_779),
.A2(n_782),
.B(n_746),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_843),
.B(n_857),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_774),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_763),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_787),
.A2(n_771),
.B(n_830),
.C(n_779),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_814),
.Y(n_906)
);

BUFx10_ASAP7_75t_L g907 ( 
.A(n_872),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_851),
.B(n_759),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_861),
.B(n_739),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_863),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_878),
.Y(n_911)
);

OAI21x1_ASAP7_75t_L g912 ( 
.A1(n_768),
.A2(n_862),
.B(n_766),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_784),
.A2(n_791),
.B1(n_786),
.B2(n_834),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_802),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_793),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_846),
.B(n_873),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_856),
.A2(n_768),
.B(n_862),
.Y(n_917)
);

NAND2x1p5_ASAP7_75t_L g918 ( 
.A(n_763),
.B(n_881),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_866),
.B(n_752),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_854),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_841),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_821),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_881),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_803),
.A2(n_827),
.B(n_845),
.C(n_838),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_817),
.B(n_805),
.Y(n_925)
);

AO21x2_ASAP7_75t_L g926 ( 
.A1(n_794),
.A2(n_778),
.B(n_755),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_785),
.B(n_788),
.Y(n_927)
);

AOI221xp5_ASAP7_75t_SL g928 ( 
.A1(n_838),
.A2(n_845),
.B1(n_847),
.B2(n_860),
.C(n_824),
.Y(n_928)
);

AOI21xp33_ASAP7_75t_L g929 ( 
.A1(n_780),
.A2(n_807),
.B(n_799),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_827),
.A2(n_842),
.B(n_847),
.C(n_835),
.Y(n_930)
);

AO31x2_ASAP7_75t_L g931 ( 
.A1(n_829),
.A2(n_849),
.A3(n_848),
.B(n_823),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_795),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_818),
.B(n_839),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_785),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_819),
.A2(n_809),
.B(n_772),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_806),
.A2(n_828),
.B(n_820),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_855),
.Y(n_937)
);

AOI21xp33_ASAP7_75t_L g938 ( 
.A1(n_780),
.A2(n_792),
.B(n_810),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_840),
.Y(n_939)
);

INVx6_ASAP7_75t_SL g940 ( 
.A(n_817),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_737),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_822),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_751),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_797),
.B(n_800),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_836),
.B(n_876),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_788),
.A2(n_831),
.B(n_826),
.Y(n_946)
);

AO31x2_ASAP7_75t_L g947 ( 
.A1(n_848),
.A2(n_867),
.A3(n_812),
.B(n_813),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_867),
.B(n_781),
.Y(n_948)
);

AOI21x1_ASAP7_75t_L g949 ( 
.A1(n_816),
.A2(n_825),
.B(n_773),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_836),
.B(n_876),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_789),
.A2(n_815),
.B1(n_826),
.B2(n_831),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_736),
.B(n_783),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_798),
.B(n_865),
.Y(n_953)
);

NOR2xp67_ASAP7_75t_L g954 ( 
.A(n_802),
.B(n_815),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_737),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_859),
.B(n_836),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_859),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_810),
.B(n_876),
.Y(n_958)
);

AO21x1_ASAP7_75t_L g959 ( 
.A1(n_790),
.A2(n_804),
.B(n_740),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_767),
.B(n_776),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_853),
.A2(n_767),
.B1(n_776),
.B2(n_777),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_776),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_832),
.A2(n_777),
.B(n_853),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_777),
.B(n_770),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_SL g965 ( 
.A1(n_754),
.A2(n_765),
.B(n_880),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_868),
.A2(n_760),
.B(n_748),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_868),
.A2(n_760),
.B(n_748),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_875),
.B(n_877),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_875),
.B(n_877),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_869),
.A2(n_619),
.B(n_870),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_875),
.B(n_877),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_875),
.B(n_877),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_875),
.B(n_877),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_763),
.B(n_881),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_837),
.Y(n_975)
);

NOR2x1_ASAP7_75t_SL g976 ( 
.A(n_763),
.B(n_881),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_875),
.B(n_877),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_875),
.B(n_613),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_868),
.A2(n_760),
.B(n_748),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_869),
.A2(n_619),
.B(n_870),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_869),
.A2(n_619),
.B(n_870),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_765),
.A2(n_718),
.B1(n_723),
.B2(n_701),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_869),
.A2(n_619),
.B(n_870),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_754),
.A2(n_879),
.B(n_874),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_754),
.A2(n_879),
.B(n_874),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_SL g986 ( 
.A(n_753),
.B(n_557),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_868),
.A2(n_760),
.B(n_748),
.Y(n_987)
);

AO31x2_ASAP7_75t_L g988 ( 
.A1(n_754),
.A2(n_741),
.A3(n_745),
.B(n_769),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_874),
.A2(n_879),
.B1(n_754),
.B2(n_619),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_869),
.A2(n_619),
.B(n_870),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_868),
.A2(n_871),
.B(n_748),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_875),
.B(n_877),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_802),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_868),
.A2(n_871),
.B(n_748),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_754),
.A2(n_879),
.B(n_874),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_754),
.A2(n_879),
.B(n_874),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_875),
.B(n_877),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_869),
.A2(n_619),
.B(n_870),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_875),
.B(n_877),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_875),
.B(n_877),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_869),
.A2(n_619),
.B(n_870),
.Y(n_1001)
);

AOI21x1_ASAP7_75t_SL g1002 ( 
.A1(n_874),
.A2(n_879),
.B(n_648),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_753),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_754),
.B(n_880),
.Y(n_1004)
);

BUFx4_ASAP7_75t_SL g1005 ( 
.A(n_841),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_875),
.B(n_613),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_875),
.B(n_877),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_869),
.A2(n_619),
.B(n_870),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_875),
.B(n_877),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_802),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_875),
.B(n_877),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_868),
.A2(n_871),
.B(n_748),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_868),
.A2(n_871),
.B(n_748),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_868),
.A2(n_871),
.B(n_748),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_775),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_744),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_875),
.B(n_877),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_868),
.A2(n_871),
.B(n_748),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_978),
.B(n_1006),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_992),
.A2(n_999),
.B1(n_1017),
.B2(n_1011),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_884),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_992),
.B(n_999),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_974),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_989),
.A2(n_980),
.B(n_970),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_1017),
.A2(n_882),
.B1(n_982),
.B2(n_972),
.Y(n_1025)
);

INVx8_ASAP7_75t_L g1026 ( 
.A(n_888),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_968),
.B(n_969),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_981),
.A2(n_990),
.B(n_983),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_971),
.B(n_973),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_977),
.B(n_997),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_1003),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1000),
.B(n_1007),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_998),
.A2(n_1008),
.B(n_1001),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1009),
.B(n_886),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_884),
.Y(n_1035)
);

CKINVDCx8_ASAP7_75t_R g1036 ( 
.A(n_932),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_920),
.Y(n_1037)
);

INVx4_ASAP7_75t_SL g1038 ( 
.A(n_888),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_907),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_909),
.B(n_908),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_893),
.B(n_909),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_882),
.B(n_891),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_982),
.A2(n_924),
.B1(n_965),
.B2(n_905),
.Y(n_1043)
);

AOI21xp33_ASAP7_75t_SL g1044 ( 
.A1(n_911),
.A2(n_932),
.B(n_975),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_SL g1045 ( 
.A(n_953),
.B(n_945),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_974),
.B(n_892),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_938),
.A2(n_943),
.B1(n_929),
.B2(n_940),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_924),
.A2(n_928),
.B1(n_995),
.B2(n_996),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_974),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_919),
.B(n_902),
.Y(n_1050)
);

INVx3_ASAP7_75t_SL g1051 ( 
.A(n_883),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_899),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_905),
.A2(n_901),
.B(n_898),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_913),
.A2(n_1004),
.B1(n_944),
.B2(n_930),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_885),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_925),
.B(n_915),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1004),
.A2(n_930),
.B1(n_897),
.B2(n_933),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_903),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_954),
.B(n_921),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_916),
.B(n_943),
.Y(n_1060)
);

BUFx12f_ASAP7_75t_L g1061 ( 
.A(n_911),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_986),
.A2(n_936),
.B(n_948),
.C(n_952),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_957),
.B(n_914),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_SL g1064 ( 
.A(n_907),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_918),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_SL g1066 ( 
.A(n_904),
.B(n_923),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_940),
.A2(n_939),
.B1(n_922),
.B2(n_906),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_1003),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_914),
.B(n_993),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_894),
.A2(n_887),
.B(n_1018),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_1005),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_910),
.B(n_1016),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_937),
.B(n_907),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_914),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_SL g1075 ( 
.A1(n_926),
.A2(n_942),
.B1(n_958),
.B2(n_940),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_960),
.B(n_942),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_918),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_993),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_991),
.A2(n_1018),
.B(n_1014),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_1005),
.Y(n_1080)
);

NAND2x1_ASAP7_75t_L g1081 ( 
.A(n_927),
.B(n_923),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_890),
.B(n_1015),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_904),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_993),
.B(n_1010),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_1010),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_941),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_941),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_955),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_927),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_956),
.B(n_1010),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_976),
.B(n_927),
.Y(n_1091)
);

BUFx4f_ASAP7_75t_L g1092 ( 
.A(n_934),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_962),
.B(n_961),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_945),
.B(n_950),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_964),
.A2(n_951),
.B(n_926),
.C(n_963),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_946),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_950),
.B(n_900),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_964),
.A2(n_959),
.B(n_1002),
.C(n_895),
.Y(n_1098)
);

CKINVDCx14_ASAP7_75t_R g1099 ( 
.A(n_947),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_994),
.A2(n_1013),
.B(n_1012),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_900),
.B(n_988),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_988),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_917),
.A2(n_912),
.B1(n_935),
.B2(n_987),
.Y(n_1103)
);

NAND2xp33_ASAP7_75t_L g1104 ( 
.A(n_947),
.B(n_949),
.Y(n_1104)
);

INVx5_ASAP7_75t_L g1105 ( 
.A(n_900),
.Y(n_1105)
);

OAI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_966),
.A2(n_967),
.B(n_979),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_947),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_988),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_947),
.B(n_895),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_889),
.B(n_895),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_889),
.B(n_895),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_931),
.B(n_889),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_889),
.A2(n_992),
.B1(n_1017),
.B2(n_999),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_992),
.A2(n_999),
.B1(n_1017),
.B2(n_882),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_968),
.B(n_969),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_SL g1116 ( 
.A1(n_984),
.A2(n_995),
.B(n_985),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_974),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_978),
.B(n_1006),
.Y(n_1118)
);

CKINVDCx8_ASAP7_75t_R g1119 ( 
.A(n_932),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_974),
.Y(n_1120)
);

NOR2xp67_ASAP7_75t_L g1121 ( 
.A(n_961),
.B(n_621),
.Y(n_1121)
);

OR2x6_ASAP7_75t_L g1122 ( 
.A(n_965),
.B(n_670),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1003),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_920),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_992),
.B(n_1017),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_883),
.Y(n_1126)
);

BUFx2_ASAP7_75t_SL g1127 ( 
.A(n_1003),
.Y(n_1127)
);

OR2x6_ASAP7_75t_L g1128 ( 
.A(n_965),
.B(n_670),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_920),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_992),
.A2(n_1017),
.B(n_999),
.C(n_875),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_885),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_992),
.B(n_1017),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_SL g1133 ( 
.A1(n_992),
.A2(n_606),
.B(n_1017),
.C(n_999),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_992),
.B(n_1017),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_885),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_974),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_914),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_989),
.A2(n_754),
.B(n_869),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_992),
.B(n_1017),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_974),
.B(n_892),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_989),
.A2(n_754),
.B(n_869),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_SL g1142 ( 
.A1(n_992),
.A2(n_999),
.B1(n_1017),
.B2(n_452),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_974),
.Y(n_1143)
);

O2A1O1Ixp5_ASAP7_75t_L g1144 ( 
.A1(n_992),
.A2(n_999),
.B(n_1017),
.C(n_875),
.Y(n_1144)
);

AOI222xp33_ASAP7_75t_L g1145 ( 
.A1(n_992),
.A2(n_999),
.B1(n_1017),
.B2(n_982),
.C1(n_1009),
.C2(n_1011),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_989),
.A2(n_754),
.B(n_869),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_884),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_974),
.B(n_892),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_896),
.Y(n_1149)
);

BUFx12f_ASAP7_75t_L g1150 ( 
.A(n_911),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_978),
.B(n_1006),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_896),
.Y(n_1152)
);

NOR2x1_ASAP7_75t_SL g1153 ( 
.A(n_953),
.B(n_945),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_896),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1145),
.A2(n_1142),
.B1(n_1025),
.B2(n_1114),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_SL g1156 ( 
.A(n_1031),
.Y(n_1156)
);

CKINVDCx11_ASAP7_75t_R g1157 ( 
.A(n_1080),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1055),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1058),
.Y(n_1159)
);

AOI222xp33_ASAP7_75t_L g1160 ( 
.A1(n_1025),
.A2(n_1043),
.B1(n_1139),
.B2(n_1125),
.C1(n_1134),
.C2(n_1022),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1023),
.B(n_1049),
.Y(n_1161)
);

AO21x1_ASAP7_75t_L g1162 ( 
.A1(n_1043),
.A2(n_1113),
.B(n_1114),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1145),
.A2(n_1113),
.B1(n_1020),
.B2(n_1042),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1046),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_SL g1165 ( 
.A1(n_1107),
.A2(n_1099),
.B1(n_1132),
.B2(n_1057),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1019),
.B(n_1118),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_1068),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1085),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1097),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_SL g1170 ( 
.A1(n_1057),
.A2(n_1116),
.B1(n_1041),
.B2(n_1153),
.Y(n_1170)
);

INVx6_ASAP7_75t_L g1171 ( 
.A(n_1039),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_1037),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1124),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_SL g1174 ( 
.A1(n_1045),
.A2(n_1040),
.B1(n_1105),
.B2(n_1027),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1140),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1102),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1020),
.A2(n_1054),
.B1(n_1151),
.B2(n_1047),
.Y(n_1177)
);

BUFx4f_ASAP7_75t_SL g1178 ( 
.A(n_1061),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1130),
.A2(n_1054),
.B1(n_1048),
.B2(n_1115),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1060),
.B(n_1056),
.Y(n_1180)
);

INVx6_ASAP7_75t_L g1181 ( 
.A(n_1039),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1029),
.B(n_1144),
.Y(n_1182)
);

BUFx2_ASAP7_75t_R g1183 ( 
.A(n_1071),
.Y(n_1183)
);

INVx6_ASAP7_75t_L g1184 ( 
.A(n_1039),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1048),
.A2(n_1034),
.B1(n_1030),
.B2(n_1032),
.Y(n_1185)
);

OAI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1122),
.A2(n_1128),
.B1(n_1050),
.B2(n_1146),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1149),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1131),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1108),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1135),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1140),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1082),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1087),
.Y(n_1193)
);

OAI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1122),
.A2(n_1128),
.B1(n_1138),
.B2(n_1141),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1086),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1075),
.A2(n_1110),
.B1(n_1072),
.B2(n_1101),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1129),
.B(n_1023),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1088),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_SL g1199 ( 
.A1(n_1105),
.A2(n_1110),
.B1(n_1122),
.B2(n_1128),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_SL g1200 ( 
.A1(n_1105),
.A2(n_1154),
.B1(n_1152),
.B2(n_1149),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1076),
.A2(n_1067),
.B1(n_1111),
.B2(n_1147),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1035),
.A2(n_1053),
.B1(n_1152),
.B2(n_1154),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1133),
.B(n_1021),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1127),
.B(n_1052),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1073),
.A2(n_1148),
.B1(n_1126),
.B2(n_1059),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1049),
.B(n_1117),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1074),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1094),
.Y(n_1208)
);

AOI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1079),
.A2(n_1100),
.B(n_1121),
.Y(n_1209)
);

INVx6_ASAP7_75t_L g1210 ( 
.A(n_1150),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1112),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_R g1212 ( 
.A1(n_1036),
.A2(n_1119),
.B1(n_1123),
.B2(n_1038),
.Y(n_1212)
);

INVxp67_ASAP7_75t_SL g1213 ( 
.A(n_1104),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1090),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1026),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_SL g1216 ( 
.A1(n_1053),
.A2(n_1093),
.B1(n_1059),
.B2(n_1064),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1026),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1064),
.A2(n_1143),
.B1(n_1136),
.B2(n_1120),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1084),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1026),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1038),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_1063),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1109),
.A2(n_1143),
.B1(n_1136),
.B2(n_1120),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1063),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_R g1225 ( 
.A(n_1117),
.B(n_1092),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1078),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1089),
.B(n_1092),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1062),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1078),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1089),
.A2(n_1091),
.B1(n_1065),
.B2(n_1077),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1070),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1121),
.A2(n_1091),
.B1(n_1065),
.B2(n_1077),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1078),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1083),
.B(n_1066),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1069),
.Y(n_1235)
);

AOI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1070),
.A2(n_1081),
.B(n_1069),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1069),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1137),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_1137),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1137),
.Y(n_1240)
);

BUFx12f_ASAP7_75t_L g1241 ( 
.A(n_1044),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1083),
.Y(n_1242)
);

INVx8_ASAP7_75t_L g1243 ( 
.A(n_1096),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1098),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1103),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1106),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1095),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1097),
.Y(n_1248)
);

NAND2x1p5_ASAP7_75t_L g1249 ( 
.A(n_1023),
.B(n_1049),
.Y(n_1249)
);

CKINVDCx6p67_ASAP7_75t_R g1250 ( 
.A(n_1051),
.Y(n_1250)
);

AOI222xp33_ASAP7_75t_L g1251 ( 
.A1(n_1025),
.A2(n_999),
.B1(n_992),
.B2(n_1017),
.C1(n_982),
.C2(n_997),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1023),
.B(n_1049),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1026),
.Y(n_1253)
);

BUFx2_ASAP7_75t_SL g1254 ( 
.A(n_1080),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1130),
.A2(n_1020),
.B1(n_999),
.B2(n_1017),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1055),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1055),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1019),
.B(n_1118),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1097),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1074),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1026),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1130),
.A2(n_1020),
.B1(n_999),
.B2(n_1017),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1028),
.A2(n_1033),
.B(n_1024),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1074),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1055),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_1122),
.B(n_1128),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1085),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1041),
.B(n_1035),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1025),
.A2(n_992),
.B1(n_1017),
.B2(n_999),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1055),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1157),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1169),
.B(n_1248),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1236),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1168),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1158),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1176),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1176),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1162),
.A2(n_1245),
.A3(n_1247),
.B(n_1246),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1166),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1193),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1243),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1243),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1259),
.B(n_1182),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1259),
.B(n_1231),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1208),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1189),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1157),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1213),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1270),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1209),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1231),
.B(n_1180),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1159),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1268),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1213),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1168),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1188),
.Y(n_1296)
);

AOI21xp33_ASAP7_75t_L g1297 ( 
.A1(n_1251),
.A2(n_1228),
.B(n_1155),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1185),
.B(n_1160),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1266),
.A2(n_1179),
.B(n_1186),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1190),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1256),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1185),
.B(n_1269),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1257),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1219),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1265),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1163),
.B(n_1155),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1244),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1195),
.B(n_1202),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1202),
.B(n_1163),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1211),
.A2(n_1196),
.B(n_1203),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1224),
.B(n_1175),
.Y(n_1311)
);

NAND2x1_ASAP7_75t_L g1312 ( 
.A(n_1171),
.B(n_1181),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1220),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1258),
.B(n_1165),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1192),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1255),
.B(n_1262),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1242),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1214),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1198),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1221),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1242),
.Y(n_1321)
);

AO21x2_ASAP7_75t_L g1322 ( 
.A1(n_1186),
.A2(n_1194),
.B(n_1218),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1263),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1196),
.A2(n_1201),
.B1(n_1177),
.B2(n_1174),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1263),
.A2(n_1232),
.B(n_1249),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1194),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1232),
.A2(n_1249),
.B(n_1234),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1199),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1229),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1233),
.Y(n_1330)
);

OAI21xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1177),
.A2(n_1239),
.B(n_1197),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1238),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1240),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1170),
.B(n_1252),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1223),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1161),
.B(n_1206),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1161),
.Y(n_1337)
);

OAI221xp5_ASAP7_75t_L g1338 ( 
.A1(n_1205),
.A2(n_1216),
.B1(n_1167),
.B2(n_1187),
.C(n_1201),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1161),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1206),
.Y(n_1340)
);

AND2x6_ASAP7_75t_L g1341 ( 
.A(n_1206),
.B(n_1252),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1235),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_SL g1343 ( 
.A1(n_1227),
.A2(n_1225),
.B(n_1164),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1197),
.B(n_1173),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1172),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1200),
.A2(n_1222),
.B1(n_1156),
.B2(n_1230),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1204),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1237),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1280),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1280),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1307),
.B(n_1264),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1283),
.B(n_1267),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1283),
.B(n_1226),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_1307),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1291),
.B(n_1226),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1306),
.A2(n_1156),
.B1(n_1210),
.B2(n_1212),
.Y(n_1356)
);

OAI222xp33_ASAP7_75t_L g1357 ( 
.A1(n_1309),
.A2(n_1227),
.B1(n_1221),
.B2(n_1220),
.C1(n_1178),
.C2(n_1215),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1289),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1291),
.B(n_1207),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1289),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1284),
.B(n_1260),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1292),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1284),
.B(n_1164),
.Y(n_1363)
);

INVxp67_ASAP7_75t_SL g1364 ( 
.A(n_1323),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_SL g1365 ( 
.A1(n_1316),
.A2(n_1261),
.B(n_1253),
.Y(n_1365)
);

AOI33xp33_ASAP7_75t_L g1366 ( 
.A1(n_1306),
.A2(n_1241),
.A3(n_1250),
.B1(n_1254),
.B2(n_1178),
.B3(n_1183),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1276),
.Y(n_1367)
);

OR2x6_ASAP7_75t_L g1368 ( 
.A(n_1299),
.B(n_1325),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1276),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1285),
.B(n_1184),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1285),
.B(n_1184),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1297),
.A2(n_1298),
.B1(n_1302),
.B2(n_1309),
.Y(n_1372)
);

INVx5_ASAP7_75t_L g1373 ( 
.A(n_1341),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1277),
.B(n_1272),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1288),
.B(n_1191),
.Y(n_1375)
);

AND2x4_ASAP7_75t_SL g1376 ( 
.A(n_1311),
.B(n_1225),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1317),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1293),
.B(n_1308),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1296),
.B(n_1210),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1303),
.B(n_1210),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1312),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1303),
.B(n_1217),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1305),
.B(n_1217),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1308),
.B(n_1241),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1315),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1271),
.B(n_1287),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1344),
.B(n_1337),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1344),
.B(n_1339),
.Y(n_1388)
);

AOI211xp5_ASAP7_75t_L g1389 ( 
.A1(n_1338),
.A2(n_1331),
.B(n_1335),
.C(n_1334),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1317),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1278),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1318),
.B(n_1278),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1378),
.B(n_1347),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1369),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1386),
.B(n_1271),
.Y(n_1395)
);

AOI221xp5_ASAP7_75t_L g1396 ( 
.A1(n_1372),
.A2(n_1314),
.B1(n_1301),
.B2(n_1300),
.C(n_1275),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1372),
.A2(n_1324),
.B1(n_1328),
.B2(n_1335),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1389),
.B(n_1329),
.C(n_1330),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1387),
.B(n_1288),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1389),
.A2(n_1326),
.B1(n_1279),
.B2(n_1314),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1356),
.A2(n_1334),
.B1(n_1294),
.B2(n_1345),
.Y(n_1401)
);

OAI221xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1356),
.A2(n_1346),
.B1(n_1328),
.B2(n_1294),
.C(n_1304),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1365),
.A2(n_1313),
.B1(n_1295),
.B2(n_1274),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1387),
.B(n_1339),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1378),
.B(n_1354),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1354),
.B(n_1321),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1374),
.B(n_1321),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1365),
.A2(n_1295),
.B1(n_1274),
.B2(n_1287),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1374),
.B(n_1329),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1367),
.B(n_1330),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1388),
.B(n_1361),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1361),
.B(n_1340),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1367),
.B(n_1333),
.Y(n_1413)
);

NAND4xp25_ASAP7_75t_L g1414 ( 
.A(n_1382),
.B(n_1383),
.C(n_1366),
.D(n_1351),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1352),
.B(n_1333),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1357),
.A2(n_1282),
.B(n_1281),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1361),
.B(n_1336),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1352),
.B(n_1278),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1363),
.B(n_1336),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_L g1420 ( 
.A(n_1391),
.B(n_1332),
.C(n_1342),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1355),
.B(n_1278),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1384),
.A2(n_1310),
.B1(n_1391),
.B2(n_1322),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1363),
.B(n_1278),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1355),
.B(n_1332),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1359),
.B(n_1310),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1353),
.B(n_1310),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1353),
.B(n_1310),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1359),
.B(n_1286),
.Y(n_1428)
);

OAI221xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1368),
.A2(n_1348),
.B1(n_1342),
.B2(n_1273),
.C(n_1323),
.Y(n_1429)
);

NOR3xp33_ASAP7_75t_L g1430 ( 
.A(n_1357),
.B(n_1351),
.C(n_1370),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1368),
.A2(n_1343),
.B(n_1312),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1376),
.A2(n_1383),
.B(n_1382),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1373),
.B(n_1273),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1369),
.B(n_1286),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_1392),
.B(n_1348),
.C(n_1319),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1375),
.B(n_1290),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1381),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1385),
.B(n_1327),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1392),
.B(n_1370),
.C(n_1371),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1394),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1433),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1438),
.Y(n_1442)
);

INVxp67_ASAP7_75t_SL g1443 ( 
.A(n_1435),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1426),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1434),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1426),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1427),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1418),
.B(n_1364),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1423),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1425),
.B(n_1364),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1423),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1439),
.B(n_1385),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1405),
.B(n_1377),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1421),
.B(n_1390),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1439),
.B(n_1390),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1393),
.B(n_1349),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1433),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1411),
.B(n_1417),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1412),
.B(n_1404),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1407),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1410),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1409),
.B(n_1413),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1435),
.B(n_1350),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1433),
.B(n_1373),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1406),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1428),
.B(n_1350),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1433),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1430),
.B(n_1358),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1399),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1437),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1420),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1437),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1420),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1458),
.B(n_1419),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1458),
.B(n_1419),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1458),
.B(n_1459),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1458),
.B(n_1436),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1459),
.B(n_1436),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1444),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1464),
.B(n_1441),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1459),
.B(n_1432),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_L g1482 ( 
.A(n_1455),
.B(n_1414),
.C(n_1408),
.D(n_1403),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1459),
.B(n_1432),
.Y(n_1483)
);

NAND4xp25_ASAP7_75t_L g1484 ( 
.A(n_1455),
.B(n_1414),
.C(n_1398),
.D(n_1416),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1463),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1443),
.Y(n_1486)
);

OR2x6_ASAP7_75t_L g1487 ( 
.A(n_1464),
.B(n_1431),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1460),
.B(n_1415),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1463),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1456),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1444),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1468),
.B(n_1424),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1468),
.B(n_1398),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1460),
.B(n_1396),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1456),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1444),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1462),
.B(n_1416),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1469),
.B(n_1379),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1456),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1470),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1443),
.B(n_1360),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1469),
.B(n_1379),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1464),
.B(n_1373),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1466),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1471),
.A2(n_1400),
.B(n_1401),
.Y(n_1505)
);

NOR2x1_ASAP7_75t_SL g1506 ( 
.A(n_1470),
.B(n_1373),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1466),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1470),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1471),
.A2(n_1400),
.B1(n_1402),
.B2(n_1401),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1462),
.B(n_1429),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1461),
.B(n_1362),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1453),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1462),
.B(n_1362),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1509),
.A2(n_1397),
.B1(n_1473),
.B2(n_1471),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1493),
.Y(n_1515)
);

NAND2x1_ASAP7_75t_L g1516 ( 
.A(n_1480),
.B(n_1441),
.Y(n_1516)
);

NAND4xp25_ASAP7_75t_L g1517 ( 
.A(n_1486),
.B(n_1455),
.C(n_1473),
.D(n_1395),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1493),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1486),
.B(n_1473),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1485),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1481),
.B(n_1483),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1513),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1513),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1476),
.B(n_1441),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1511),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1492),
.B(n_1461),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1481),
.B(n_1441),
.Y(n_1527)
);

OAI211xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1505),
.A2(n_1440),
.B(n_1445),
.C(n_1452),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1479),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1492),
.B(n_1484),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1512),
.B(n_1461),
.Y(n_1531)
);

AND3x2_ASAP7_75t_L g1532 ( 
.A(n_1494),
.B(n_1447),
.C(n_1449),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1483),
.B(n_1476),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1474),
.B(n_1475),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1500),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1490),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1474),
.B(n_1447),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1490),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1495),
.B(n_1452),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1475),
.B(n_1457),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1480),
.B(n_1457),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1485),
.B(n_1465),
.Y(n_1542)
);

NAND2x1_ASAP7_75t_L g1543 ( 
.A(n_1480),
.B(n_1472),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1495),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1499),
.B(n_1448),
.Y(n_1545)
);

NAND2x1p5_ASAP7_75t_L g1546 ( 
.A(n_1500),
.B(n_1373),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1508),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1499),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1482),
.A2(n_1422),
.B1(n_1449),
.B2(n_1451),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1480),
.B(n_1477),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1504),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1479),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1491),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1489),
.B(n_1488),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1504),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1507),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1491),
.Y(n_1557)
);

INVxp33_ASAP7_75t_L g1558 ( 
.A(n_1521),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1535),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1521),
.B(n_1508),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1514),
.B(n_1489),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1530),
.B(n_1507),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1533),
.B(n_1477),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1535),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1544),
.Y(n_1565)
);

INVxp33_ASAP7_75t_L g1566 ( 
.A(n_1517),
.Y(n_1566)
);

AO21x2_ASAP7_75t_L g1567 ( 
.A1(n_1519),
.A2(n_1501),
.B(n_1510),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1547),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1544),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1548),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1532),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1529),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1548),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1530),
.B(n_1510),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1533),
.B(n_1478),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1527),
.B(n_1478),
.Y(n_1576)
);

BUFx4f_ASAP7_75t_SL g1577 ( 
.A(n_1527),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1534),
.B(n_1497),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1515),
.B(n_1497),
.Y(n_1579)
);

AO21x1_ASAP7_75t_L g1580 ( 
.A1(n_1549),
.A2(n_1496),
.B(n_1450),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1516),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1534),
.B(n_1498),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1516),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1518),
.B(n_1465),
.Y(n_1584)
);

NOR2xp67_ASAP7_75t_SL g1585 ( 
.A(n_1520),
.B(n_1320),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1536),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1538),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1528),
.A2(n_1448),
.B(n_1450),
.Y(n_1588)
);

CKINVDCx16_ASAP7_75t_R g1589 ( 
.A(n_1550),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1551),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1526),
.B(n_1320),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1555),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1550),
.B(n_1498),
.Y(n_1593)
);

NAND2xp33_ASAP7_75t_SL g1594 ( 
.A(n_1566),
.B(n_1543),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1565),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1558),
.B(n_1559),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1571),
.A2(n_1524),
.B1(n_1543),
.B2(n_1537),
.Y(n_1597)
);

NAND2x1_ASAP7_75t_L g1598 ( 
.A(n_1581),
.B(n_1524),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1561),
.A2(n_1542),
.B(n_1539),
.C(n_1554),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1574),
.A2(n_1557),
.B1(n_1529),
.B2(n_1553),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1574),
.B(n_1531),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1565),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1571),
.B(n_1524),
.Y(n_1603)
);

AOI21xp33_ASAP7_75t_L g1604 ( 
.A1(n_1571),
.A2(n_1539),
.B(n_1556),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1569),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1589),
.B(n_1537),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1589),
.B(n_1541),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1577),
.Y(n_1608)
);

NAND2x1_ASAP7_75t_L g1609 ( 
.A(n_1581),
.B(n_1541),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1578),
.B(n_1540),
.Y(n_1610)
);

AOI211xp5_ASAP7_75t_L g1611 ( 
.A1(n_1571),
.A2(n_1545),
.B(n_1522),
.C(n_1523),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1569),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1559),
.B(n_1525),
.Y(n_1613)
);

INVxp67_ASAP7_75t_SL g1614 ( 
.A(n_1571),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1579),
.B(n_1545),
.Y(n_1615)
);

NAND2xp33_ASAP7_75t_SL g1616 ( 
.A(n_1571),
.B(n_1540),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1561),
.A2(n_1506),
.B(n_1487),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1578),
.B(n_1502),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1564),
.B(n_1454),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1608),
.B(n_1564),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1595),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1616),
.A2(n_1580),
.B1(n_1567),
.B2(n_1600),
.Y(n_1622)
);

NOR2xp67_ASAP7_75t_L g1623 ( 
.A(n_1603),
.B(n_1581),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1602),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1610),
.B(n_1568),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1596),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1605),
.Y(n_1627)
);

AOI21xp33_ASAP7_75t_L g1628 ( 
.A1(n_1614),
.A2(n_1567),
.B(n_1562),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1606),
.B(n_1560),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1607),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1619),
.B(n_1560),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1619),
.B(n_1568),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1603),
.B(n_1564),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1616),
.A2(n_1580),
.B1(n_1567),
.B2(n_1600),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1601),
.B(n_1591),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1613),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1594),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1612),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1615),
.B(n_1579),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1622),
.A2(n_1567),
.B1(n_1611),
.B2(n_1604),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1629),
.B(n_1593),
.Y(n_1641)
);

O2A1O1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1628),
.A2(n_1599),
.B(n_1562),
.C(n_1597),
.Y(n_1642)
);

OAI21xp33_ASAP7_75t_L g1643 ( 
.A1(n_1620),
.A2(n_1634),
.B(n_1629),
.Y(n_1643)
);

AOI211xp5_ASAP7_75t_L g1644 ( 
.A1(n_1637),
.A2(n_1594),
.B(n_1617),
.C(n_1585),
.Y(n_1644)
);

OAI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1639),
.A2(n_1588),
.B1(n_1609),
.B2(n_1598),
.C(n_1584),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1633),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1631),
.B(n_1630),
.Y(n_1647)
);

AOI21xp33_ASAP7_75t_L g1648 ( 
.A1(n_1636),
.A2(n_1572),
.B(n_1570),
.Y(n_1648)
);

NOR3x1_ASAP7_75t_L g1649 ( 
.A(n_1625),
.B(n_1583),
.C(n_1618),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1623),
.B(n_1632),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1623),
.A2(n_1592),
.B(n_1583),
.Y(n_1651)
);

NAND5xp2_ASAP7_75t_L g1652 ( 
.A(n_1644),
.B(n_1631),
.C(n_1635),
.D(n_1621),
.E(n_1624),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1642),
.A2(n_1626),
.B(n_1630),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1643),
.B(n_1624),
.C(n_1621),
.Y(n_1654)
);

NOR2x1_ASAP7_75t_L g1655 ( 
.A(n_1650),
.B(n_1627),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1641),
.Y(n_1656)
);

NAND4xp75_ASAP7_75t_L g1657 ( 
.A(n_1649),
.B(n_1638),
.C(n_1627),
.D(n_1572),
.Y(n_1657)
);

NOR2x1_ASAP7_75t_L g1658 ( 
.A(n_1647),
.B(n_1638),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1646),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1640),
.A2(n_1573),
.B1(n_1570),
.B2(n_1588),
.C(n_1587),
.Y(n_1660)
);

AOI211xp5_ASAP7_75t_L g1661 ( 
.A1(n_1645),
.A2(n_1585),
.B(n_1573),
.C(n_1587),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1648),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1656),
.B(n_1651),
.Y(n_1663)
);

AOI21xp33_ASAP7_75t_L g1664 ( 
.A1(n_1658),
.A2(n_1572),
.B(n_1586),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1655),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1652),
.B(n_1581),
.Y(n_1666)
);

NOR4xp25_ASAP7_75t_L g1667 ( 
.A(n_1662),
.B(n_1590),
.C(n_1586),
.D(n_1575),
.Y(n_1667)
);

OAI211xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1653),
.A2(n_1660),
.B(n_1661),
.C(n_1654),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1659),
.B(n_1582),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1657),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1669),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1665),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1664),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1663),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1667),
.B(n_1576),
.Y(n_1675)
);

INVxp67_ASAP7_75t_SL g1676 ( 
.A(n_1670),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1666),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1668),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1677),
.B(n_1590),
.Y(n_1679)
);

OAI211xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1678),
.A2(n_1472),
.B(n_1467),
.C(n_1457),
.Y(n_1680)
);

AND3x4_ASAP7_75t_L g1681 ( 
.A(n_1671),
.B(n_1470),
.C(n_1503),
.Y(n_1681)
);

AND3x4_ASAP7_75t_L g1682 ( 
.A(n_1675),
.B(n_1503),
.C(n_1464),
.Y(n_1682)
);

NOR2x1_ASAP7_75t_L g1683 ( 
.A(n_1674),
.B(n_1673),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1672),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1681),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1684),
.Y(n_1686)
);

OAI22x1_ASAP7_75t_L g1687 ( 
.A1(n_1683),
.A2(n_1676),
.B1(n_1673),
.B2(n_1672),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1687),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1688),
.B(n_1686),
.C(n_1676),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1689),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1689),
.A2(n_1679),
.B(n_1685),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1690),
.Y(n_1692)
);

AOI21xp33_ASAP7_75t_SL g1693 ( 
.A1(n_1691),
.A2(n_1682),
.B(n_1680),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1692),
.B1(n_1552),
.B2(n_1557),
.C(n_1553),
.Y(n_1694)
);

OA21x2_ASAP7_75t_L g1695 ( 
.A1(n_1692),
.A2(n_1575),
.B(n_1563),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1695),
.B(n_1563),
.Y(n_1696)
);

AOI322xp5_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1694),
.A3(n_1552),
.B1(n_1576),
.B2(n_1593),
.C1(n_1582),
.C2(n_1496),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1697),
.A2(n_1546),
.B1(n_1442),
.B2(n_1444),
.C(n_1446),
.Y(n_1698)
);

AOI211xp5_ASAP7_75t_L g1699 ( 
.A1(n_1698),
.A2(n_1380),
.B(n_1503),
.C(n_1467),
.Y(n_1699)
);


endmodule