module real_jpeg_16934_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_556;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_SL g36 ( 
.A(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_0),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_0),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_0),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_0),
.B(n_164),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_20),
.B(n_560),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_1),
.B(n_561),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_2),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_2),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_2),
.B(n_152),
.Y(n_151)
);

NAND2x1_ASAP7_75t_L g220 ( 
.A(n_2),
.B(n_70),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_2),
.B(n_267),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_2),
.B(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_2),
.B(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_3),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g294 ( 
.A(n_3),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g359 ( 
.A(n_3),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_5),
.Y(n_270)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_5),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_5),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_5),
.Y(n_494)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_6),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_6),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_6),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_6),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_6),
.B(n_368),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_6),
.B(n_267),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_6),
.B(n_261),
.Y(n_475)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_7),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_7),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_7),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_8),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_8),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_8),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_8),
.B(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_8),
.B(n_503),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_8),
.B(n_512),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_8),
.B(n_520),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_9),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_9),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_9),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_9),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_9),
.B(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_9),
.B(n_293),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_9),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_9),
.B(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_10),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_10),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_10),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_10),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_10),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_10),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_10),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_11),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_11),
.B(n_245),
.Y(n_244)
);

AOI22x1_ASAP7_75t_L g290 ( 
.A1(n_11),
.A2(n_15),
.B1(n_291),
.B2(n_295),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_11),
.B(n_362),
.Y(n_361)
);

AOI31xp67_ASAP7_75t_L g404 ( 
.A1(n_11),
.A2(n_290),
.A3(n_405),
.B(n_408),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_11),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_11),
.B(n_462),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_11),
.B(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_11),
.B(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_12),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_13),
.Y(n_149)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_13),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_14),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_14),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_14),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_14),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_14),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_14),
.B(n_312),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_14),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_14),
.B(n_294),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_15),
.B(n_47),
.Y(n_46)
);

NAND2x1_ASAP7_75t_L g64 ( 
.A(n_15),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_15),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_15),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_15),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_15),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_15),
.B(n_269),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_15),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_16),
.Y(n_251)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_16),
.Y(n_375)
);

BUFx5_ASAP7_75t_L g440 ( 
.A(n_16),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_17),
.Y(n_139)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_18),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_18),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_18),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_182),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_180),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_155),
.Y(n_22)
);

NOR2xp67_ASAP7_75t_R g181 ( 
.A(n_23),
.B(n_155),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_113),
.C(n_128),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_24),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_72),
.C(n_93),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_26),
.B(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_45),
.C(n_58),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_27),
.B(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_28),
.B(n_35),
.C(n_41),
.Y(n_126)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_30),
.Y(n_437)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_32),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_32),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_34),
.A2(n_35),
.B1(n_116),
.B2(n_119),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_35),
.B(n_116),
.C(n_120),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_40),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_41),
.A2(n_42),
.B1(n_96),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_42),
.B(n_96),
.C(n_99),
.Y(n_95)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_43),
.Y(n_474)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_44),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_45),
.B(n_58),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.C(n_54),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_46),
.B(n_54),
.Y(n_214)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_50),
.B(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_59),
.B(n_64),
.C(n_69),
.Y(n_127)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_62),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_73),
.B(n_93),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_84),
.C(n_92),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_91),
.B2(n_92),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_83),
.Y(n_273)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_87),
.Y(n_301)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_89),
.Y(n_254)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_89),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.C(n_109),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_94),
.A2(n_95),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_96),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_96),
.B(n_204),
.C(n_208),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_96),
.A2(n_202),
.B1(n_209),
.B2(n_257),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_97),
.Y(n_411)
);

INVx6_ASAP7_75t_L g508 ( 
.A(n_97),
.Y(n_508)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_98),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_99),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_99),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_99),
.A2(n_199),
.B1(n_302),
.B2(n_351),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_102),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_102),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_103),
.B(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_104),
.B(n_109),
.Y(n_229)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_105),
.B(n_260),
.C(n_264),
.Y(n_259)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_109),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_SL g276 ( 
.A(n_109),
.B(n_224),
.Y(n_276)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_113),
.A2(n_128),
.B1(n_129),
.B2(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_113),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_126),
.C(n_127),
.Y(n_113)
);

XNOR2x2_ASAP7_75t_SL g193 ( 
.A(n_114),
.B(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_116),
.Y(n_119)
);

AOI22x1_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_119),
.B1(n_145),
.B2(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_145),
.C(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_126),
.B(n_127),
.Y(n_194)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_141),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_130),
.B(n_142),
.C(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_140),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_135),
.C(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_139),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

XOR2x1_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_145),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_150),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_149),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_178),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_171),
.B2(n_172),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_231),
.B(n_556),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_184),
.A2(n_558),
.B(n_559),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_185),
.B(n_188),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.C(n_195),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_193),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_195),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_215),
.C(n_228),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.C(n_213),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_198),
.B(n_334),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_199),
.B(n_300),
.C(n_302),
.Y(n_299)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_203),
.B(n_213),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_204),
.B(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_228),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_224),
.C(n_227),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.C(n_221),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_221),
.Y(n_242)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2x1_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_242),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_280),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_277),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_SL g558 ( 
.A(n_234),
.B(n_277),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.C(n_239),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g385 ( 
.A(n_235),
.B(n_237),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_239),
.B(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_258),
.C(n_274),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_240),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.C(n_255),
.Y(n_240)
);

XNOR2x2_ASAP7_75t_SL g343 ( 
.A(n_241),
.B(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_243),
.B(n_255),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.C(n_252),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_244),
.A2(n_252),
.B1(n_253),
.B2(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_244),
.Y(n_382)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_247),
.B(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_251),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_252),
.B(n_436),
.C(n_438),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_252),
.A2(n_253),
.B1(n_436),
.B2(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_258),
.B(n_275),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_268),
.C(n_271),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_259),
.B(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_264),
.Y(n_288)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_267),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_268),
.A2(n_271),
.B1(n_272),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx8_ASAP7_75t_L g515 ( 
.A(n_270),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_271),
.A2(n_272),
.B1(n_417),
.B2(n_418),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_272),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

AO21x2_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_389),
.B(n_553),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_383),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_337),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_283),
.B(n_337),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_330),
.Y(n_283)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_284),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_303),
.C(n_325),
.Y(n_284)
);

INVxp33_ASAP7_75t_SL g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.C(n_299),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_287),
.B(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_289),
.A2(n_290),
.B1(n_299),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx12f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_299),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_350),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_302),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_304),
.A2(n_326),
.B1(n_327),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_315),
.C(n_320),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_305),
.B(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_309),
.C(n_311),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_306),
.A2(n_311),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_306),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_306),
.B(n_456),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_308),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_309),
.B(n_401),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_311),
.Y(n_403)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_313),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_315),
.A2(n_316),
.B1(n_320),
.B2(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_320),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_333),
.B1(n_335),
.B2(n_336),
.Y(n_330)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_333),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_333),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_335),
.B(n_387),
.C(n_388),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_343),
.C(n_345),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_339),
.A2(n_340),
.B1(n_343),
.B2(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_343),
.Y(n_394)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_346),
.B(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_376),
.C(n_380),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_398),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_352),
.C(n_360),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2x1_ASAP7_75t_SL g443 ( 
.A(n_349),
.B(n_444),
.Y(n_443)
);

XNOR2x1_ASAP7_75t_L g444 ( 
.A(n_352),
.B(n_360),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_357),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_353),
.B(n_357),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_367),
.C(n_371),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_361),
.A2(n_367),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_361),
.Y(n_432)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_367),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_367),
.A2(n_433),
.B1(n_501),
.B2(n_502),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_367),
.B(n_501),
.C(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XOR2x1_ASAP7_75t_SL g430 ( 
.A(n_371),
.B(n_431),
.Y(n_430)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_380),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_383),
.A2(n_554),
.B(n_555),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_384),
.B(n_386),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_447),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_395),
.C(n_424),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_392),
.B(n_396),
.Y(n_449)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_399),
.C(n_420),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_421),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_404),
.C(n_412),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_404),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_402),
.B(n_457),
.C(n_461),
.Y(n_480)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx6_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_427),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_416),
.C(n_417),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g541 ( 
.A(n_413),
.B(n_542),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

XNOR2x1_ASAP7_75t_SL g487 ( 
.A(n_414),
.B(n_415),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_414),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_414),
.A2(n_505),
.B1(n_506),
.B2(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NOR2x1_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_445),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_445),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.C(n_443),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_426),
.B(n_551),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_429),
.B(n_443),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_434),
.C(n_441),
.Y(n_429)
);

XOR2x1_ASAP7_75t_L g536 ( 
.A(n_430),
.B(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_435),
.B(n_442),
.Y(n_537)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_436),
.Y(n_483)
);

XOR2x2_ASAP7_75t_L g481 ( 
.A(n_438),
.B(n_482),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.C(n_450),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_451),
.A2(n_548),
.B(n_552),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_533),
.B(n_547),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_495),
.B(n_532),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_478),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_454),
.B(n_478),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_463),
.C(n_472),
.Y(n_454)
);

XOR2x1_ASAP7_75t_SL g526 ( 
.A(n_455),
.B(n_527),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_461),
.Y(n_456)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_463),
.A2(n_464),
.B1(n_472),
.B2(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_471),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_471),
.Y(n_499)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_472),
.Y(n_528)
);

AO22x1_ASAP7_75t_SL g472 ( 
.A1(n_473),
.A2(n_475),
.B1(n_476),
.B2(n_477),
.Y(n_472)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_473),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_475),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_475),
.B(n_476),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_477),
.B(n_519),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_484),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_480),
.B(n_481),
.C(n_546),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_484),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

MAJx2_ASAP7_75t_L g544 ( 
.A(n_485),
.B(n_487),
.C(n_488),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

AOI21x1_ASAP7_75t_L g495 ( 
.A1(n_496),
.A2(n_525),
.B(n_531),
.Y(n_495)
);

OAI21x1_ASAP7_75t_SL g496 ( 
.A1(n_497),
.A2(n_509),
.B(n_524),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_504),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_498),
.B(n_504),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_499),
.Y(n_530)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_505),
.B(n_506),
.Y(n_504)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_506),
.Y(n_517)
);

INVx6_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_518),
.B(n_523),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_516),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_516),
.Y(n_523)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_526),
.B(n_529),
.Y(n_525)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_526),
.B(n_529),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_534),
.B(n_545),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_545),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_535),
.A2(n_536),
.B1(n_538),
.B2(n_539),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_535),
.B(n_540),
.C(n_544),
.Y(n_549)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_540),
.A2(n_541),
.B1(n_543),
.B2(n_544),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_550),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_549),
.B(n_550),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);


endmodule