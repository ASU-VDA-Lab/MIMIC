module real_aes_12134_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_552;
wire n_590;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1250;
wire n_1095;
wire n_360;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_315;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1014;
wire n_742;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_265;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1162;
wire n_762;
wire n_325;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_974;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_304;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_244;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_338;
wire n_698;
wire n_371;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_340;
wire n_483;
wire n_1280;
wire n_394;
wire n_729;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_0), .A2(n_203), .B1(n_468), .B2(n_470), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_0), .A2(n_203), .B1(n_450), .B2(n_454), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_1), .A2(n_11), .B1(n_435), .B2(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g686 ( .A(n_1), .Y(n_686) );
INVx1_ASAP7_75t_L g434 ( .A(n_2), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_2), .A2(n_126), .B1(n_463), .B2(n_464), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_3), .A2(n_17), .B1(n_352), .B2(n_381), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_3), .A2(n_221), .B1(n_390), .B2(n_392), .Y(n_898) );
INVx1_ASAP7_75t_L g1009 ( .A(n_4), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_5), .A2(n_8), .B1(n_327), .B2(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g491 ( .A(n_5), .Y(n_491) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_6), .Y(n_248) );
INVx1_ASAP7_75t_L g307 ( .A(n_6), .Y(n_307) );
INVx1_ASAP7_75t_L g644 ( .A(n_7), .Y(n_644) );
INVx1_ASAP7_75t_L g493 ( .A(n_8), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_9), .A2(n_38), .B1(n_838), .B2(n_840), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_9), .A2(n_38), .B1(n_577), .B2(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g754 ( .A(n_10), .Y(n_754) );
INVx1_ASAP7_75t_L g683 ( .A(n_11), .Y(n_683) );
INVx1_ASAP7_75t_L g809 ( .A(n_12), .Y(n_809) );
INVxp33_ASAP7_75t_SL g952 ( .A(n_13), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_13), .A2(n_227), .B1(n_586), .B2(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g1121 ( .A(n_14), .Y(n_1121) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_15), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_16), .Y(n_425) );
INVx1_ASAP7_75t_L g884 ( .A(n_17), .Y(n_884) );
INVx1_ASAP7_75t_L g432 ( .A(n_18), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_18), .A2(n_231), .B1(n_459), .B2(n_460), .Y(n_458) );
AO221x2_ASAP7_75t_L g1030 ( .A1(n_19), .A2(n_54), .B1(n_1007), .B2(n_1029), .C(n_1031), .Y(n_1030) );
XNOR2xp5_ASAP7_75t_L g852 ( .A(n_20), .B(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g1048 ( .A(n_20), .Y(n_1048) );
INVxp33_ASAP7_75t_L g566 ( .A(n_21), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_21), .A2(n_198), .B1(n_611), .B2(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g313 ( .A(n_22), .Y(n_313) );
INVx1_ASAP7_75t_L g1032 ( .A(n_23), .Y(n_1032) );
INVxp33_ASAP7_75t_SL g764 ( .A(n_24), .Y(n_764) );
AOI22xp5_ASAP7_75t_SL g795 ( .A1(n_24), .A2(n_63), .B1(n_796), .B2(n_798), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_25), .A2(n_200), .B1(n_444), .B2(n_914), .Y(n_913) );
INVxp67_ASAP7_75t_SL g942 ( .A(n_25), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_26), .A2(n_177), .B1(n_528), .B2(n_924), .Y(n_923) );
OAI211xp5_ASAP7_75t_SL g927 ( .A1(n_26), .A2(n_399), .B(n_928), .C(n_931), .Y(n_927) );
BUFx2_ASAP7_75t_L g269 ( .A(n_27), .Y(n_269) );
BUFx2_ASAP7_75t_L g335 ( .A(n_27), .Y(n_335) );
INVx1_ASAP7_75t_L g608 ( .A(n_27), .Y(n_608) );
AO22x1_ASAP7_75t_L g746 ( .A1(n_28), .A2(n_747), .B1(n_748), .B2(n_800), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_28), .Y(n_747) );
INVx1_ASAP7_75t_L g1225 ( .A(n_29), .Y(n_1225) );
AOI22xp33_ASAP7_75t_SL g1239 ( .A1(n_29), .A2(n_191), .B1(n_463), .B2(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1119 ( .A(n_30), .Y(n_1119) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_31), .A2(n_100), .B1(n_531), .B2(n_532), .Y(n_530) );
INVxp67_ASAP7_75t_L g544 ( .A(n_31), .Y(n_544) );
INVx1_ASAP7_75t_L g957 ( .A(n_32), .Y(n_957) );
AOI22xp33_ASAP7_75t_SL g971 ( .A1(n_32), .A2(n_70), .B1(n_592), .B2(n_972), .Y(n_971) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_33), .A2(n_190), .B1(n_592), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_33), .A2(n_190), .B1(n_435), .B2(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g812 ( .A(n_34), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_34), .A2(n_90), .B1(n_464), .B2(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g1004 ( .A(n_35), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_35), .B(n_1014), .Y(n_1017) );
AOI22xp33_ASAP7_75t_SL g773 ( .A1(n_36), .A2(n_159), .B1(n_603), .B2(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_36), .A2(n_159), .B1(n_791), .B2(n_794), .Y(n_790) );
INVx1_ASAP7_75t_L g814 ( .A(n_37), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_37), .A2(n_136), .B1(n_541), .B2(n_710), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_39), .A2(n_166), .B1(n_464), .B2(n_524), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_39), .A2(n_166), .B1(n_470), .B2(n_527), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_40), .A2(n_49), .B1(n_459), .B2(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_40), .A2(n_49), .B1(n_474), .B2(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g896 ( .A(n_41), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_42), .A2(n_139), .B1(n_966), .B2(n_967), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_42), .A2(n_139), .B1(n_734), .B2(n_977), .Y(n_976) );
INVxp67_ASAP7_75t_L g712 ( .A(n_43), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_43), .A2(n_111), .B1(n_740), .B2(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g575 ( .A(n_44), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_44), .A2(n_127), .B1(n_592), .B2(n_603), .Y(n_602) );
CKINVDCx16_ASAP7_75t_R g1045 ( .A(n_45), .Y(n_1045) );
INVx1_ASAP7_75t_L g1115 ( .A(n_46), .Y(n_1115) );
OAI211xp5_ASAP7_75t_L g641 ( .A1(n_47), .A2(n_341), .B(n_374), .C(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_SL g659 ( .A1(n_47), .A2(n_189), .B1(n_593), .B2(n_651), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_48), .A2(n_223), .B1(n_330), .B2(n_345), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_48), .A2(n_168), .B1(n_390), .B2(n_392), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_50), .A2(n_129), .B1(n_464), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_50), .A2(n_129), .B1(n_528), .B2(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g959 ( .A(n_51), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_51), .A2(n_208), .B1(n_488), .B2(n_541), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_52), .A2(n_167), .B1(n_599), .B2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_52), .A2(n_167), .B1(n_665), .B2(n_667), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g1218 ( .A(n_53), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_55), .A2(n_205), .B1(n_527), .B2(n_528), .Y(n_526) );
INVxp33_ASAP7_75t_L g546 ( .A(n_55), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_56), .A2(n_194), .B1(n_450), .B2(n_464), .Y(n_915) );
INVx1_ASAP7_75t_L g938 ( .A(n_56), .Y(n_938) );
AOI22xp33_ASAP7_75t_SL g964 ( .A1(n_57), .A2(n_120), .B1(n_592), .B2(n_782), .Y(n_964) );
AOI22xp33_ASAP7_75t_SL g978 ( .A1(n_57), .A2(n_120), .B1(n_435), .B2(n_673), .Y(n_978) );
INVx1_ASAP7_75t_L g767 ( .A(n_58), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_58), .A2(n_130), .B1(n_509), .B2(n_791), .Y(n_799) );
INVx1_ASAP7_75t_L g297 ( .A(n_59), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_59), .A2(n_168), .B1(n_348), .B2(n_352), .Y(n_347) );
INVx1_ASAP7_75t_L g699 ( .A(n_60), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_60), .A2(n_76), .B1(n_651), .B2(n_720), .Y(n_727) );
INVx1_ASAP7_75t_L g1057 ( .A(n_61), .Y(n_1057) );
CKINVDCx16_ASAP7_75t_R g1062 ( .A(n_62), .Y(n_1062) );
INVxp33_ASAP7_75t_SL g765 ( .A(n_63), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_64), .A2(n_222), .B1(n_468), .B2(n_470), .Y(n_477) );
INVx1_ASAP7_75t_L g484 ( .A(n_64), .Y(n_484) );
INVx1_ASAP7_75t_L g895 ( .A(n_65), .Y(n_895) );
INVx1_ASAP7_75t_L g696 ( .A(n_66), .Y(n_696) );
INVx1_ASAP7_75t_L g865 ( .A(n_67), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_68), .A2(n_209), .B1(n_586), .B2(n_589), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_68), .A2(n_209), .B1(n_614), .B2(n_616), .Y(n_613) );
INVxp67_ASAP7_75t_SL g822 ( .A(n_69), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_69), .A2(n_135), .B1(n_740), .B2(n_796), .Y(n_848) );
INVxp33_ASAP7_75t_SL g950 ( .A(n_70), .Y(n_950) );
INVx1_ASAP7_75t_L g1015 ( .A(n_71), .Y(n_1015) );
AOI22xp33_ASAP7_75t_SL g1235 ( .A1(n_72), .A2(n_229), .B1(n_444), .B2(n_448), .Y(n_1235) );
AOI22xp33_ASAP7_75t_SL g1243 ( .A1(n_72), .A2(n_229), .B1(n_327), .B2(n_919), .Y(n_1243) );
INVx1_ASAP7_75t_L g563 ( .A(n_73), .Y(n_563) );
INVx1_ASAP7_75t_L g291 ( .A(n_74), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_74), .A2(n_155), .B1(n_379), .B2(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g870 ( .A(n_75), .Y(n_870) );
OAI211xp5_ASAP7_75t_SL g899 ( .A1(n_75), .A2(n_397), .B(n_399), .C(n_900), .Y(n_899) );
INVxp33_ASAP7_75t_SL g693 ( .A(n_76), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_77), .A2(n_196), .B1(n_586), .B2(n_777), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_77), .A2(n_196), .B1(n_787), .B2(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g761 ( .A(n_78), .Y(n_761) );
INVxp33_ASAP7_75t_SL g807 ( .A(n_79), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_79), .A2(n_153), .B1(n_459), .B2(n_828), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g1022 ( .A1(n_80), .A2(n_124), .B1(n_1023), .B2(n_1026), .Y(n_1022) );
AOI222xp33_ASAP7_75t_L g1208 ( .A1(n_80), .A2(n_1209), .B1(n_1268), .B2(n_1272), .C1(n_1276), .C2(n_1280), .Y(n_1208) );
AO22x2_ASAP7_75t_L g1210 ( .A1(n_80), .A2(n_1211), .B1(n_1250), .B2(n_1251), .Y(n_1210) );
INVxp67_ASAP7_75t_L g1250 ( .A(n_80), .Y(n_1250) );
CKINVDCx16_ASAP7_75t_R g1064 ( .A(n_81), .Y(n_1064) );
INVx1_ASAP7_75t_L g511 ( .A(n_82), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_82), .A2(n_86), .B1(n_488), .B2(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g945 ( .A(n_83), .Y(n_945) );
INVx1_ASAP7_75t_L g312 ( .A(n_84), .Y(n_312) );
INVx1_ASAP7_75t_L g933 ( .A(n_85), .Y(n_933) );
INVx1_ASAP7_75t_L g512 ( .A(n_86), .Y(n_512) );
INVx1_ASAP7_75t_L g343 ( .A(n_87), .Y(n_343) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_87), .A2(n_397), .B(n_399), .C(n_405), .Y(n_396) );
INVx1_ASAP7_75t_L g859 ( .A(n_88), .Y(n_859) );
INVxp67_ASAP7_75t_SL g706 ( .A(n_89), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_89), .A2(n_119), .B1(n_730), .B2(n_738), .Y(n_737) );
INVxp33_ASAP7_75t_SL g806 ( .A(n_90), .Y(n_806) );
INVx1_ASAP7_75t_L g888 ( .A(n_91), .Y(n_888) );
INVx1_ASAP7_75t_L g439 ( .A(n_92), .Y(n_439) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_92), .A2(n_174), .B1(n_487), .B2(n_488), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_93), .A2(n_133), .B1(n_327), .B2(n_474), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_93), .A2(n_133), .B1(n_392), .B2(n_413), .Y(n_926) );
INVx1_ASAP7_75t_L g1214 ( .A(n_94), .Y(n_1214) );
AOI22xp33_ASAP7_75t_SL g1249 ( .A1(n_94), .A2(n_148), .B1(n_520), .B2(n_531), .Y(n_1249) );
AOI22xp5_ASAP7_75t_L g1273 ( .A1(n_95), .A2(n_1251), .B1(n_1274), .B2(n_1275), .Y(n_1273) );
CKINVDCx5p33_ASAP7_75t_R g1274 ( .A(n_95), .Y(n_1274) );
INVxp67_ASAP7_75t_SL g284 ( .A(n_96), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_96), .A2(n_178), .B1(n_327), .B2(n_330), .Y(n_326) );
INVx1_ASAP7_75t_L g1047 ( .A(n_97), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_98), .A2(n_185), .B1(n_450), .B2(n_707), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1242 ( .A1(n_98), .A2(n_185), .B1(n_629), .B2(n_738), .Y(n_1242) );
INVxp33_ASAP7_75t_SL g751 ( .A(n_99), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g781 ( .A1(n_99), .A2(n_232), .B1(n_774), .B2(n_782), .Y(n_781) );
INVxp33_ASAP7_75t_L g543 ( .A(n_100), .Y(n_543) );
AO221x2_ASAP7_75t_L g1000 ( .A1(n_101), .A2(n_165), .B1(n_1001), .B2(n_1007), .C(n_1008), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_102), .A2(n_211), .B1(n_667), .B2(n_676), .Y(n_980) );
INVxp67_ASAP7_75t_SL g987 ( .A(n_102), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_103), .A2(n_202), .B1(n_444), .B2(n_448), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_103), .A2(n_202), .B1(n_472), .B2(n_474), .Y(n_471) );
INVx1_ASAP7_75t_L g869 ( .A(n_104), .Y(n_869) );
OAI22xp33_ASAP7_75t_SL g901 ( .A1(n_104), .A2(n_137), .B1(n_249), .B2(n_413), .Y(n_901) );
AO22x2_ASAP7_75t_L g501 ( .A1(n_105), .A2(n_502), .B1(n_549), .B2(n_550), .Y(n_501) );
INVx1_ASAP7_75t_L g549 ( .A(n_105), .Y(n_549) );
INVx1_ASAP7_75t_L g240 ( .A(n_106), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_107), .A2(n_158), .B1(n_676), .B2(n_678), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_107), .A2(n_158), .B1(n_392), .B2(n_413), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_108), .A2(n_177), .B1(n_249), .B2(n_390), .Y(n_934) );
OAI22xp33_ASAP7_75t_L g944 ( .A1(n_108), .A2(n_194), .B1(n_348), .B2(n_352), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g1028 ( .A1(n_109), .A2(n_157), .B1(n_1007), .B2(n_1029), .Y(n_1028) );
XNOR2xp5_ASAP7_75t_L g636 ( .A(n_110), .B(n_637), .Y(n_636) );
INVxp67_ASAP7_75t_L g713 ( .A(n_111), .Y(n_713) );
INVx1_ASAP7_75t_L g514 ( .A(n_112), .Y(n_514) );
INVx1_ASAP7_75t_L g758 ( .A(n_113), .Y(n_758) );
AOI22xp33_ASAP7_75t_SL g979 ( .A1(n_114), .A2(n_224), .B1(n_577), .B2(n_611), .Y(n_979) );
INVxp67_ASAP7_75t_SL g983 ( .A(n_114), .Y(n_983) );
CKINVDCx5p33_ASAP7_75t_R g1222 ( .A(n_115), .Y(n_1222) );
INVxp67_ASAP7_75t_SL g701 ( .A(n_116), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_116), .A2(n_233), .B1(n_541), .B2(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_117), .A2(n_122), .B1(n_519), .B2(n_520), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_117), .A2(n_122), .B1(n_444), .B2(n_448), .Y(n_535) );
INVx1_ASAP7_75t_L g554 ( .A(n_118), .Y(n_554) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_119), .Y(n_704) );
XOR2xp5_ASAP7_75t_L g261 ( .A(n_121), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g954 ( .A(n_123), .Y(n_954) );
INVxp33_ASAP7_75t_SL g505 ( .A(n_125), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_125), .A2(n_142), .B1(n_454), .B2(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g431 ( .A(n_126), .Y(n_431) );
INVxp33_ASAP7_75t_L g570 ( .A(n_127), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_128), .A2(n_215), .B1(n_352), .B2(n_381), .Y(n_640) );
INVxp33_ASAP7_75t_SL g687 ( .A(n_128), .Y(n_687) );
INVxp33_ASAP7_75t_SL g769 ( .A(n_130), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_131), .A2(n_189), .B1(n_348), .B2(n_379), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_131), .A2(n_215), .B1(n_599), .B2(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_132), .A2(n_138), .B1(n_444), .B2(n_910), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_132), .A2(n_138), .B1(n_345), .B2(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g862 ( .A(n_134), .Y(n_862) );
INVxp33_ASAP7_75t_L g821 ( .A(n_135), .Y(n_821) );
INVx1_ASAP7_75t_L g813 ( .A(n_136), .Y(n_813) );
INVx1_ASAP7_75t_L g872 ( .A(n_137), .Y(n_872) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_140), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_140), .A2(n_182), .B1(n_599), .B2(n_600), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g1035 ( .A1(n_141), .A2(n_149), .B1(n_1023), .B2(n_1026), .Y(n_1035) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_142), .Y(n_508) );
INVxp33_ASAP7_75t_SL g515 ( .A(n_143), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_143), .A2(n_162), .B1(n_444), .B2(n_448), .Y(n_522) );
INVxp33_ASAP7_75t_SL g694 ( .A(n_144), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_144), .A2(n_219), .B1(n_717), .B2(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g883 ( .A(n_145), .Y(n_883) );
OAI22xp33_ASAP7_75t_L g890 ( .A1(n_145), .A2(n_161), .B1(n_348), .B2(n_379), .Y(n_890) );
INVx1_ASAP7_75t_L g277 ( .A(n_146), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_147), .A2(n_216), .B1(n_450), .B2(n_454), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_147), .A2(n_216), .B1(n_468), .B2(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g1215 ( .A(n_148), .Y(n_1215) );
XNOR2xp5_ASAP7_75t_L g689 ( .A(n_149), .B(n_690), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_150), .A2(n_186), .B1(n_1001), .B2(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g558 ( .A(n_151), .Y(n_558) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_152), .Y(n_242) );
AND3x2_ASAP7_75t_L g1005 ( .A(n_152), .B(n_240), .C(n_1006), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_152), .B(n_240), .Y(n_1012) );
INVxp33_ASAP7_75t_SL g810 ( .A(n_153), .Y(n_810) );
INVxp33_ASAP7_75t_SL g824 ( .A(n_154), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_154), .A2(n_199), .B1(n_577), .B2(n_843), .Y(n_847) );
INVx1_ASAP7_75t_L g294 ( .A(n_155), .Y(n_294) );
INVx2_ASAP7_75t_L g253 ( .A(n_156), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_160), .A2(n_204), .B1(n_658), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_160), .A2(n_204), .B1(n_733), .B2(n_734), .Y(n_732) );
INVx1_ASAP7_75t_L g886 ( .A(n_161), .Y(n_886) );
INVxp33_ASAP7_75t_SL g506 ( .A(n_162), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_163), .A2(n_170), .B1(n_1007), .B2(n_1029), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_164), .A2(n_175), .B1(n_720), .B2(n_722), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_164), .A2(n_175), .B1(n_662), .B2(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g1006 ( .A(n_169), .Y(n_1006) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_171), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_171), .A2(n_193), .B1(n_520), .B2(n_624), .Y(n_623) );
CKINVDCx16_ASAP7_75t_R g1043 ( .A(n_172), .Y(n_1043) );
INVx1_ASAP7_75t_L g1117 ( .A(n_173), .Y(n_1117) );
INVx1_ASAP7_75t_L g436 ( .A(n_174), .Y(n_436) );
INVx1_ASAP7_75t_L g1231 ( .A(n_176), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_176), .A2(n_214), .B1(n_459), .B2(n_777), .Y(n_1238) );
INVxp67_ASAP7_75t_SL g279 ( .A(n_178), .Y(n_279) );
INVx1_ASAP7_75t_L g272 ( .A(n_179), .Y(n_272) );
INVx1_ASAP7_75t_L g255 ( .A(n_180), .Y(n_255) );
INVx2_ASAP7_75t_L g268 ( .A(n_180), .Y(n_268) );
XOR2x2_ASAP7_75t_L g946 ( .A(n_181), .B(n_947), .Y(n_946) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_182), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g1073 ( .A1(n_183), .A2(n_212), .B1(n_1023), .B2(n_1026), .Y(n_1073) );
INVx1_ASAP7_75t_L g1217 ( .A(n_184), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_184), .A2(n_228), .B1(n_1246), .B2(n_1247), .Y(n_1245) );
OAI211xp5_ASAP7_75t_L g1254 ( .A1(n_184), .A2(n_399), .B(n_1255), .C(n_1257), .Y(n_1254) );
XNOR2xp5_ASAP7_75t_L g421 ( .A(n_187), .B(n_422), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_188), .Y(n_561) );
INVx1_ASAP7_75t_L g1229 ( .A(n_191), .Y(n_1229) );
OAI211xp5_ASAP7_75t_L g1263 ( .A1(n_191), .A2(n_374), .B(n_1264), .C(n_1266), .Y(n_1263) );
INVx1_ASAP7_75t_L g340 ( .A(n_192), .Y(n_340) );
OAI22xp33_ASAP7_75t_SL g412 ( .A1(n_192), .A2(n_223), .B1(n_249), .B2(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_193), .Y(n_567) );
INVxp33_ASAP7_75t_SL g755 ( .A(n_195), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_195), .A2(n_218), .B1(n_586), .B2(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g1058 ( .A(n_197), .Y(n_1058) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_198), .Y(n_562) );
INVxp67_ASAP7_75t_SL g818 ( .A(n_199), .Y(n_818) );
INVx1_ASAP7_75t_L g943 ( .A(n_200), .Y(n_943) );
INVx1_ASAP7_75t_L g643 ( .A(n_201), .Y(n_643) );
INVxp67_ASAP7_75t_SL g539 ( .A(n_205), .Y(n_539) );
XOR2x2_ASAP7_75t_L g802 ( .A(n_206), .B(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g857 ( .A(n_207), .Y(n_857) );
INVx1_ASAP7_75t_L g960 ( .A(n_208), .Y(n_960) );
INVx1_ASAP7_75t_L g932 ( .A(n_210), .Y(n_932) );
INVxp33_ASAP7_75t_SL g986 ( .A(n_211), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g1219 ( .A(n_213), .Y(n_1219) );
INVx1_ASAP7_75t_L g1226 ( .A(n_214), .Y(n_1226) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_217), .Y(n_370) );
INVxp33_ASAP7_75t_SL g752 ( .A(n_218), .Y(n_752) );
INVxp67_ASAP7_75t_SL g697 ( .A(n_219), .Y(n_697) );
INVx2_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
INVx1_ASAP7_75t_L g874 ( .A(n_221), .Y(n_874) );
INVx1_ASAP7_75t_L g496 ( .A(n_222), .Y(n_496) );
INVxp33_ASAP7_75t_SL g989 ( .A(n_224), .Y(n_989) );
INVx1_ASAP7_75t_L g319 ( .A(n_225), .Y(n_319) );
BUFx3_ASAP7_75t_L g329 ( .A(n_225), .Y(n_329) );
INVx1_ASAP7_75t_L g321 ( .A(n_226), .Y(n_321) );
BUFx3_ASAP7_75t_L g332 ( .A(n_226), .Y(n_332) );
INVxp67_ASAP7_75t_SL g955 ( .A(n_227), .Y(n_955) );
INVx1_ASAP7_75t_L g1221 ( .A(n_228), .Y(n_1221) );
INVx1_ASAP7_75t_L g300 ( .A(n_230), .Y(n_300) );
INVx1_ASAP7_75t_L g426 ( .A(n_231), .Y(n_426) );
INVx1_ASAP7_75t_L g757 ( .A(n_232), .Y(n_757) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_233), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_256), .B(n_992), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_243), .Y(n_237) );
AND2x4_ASAP7_75t_L g1271 ( .A(n_238), .B(n_244), .Y(n_1271) );
NOR2xp33_ASAP7_75t_SL g238 ( .A(n_239), .B(n_241), .Y(n_238) );
INVx1_ASAP7_75t_SL g1279 ( .A(n_239), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_239), .B(n_241), .Y(n_1282) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_241), .B(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_249), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x6_ASAP7_75t_L g417 ( .A(n_246), .B(n_335), .Y(n_417) );
OR2x2_ASAP7_75t_L g548 ( .A(n_246), .B(n_335), .Y(n_548) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g456 ( .A(n_247), .B(n_255), .Y(n_456) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g266 ( .A(n_248), .B(n_267), .Y(n_266) );
INVx8_ASAP7_75t_L g495 ( .A(n_249), .Y(n_495) );
OR2x6_ASAP7_75t_L g249 ( .A(n_250), .B(n_254), .Y(n_249) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_250), .Y(n_271) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_250), .Y(n_296) );
OR2x6_ASAP7_75t_L g390 ( .A(n_250), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_SL g879 ( .A(n_250), .Y(n_879) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g276 ( .A(n_252), .Y(n_276) );
INVx2_ASAP7_75t_L g283 ( .A(n_252), .Y(n_283) );
AND2x4_ASAP7_75t_L g288 ( .A(n_252), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g404 ( .A(n_252), .Y(n_404) );
AND2x2_ASAP7_75t_L g453 ( .A(n_252), .B(n_253), .Y(n_453) );
INVx1_ASAP7_75t_L g275 ( .A(n_253), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_253), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g289 ( .A(n_253), .Y(n_289) );
INVx1_ASAP7_75t_L g407 ( .A(n_253), .Y(n_407) );
INVx1_ASAP7_75t_L g447 ( .A(n_253), .Y(n_447) );
AND2x4_ASAP7_75t_L g406 ( .A(n_254), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g488 ( .A(n_255), .B(n_410), .Y(n_488) );
OR2x2_ASAP7_75t_L g710 ( .A(n_255), .B(n_410), .Y(n_710) );
XNOR2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_632), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_499), .B1(n_630), .B2(n_631), .Y(n_257) );
INVx1_ASAP7_75t_L g630 ( .A(n_258), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_418), .B1(n_419), .B2(n_498), .Y(n_258) );
INVx2_ASAP7_75t_SL g498 ( .A(n_259), .Y(n_498) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND3xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_346), .C(n_388), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_308), .Y(n_263) );
OAI33xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_270), .A3(n_278), .B1(n_290), .B2(n_295), .B3(n_301), .Y(n_264) );
OAI33xp33_ASAP7_75t_L g876 ( .A1(n_265), .A2(n_301), .A3(n_877), .B1(n_880), .B2(n_881), .B3(n_885), .Y(n_876) );
OR2x6_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
INVx1_ASAP7_75t_L g391 ( .A(n_267), .Y(n_391) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g306 ( .A(n_268), .Y(n_306) );
INVx2_ASAP7_75t_L g303 ( .A(n_269), .Y(n_303) );
BUFx2_ASAP7_75t_L g387 ( .A(n_269), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B1(n_273), .B2(n_277), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g314 ( .A1(n_272), .A2(n_277), .B1(n_315), .B2(n_322), .C(n_326), .Y(n_314) );
OAI22xp33_ASAP7_75t_L g877 ( .A1(n_273), .A2(n_862), .B1(n_865), .B2(n_878), .Y(n_877) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g299 ( .A(n_275), .B(n_276), .Y(n_299) );
INVx1_ASAP7_75t_L g410 ( .A(n_276), .Y(n_410) );
OAI22xp33_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_280), .B1(n_284), .B2(n_285), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_280), .A2(n_291), .B1(n_292), .B2(n_294), .Y(n_290) );
OAI22xp33_ASAP7_75t_L g880 ( .A1(n_280), .A2(n_292), .B1(n_857), .B2(n_859), .Y(n_880) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g882 ( .A(n_281), .Y(n_882) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx2_ASAP7_75t_L g415 ( .A(n_282), .Y(n_415) );
AND2x4_ASAP7_75t_L g445 ( .A(n_283), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g726 ( .A(n_286), .Y(n_726) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx3_ASAP7_75t_L g293 ( .A(n_287), .Y(n_293) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_287), .Y(n_461) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g395 ( .A(n_288), .Y(n_395) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_288), .Y(n_448) );
INVx1_ASAP7_75t_L g836 ( .A(n_288), .Y(n_836) );
AND2x4_ASAP7_75t_L g403 ( .A(n_289), .B(n_404), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g881 ( .A1(n_292), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_881) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g590 ( .A(n_293), .Y(n_590) );
BUFx3_ASAP7_75t_L g658 ( .A(n_293), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B1(n_298), .B2(n_300), .Y(n_295) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx2_ASAP7_75t_L g398 ( .A(n_299), .Y(n_398) );
INVx3_ASAP7_75t_L g887 ( .A(n_299), .Y(n_887) );
INVx2_ASAP7_75t_L g930 ( .A(n_299), .Y(n_930) );
AOI222xp33_ASAP7_75t_L g360 ( .A1(n_300), .A2(n_361), .B1(n_365), .B2(n_370), .C1(n_371), .C2(n_373), .Y(n_360) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_302), .B(n_458), .C(n_462), .Y(n_457) );
AOI33xp33_ASAP7_75t_L g517 ( .A1(n_302), .A2(n_475), .A3(n_518), .B1(n_521), .B2(n_522), .B3(n_523), .Y(n_517) );
NAND3xp33_ASAP7_75t_L g1237 ( .A(n_302), .B(n_1238), .C(n_1239), .Y(n_1237) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
OR2x2_ASAP7_75t_L g309 ( .A(n_303), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g455 ( .A(n_303), .B(n_456), .Y(n_455) );
OR2x6_ASAP7_75t_L g619 ( .A(n_303), .B(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g655 ( .A(n_303), .B(n_456), .Y(n_655) );
OR2x2_ASAP7_75t_L g670 ( .A(n_303), .B(n_620), .Y(n_670) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x6_ASAP7_75t_L g606 ( .A(n_305), .B(n_607), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g402 ( .A(n_306), .Y(n_402) );
OAI22xp5_ASAP7_75t_SL g308 ( .A1(n_309), .A2(n_314), .B1(n_333), .B2(n_338), .Y(n_308) );
INVx3_ASAP7_75t_L g475 ( .A(n_309), .Y(n_475) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g620 ( .A(n_311), .Y(n_620) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x4_ASAP7_75t_L g336 ( .A(n_312), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g386 ( .A(n_312), .Y(n_386) );
INVx2_ASAP7_75t_L g337 ( .A(n_313), .Y(n_337) );
INVx1_ASAP7_75t_L g351 ( .A(n_313), .Y(n_351) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_313), .Y(n_355) );
INVx1_ASAP7_75t_L g366 ( .A(n_313), .Y(n_366) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g339 ( .A(n_316), .Y(n_339) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g348 ( .A(n_317), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g864 ( .A(n_317), .Y(n_864) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
AND2x2_ASAP7_75t_L g325 ( .A(n_318), .B(n_320), .Y(n_325) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g331 ( .A(n_319), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g328 ( .A(n_321), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g342 ( .A(n_325), .Y(n_342) );
BUFx4f_ASAP7_75t_L g867 ( .A(n_325), .Y(n_867) );
INVx1_ASAP7_75t_L g1265 ( .A(n_325), .Y(n_1265) );
INVx2_ASAP7_75t_L g666 ( .A(n_327), .Y(n_666) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_328), .Y(n_345) );
AND2x6_ASAP7_75t_L g380 ( .A(n_328), .B(n_350), .Y(n_380) );
INVx2_ASAP7_75t_SL g473 ( .A(n_328), .Y(n_473) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_328), .Y(n_519) );
BUFx3_ASAP7_75t_L g531 ( .A(n_328), .Y(n_531) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_328), .Y(n_733) );
BUFx2_ASAP7_75t_L g845 ( .A(n_328), .Y(n_845) );
INVx2_ASAP7_75t_L g357 ( .A(n_329), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_329), .B(n_332), .Y(n_364) );
INVx1_ASAP7_75t_L g668 ( .A(n_330), .Y(n_668) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_330), .Y(n_734) );
INVx1_ASAP7_75t_L g860 ( .A(n_330), .Y(n_860) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_331), .Y(n_384) );
INVx2_ASAP7_75t_L g534 ( .A(n_331), .Y(n_534) );
INVx1_ASAP7_75t_L g617 ( .A(n_331), .Y(n_617) );
INVx1_ASAP7_75t_L g920 ( .A(n_331), .Y(n_920) );
INVx2_ASAP7_75t_L g358 ( .A(n_332), .Y(n_358) );
INVx1_ASAP7_75t_L g622 ( .A(n_333), .Y(n_622) );
INVx4_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx4f_ASAP7_75t_L g679 ( .A(n_334), .Y(n_679) );
BUFx4f_ASAP7_75t_L g743 ( .A(n_334), .Y(n_743) );
AOI33xp33_ASAP7_75t_L g784 ( .A1(n_334), .A2(n_785), .A3(n_786), .B1(n_790), .B2(n_795), .B3(n_799), .Y(n_784) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
AND2x4_ASAP7_75t_L g481 ( .A(n_335), .B(n_336), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_341), .B2(n_343), .C(n_344), .Y(n_338) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g677 ( .A(n_345), .Y(n_677) );
OAI31xp33_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_359), .A3(n_378), .B(n_385), .Y(n_346) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g376 ( .A(n_350), .Y(n_376) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x6_ASAP7_75t_L g371 ( .A(n_351), .B(n_372), .Y(n_371) );
INVx4_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_353), .A2(n_382), .B1(n_425), .B2(n_426), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_353), .A2(n_382), .B1(n_514), .B2(n_515), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_353), .A2(n_382), .B1(n_558), .B2(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_353), .A2(n_382), .B1(n_696), .B2(n_697), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_353), .A2(n_382), .B1(n_754), .B2(n_755), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_353), .A2(n_382), .B1(n_809), .B2(n_810), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_353), .A2(n_382), .B1(n_954), .B2(n_955), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g1230 ( .A1(n_353), .A2(n_382), .B1(n_1222), .B2(n_1231), .Y(n_1230) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
AND2x2_ASAP7_75t_SL g437 ( .A(n_354), .B(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g579 ( .A(n_354), .B(n_438), .Y(n_579) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx6_ASAP7_75t_L g430 ( .A(n_356), .Y(n_430) );
INVx2_ASAP7_75t_L g469 ( .A(n_356), .Y(n_469) );
BUFx2_ASAP7_75t_L g738 ( .A(n_356), .Y(n_738) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g372 ( .A(n_357), .Y(n_372) );
INVx1_ASAP7_75t_L g369 ( .A(n_358), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_360), .B(n_374), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
BUFx3_ASAP7_75t_L g435 ( .A(n_363), .Y(n_435) );
INVx1_ASAP7_75t_L g510 ( .A(n_363), .Y(n_510) );
BUFx4f_ASAP7_75t_L g577 ( .A(n_363), .Y(n_577) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_363), .Y(n_629) );
INVx1_ASAP7_75t_L g940 ( .A(n_363), .Y(n_940) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_364), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g893 ( .A1(n_365), .A2(n_371), .B1(n_888), .B2(n_894), .C1(n_895), .C2(n_896), .Y(n_893) );
AOI222xp33_ASAP7_75t_L g937 ( .A1(n_365), .A2(n_371), .B1(n_932), .B2(n_933), .C1(n_938), .C2(n_939), .Y(n_937) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_SL g383 ( .A(n_366), .Y(n_383) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g438 ( .A(n_368), .Y(n_438) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_370), .A2(n_373), .B1(n_406), .B2(n_408), .Y(n_405) );
AOI222xp33_ASAP7_75t_L g433 ( .A1(n_371), .A2(n_434), .B1(n_435), .B2(n_436), .C1(n_437), .C2(n_439), .Y(n_433) );
AOI222xp33_ASAP7_75t_L g507 ( .A1(n_371), .A2(n_437), .B1(n_508), .B2(n_509), .C1(n_511), .C2(n_512), .Y(n_507) );
AOI222xp33_ASAP7_75t_L g574 ( .A1(n_371), .A2(n_561), .B1(n_563), .B2(n_575), .C1(n_576), .C2(n_578), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_371), .A2(n_579), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_371), .A2(n_437), .B1(n_627), .B2(n_699), .C1(n_700), .C2(n_701), .Y(n_698) );
AOI222xp33_ASAP7_75t_L g756 ( .A1(n_371), .A2(n_435), .B1(n_757), .B2(n_758), .C1(n_759), .C2(n_761), .Y(n_756) );
AOI222xp33_ASAP7_75t_L g811 ( .A1(n_371), .A2(n_437), .B1(n_730), .B2(n_812), .C1(n_813), .C2(n_814), .Y(n_811) );
AOI222xp33_ASAP7_75t_L g956 ( .A1(n_371), .A2(n_578), .B1(n_957), .B2(n_958), .C1(n_959), .C2(n_960), .Y(n_956) );
AOI222xp33_ASAP7_75t_L g1227 ( .A1(n_371), .A2(n_578), .B1(n_1218), .B2(n_1219), .C1(n_1228), .C2(n_1229), .Y(n_1227) );
AOI22xp33_ASAP7_75t_SL g1266 ( .A1(n_371), .A2(n_579), .B1(n_1218), .B2(n_1219), .Y(n_1266) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_374), .B(n_504), .C(n_507), .D(n_513), .Y(n_503) );
NAND4xp25_ASAP7_75t_SL g691 ( .A(n_374), .B(n_692), .C(n_695), .D(n_698), .Y(n_691) );
NAND4xp25_ASAP7_75t_L g804 ( .A(n_374), .B(n_805), .C(n_808), .D(n_811), .Y(n_804) );
NAND2xp5_ASAP7_75t_SL g892 ( .A(n_374), .B(n_893), .Y(n_892) );
NAND3xp33_ASAP7_75t_SL g936 ( .A(n_374), .B(n_937), .C(n_941), .Y(n_936) );
CKINVDCx8_ASAP7_75t_R g374 ( .A(n_375), .Y(n_374) );
INVx5_ASAP7_75t_L g440 ( .A(n_375), .Y(n_440) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_377), .Y(n_470) );
INVx2_ASAP7_75t_L g529 ( .A(n_377), .Y(n_529) );
BUFx6f_ASAP7_75t_L g731 ( .A(n_377), .Y(n_731) );
INVx1_ASAP7_75t_L g1248 ( .A(n_377), .Y(n_1248) );
CKINVDCx6p67_ASAP7_75t_R g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_380), .A2(n_428), .B1(n_431), .B2(n_432), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_380), .A2(n_428), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_380), .A2(n_428), .B1(n_570), .B2(n_571), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_380), .A2(n_428), .B1(n_693), .B2(n_694), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_380), .A2(n_428), .B1(n_751), .B2(n_752), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_380), .A2(n_428), .B1(n_806), .B2(n_807), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_380), .A2(n_382), .B1(n_942), .B2(n_943), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_380), .A2(n_950), .B1(n_951), .B2(n_952), .Y(n_949) );
AOI22xp5_ASAP7_75t_SL g1224 ( .A1(n_380), .A2(n_951), .B1(n_1225), .B2(n_1226), .Y(n_1224) );
INVx4_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x6_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
AND2x4_ASAP7_75t_L g428 ( .A(n_383), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_L g951 ( .A(n_383), .B(n_429), .Y(n_951) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_384), .Y(n_474) );
INVx1_ASAP7_75t_L g480 ( .A(n_384), .Y(n_480) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_384), .Y(n_520) );
INVx1_ASAP7_75t_L g742 ( .A(n_384), .Y(n_742) );
INVx2_ASAP7_75t_L g873 ( .A(n_384), .Y(n_873) );
AOI211xp5_ASAP7_75t_L g422 ( .A1(n_385), .A2(n_423), .B(n_441), .C(n_482), .Y(n_422) );
AOI211x1_ASAP7_75t_L g502 ( .A1(n_385), .A2(n_503), .B(n_516), .C(n_537), .Y(n_502) );
OAI31xp33_ASAP7_75t_L g638 ( .A1(n_385), .A2(n_639), .A3(n_640), .B(n_641), .Y(n_638) );
OAI31xp33_ASAP7_75t_L g889 ( .A1(n_385), .A2(n_890), .A3(n_891), .B(n_892), .Y(n_889) );
OAI21xp5_ASAP7_75t_SL g935 ( .A1(n_385), .A2(n_936), .B(n_944), .Y(n_935) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AND2x4_ASAP7_75t_L g582 ( .A(n_386), .B(n_387), .Y(n_582) );
OAI31xp33_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_396), .A3(n_412), .B(n_416), .Y(n_388) );
INVx4_ASAP7_75t_L g497 ( .A(n_390), .Y(n_497) );
INVx5_ASAP7_75t_L g547 ( .A(n_390), .Y(n_547) );
AND2x4_ASAP7_75t_L g393 ( .A(n_391), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g414 ( .A(n_391), .Y(n_414) );
AND2x4_ASAP7_75t_L g490 ( .A(n_391), .B(n_445), .Y(n_490) );
AND2x4_ASAP7_75t_L g492 ( .A(n_391), .B(n_394), .Y(n_492) );
INVx5_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
AOI22xp5_ASAP7_75t_SL g711 ( .A1(n_393), .A2(n_490), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_393), .A2(n_490), .B1(n_764), .B2(n_765), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_393), .A2(n_490), .B1(n_986), .B2(n_987), .Y(n_985) );
AOI22xp5_ASAP7_75t_L g1213 ( .A1(n_393), .A2(n_490), .B1(n_1214), .B2(n_1215), .Y(n_1213) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_395), .Y(n_780) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND4xp25_ASAP7_75t_L g556 ( .A(n_399), .B(n_557), .C(n_560), .D(n_565), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_399), .B(n_682), .C(n_685), .Y(n_681) );
NAND4xp25_ASAP7_75t_SL g762 ( .A(n_399), .B(n_763), .C(n_766), .D(n_768), .Y(n_762) );
NAND4xp25_ASAP7_75t_L g1212 ( .A(n_399), .B(n_1213), .C(n_1216), .D(n_1220), .Y(n_1212) );
CKINVDCx11_ASAP7_75t_R g399 ( .A(n_400), .Y(n_399) );
AOI211xp5_ASAP7_75t_L g483 ( .A1(n_400), .A2(n_484), .B(n_485), .C(n_486), .Y(n_483) );
AOI211xp5_ASAP7_75t_L g538 ( .A1(n_400), .A2(n_485), .B(n_539), .C(n_540), .Y(n_538) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_400), .A2(n_706), .B(n_707), .C(n_709), .Y(n_705) );
AOI211xp5_ASAP7_75t_L g816 ( .A1(n_400), .A2(n_817), .B(n_818), .C(n_819), .Y(n_816) );
AOI211xp5_ASAP7_75t_SL g982 ( .A1(n_400), .A2(n_707), .B(n_983), .C(n_984), .Y(n_982) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g411 ( .A(n_402), .Y(n_411) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_403), .Y(n_454) );
BUFx3_ASAP7_75t_L g465 ( .A(n_403), .Y(n_465) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_403), .Y(n_653) );
INVx1_ASAP7_75t_L g708 ( .A(n_403), .Y(n_708) );
BUFx2_ASAP7_75t_L g974 ( .A(n_403), .Y(n_974) );
BUFx3_ASAP7_75t_L g1240 ( .A(n_403), .Y(n_1240) );
INVx2_ASAP7_75t_L g487 ( .A(n_406), .Y(n_487) );
INVx2_ASAP7_75t_L g541 ( .A(n_406), .Y(n_541) );
AOI222xp33_ASAP7_75t_L g682 ( .A1(n_406), .A2(n_643), .B1(n_644), .B2(n_653), .C1(n_683), .C2(n_684), .Y(n_682) );
AOI222xp33_ASAP7_75t_L g766 ( .A1(n_406), .A2(n_408), .B1(n_651), .B2(n_758), .C1(n_761), .C2(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_406), .A2(n_408), .B1(n_895), .B2(n_896), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_406), .A2(n_408), .B1(n_932), .B2(n_933), .Y(n_931) );
INVx2_ASAP7_75t_L g1259 ( .A(n_406), .Y(n_1259) );
AOI222xp33_ASAP7_75t_L g560 ( .A1(n_408), .A2(n_485), .B1(n_561), .B2(n_562), .C1(n_563), .C2(n_564), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_408), .A2(n_1218), .B1(n_1219), .B2(n_1258), .Y(n_1257) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
AND2x4_ASAP7_75t_L g684 ( .A(n_409), .B(n_411), .Y(n_684) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_416), .A2(n_556), .B1(n_568), .B2(n_580), .C(n_583), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_416), .A2(n_681), .B(n_688), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_416), .A2(n_582), .B1(n_749), .B2(n_762), .C(n_770), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_416), .A2(n_582), .B1(n_804), .B2(n_815), .C(n_825), .Y(n_803) );
OAI31xp33_ASAP7_75t_SL g897 ( .A1(n_416), .A2(n_898), .A3(n_899), .B(n_901), .Y(n_897) );
OAI31xp33_ASAP7_75t_SL g925 ( .A1(n_416), .A2(n_926), .A3(n_927), .B(n_934), .Y(n_925) );
AOI221x1_ASAP7_75t_L g1211 ( .A1(n_416), .A2(n_961), .B1(n_1212), .B2(n_1223), .C(n_1232), .Y(n_1211) );
OAI31xp33_ASAP7_75t_L g1252 ( .A1(n_416), .A2(n_1253), .A3(n_1254), .B(n_1260), .Y(n_1252) );
CKINVDCx16_ASAP7_75t_R g416 ( .A(n_417), .Y(n_416) );
AOI31xp33_ASAP7_75t_L g482 ( .A1(n_417), .A2(n_483), .A3(n_489), .B(n_494), .Y(n_482) );
AOI31xp33_ASAP7_75t_L g702 ( .A1(n_417), .A2(n_703), .A3(n_705), .B(n_711), .Y(n_702) );
AOI31xp33_ASAP7_75t_L g981 ( .A1(n_417), .A2(n_982), .A3(n_985), .B(n_988), .Y(n_981) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND4xp25_ASAP7_75t_L g423 ( .A(n_424), .B(n_427), .C(n_433), .D(n_440), .Y(n_423) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_425), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_494) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g612 ( .A(n_430), .Y(n_612) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_430), .Y(n_663) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_430), .Y(n_674) );
INVx2_ASAP7_75t_L g793 ( .A(n_430), .Y(n_793) );
INVx1_ASAP7_75t_L g924 ( .A(n_430), .Y(n_924) );
NAND4xp25_ASAP7_75t_L g568 ( .A(n_440), .B(n_569), .C(n_572), .D(n_574), .Y(n_568) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_440), .B(n_750), .C(n_753), .D(n_756), .Y(n_749) );
NAND4xp25_ASAP7_75t_SL g948 ( .A(n_440), .B(n_949), .C(n_953), .D(n_956), .Y(n_948) );
NAND4xp25_ASAP7_75t_L g1223 ( .A(n_440), .B(n_1224), .C(n_1227), .D(n_1230), .Y(n_1223) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_442), .B(n_457), .C(n_466), .D(n_476), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_449), .C(n_455), .Y(n_442) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_445), .Y(n_459) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_445), .Y(n_588) );
BUFx2_ASAP7_75t_L g599 ( .A(n_445), .Y(n_599) );
INVx1_ASAP7_75t_L g718 ( .A(n_445), .Y(n_718) );
BUFx2_ASAP7_75t_L g966 ( .A(n_445), .Y(n_966) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g601 ( .A(n_448), .Y(n_601) );
INVx4_ASAP7_75t_L g649 ( .A(n_448), .Y(n_649) );
INVx2_ASAP7_75t_SL g968 ( .A(n_448), .Y(n_968) );
BUFx3_ASAP7_75t_L g970 ( .A(n_448), .Y(n_970) );
INVx2_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g524 ( .A(n_451), .Y(n_524) );
INVx2_ASAP7_75t_L g830 ( .A(n_451), .Y(n_830) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g463 ( .A(n_452), .Y(n_463) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_452), .Y(n_775) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g594 ( .A(n_453), .Y(n_594) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_454), .Y(n_485) );
INVx2_ASAP7_75t_SL g604 ( .A(n_454), .Y(n_604) );
AOI33xp33_ASAP7_75t_L g525 ( .A1(n_455), .A2(n_481), .A3(n_526), .B1(n_530), .B2(n_535), .B3(n_536), .Y(n_525) );
INVx2_ASAP7_75t_L g596 ( .A(n_455), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g715 ( .A(n_455), .B(n_716), .C(n_719), .Y(n_715) );
BUFx3_ASAP7_75t_L g772 ( .A(n_455), .Y(n_772) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_455), .B(n_832), .C(n_837), .Y(n_831) );
NAND3xp33_ASAP7_75t_L g908 ( .A(n_455), .B(n_909), .C(n_911), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g1234 ( .A(n_455), .B(n_1235), .C(n_1236), .Y(n_1234) );
INVx2_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx3_ASAP7_75t_L g777 ( .A(n_461), .Y(n_777) );
INVx2_ASAP7_75t_L g828 ( .A(n_461), .Y(n_828) );
INVx2_ASAP7_75t_L g910 ( .A(n_461), .Y(n_910) );
INVx2_ASAP7_75t_L g914 ( .A(n_461), .Y(n_914) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_464), .Y(n_817) );
AOI222xp33_ASAP7_75t_L g1216 ( .A1(n_464), .A2(n_564), .B1(n_684), .B2(n_1217), .C1(n_1218), .C2(n_1219), .Y(n_1216) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .C(n_475), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_SL g527 ( .A(n_469), .Y(n_527) );
HB1xp67_ASAP7_75t_L g958 ( .A(n_470), .Y(n_958) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_470), .Y(n_1228) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_SL g798 ( .A(n_473), .Y(n_798) );
INVx1_ASAP7_75t_L g789 ( .A(n_474), .Y(n_789) );
NAND3xp33_ASAP7_75t_L g841 ( .A(n_475), .B(n_842), .C(n_844), .Y(n_841) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_475), .B(n_917), .C(n_918), .Y(n_916) );
NAND3xp33_ASAP7_75t_L g1241 ( .A(n_475), .B(n_1242), .C(n_1243), .Y(n_1241) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .C(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND3xp33_ASAP7_75t_L g846 ( .A(n_481), .B(n_847), .C(n_848), .Y(n_846) );
INVx1_ASAP7_75t_L g875 ( .A(n_481), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g921 ( .A(n_481), .B(n_922), .C(n_923), .Y(n_921) );
NAND3xp33_ASAP7_75t_L g1244 ( .A(n_481), .B(n_1245), .C(n_1249), .Y(n_1244) );
INVx1_ASAP7_75t_L g564 ( .A(n_487), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_490), .A2(n_491), .B1(n_492), .B2(n_493), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_490), .A2(n_492), .B1(n_543), .B2(n_544), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_490), .A2(n_497), .B1(n_558), .B2(n_559), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_490), .A2(n_492), .B1(n_821), .B2(n_822), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_492), .A2(n_495), .B1(n_566), .B2(n_567), .Y(n_565) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_495), .A2(n_514), .B1(n_546), .B2(n_547), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_495), .A2(n_497), .B1(n_686), .B2(n_687), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_495), .A2(n_547), .B1(n_696), .B2(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_495), .A2(n_547), .B1(n_754), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_495), .A2(n_547), .B1(n_809), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_SL g988 ( .A1(n_495), .A2(n_497), .B1(n_954), .B2(n_989), .Y(n_988) );
AOI22xp5_ASAP7_75t_L g1220 ( .A1(n_495), .A2(n_497), .B1(n_1221), .B2(n_1222), .Y(n_1220) );
INVx1_ASAP7_75t_L g631 ( .A(n_499), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_551), .B2(n_552), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g550 ( .A(n_502), .Y(n_550) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_525), .Y(n_516) );
INVx1_ASAP7_75t_L g615 ( .A(n_519), .Y(n_615) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_L g894 ( .A(n_529), .Y(n_894) );
INVx2_ASAP7_75t_SL g625 ( .A(n_531), .Y(n_625) );
BUFx3_ASAP7_75t_L g787 ( .A(n_531), .Y(n_787) );
BUFx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g797 ( .A(n_533), .Y(n_797) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AOI31xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_542), .A3(n_545), .B(n_548), .Y(n_537) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
XNOR2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_554), .A2(n_1011), .B1(n_1016), .B2(n_1032), .Y(n_1031) );
BUFx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx4f_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g760 ( .A(n_579), .Y(n_760) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AO211x2_ASAP7_75t_L g690 ( .A1(n_582), .A2(n_691), .B(n_702), .C(n_714), .Y(n_690) );
BUFx6f_ASAP7_75t_L g961 ( .A(n_582), .Y(n_961) );
NAND4xp25_ASAP7_75t_L g583 ( .A(n_584), .B(n_597), .C(n_609), .D(n_621), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_591), .C(n_595), .Y(n_584) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_SL g721 ( .A(n_594), .Y(n_721) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_602), .C(n_605), .Y(n_597) );
INVxp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g782 ( .A(n_604), .Y(n_782) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_605), .B(n_657), .C(n_659), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_605), .B(n_724), .C(n_727), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g826 ( .A(n_605), .B(n_827), .C(n_829), .Y(n_826) );
INVx5_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx6_ASAP7_75t_L g783 ( .A(n_606), .Y(n_783) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_613), .C(n_618), .Y(n_609) );
BUFx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_615), .A2(n_872), .B1(n_873), .B2(n_874), .Y(n_871) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g678 ( .A(n_617), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g735 ( .A(n_619), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_619), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .C(n_626), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g794 ( .A(n_628), .Y(n_794) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_849), .B2(n_991), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
XNOR2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_744), .Y(n_634) );
XOR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_689), .Y(n_635) );
NAND3x1_ASAP7_75t_L g637 ( .A(n_638), .B(n_645), .C(n_680), .Y(n_637) );
AND4x1_ASAP7_75t_L g645 ( .A(n_646), .B(n_656), .C(n_660), .D(n_671), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_650), .C(n_654), .Y(n_646) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g840 ( .A(n_652), .Y(n_840) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
BUFx2_ASAP7_75t_L g722 ( .A(n_653), .Y(n_722) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI33xp33_ASAP7_75t_L g963 ( .A1(n_655), .A2(n_783), .A3(n_964), .B1(n_965), .B2(n_969), .B3(n_971), .Y(n_963) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_664), .C(n_669), .Y(n_660) );
INVx4_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g843 ( .A(n_663), .Y(n_843) );
INVx1_ASAP7_75t_L g1246 ( .A(n_663), .Y(n_1246) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
OAI33xp33_ASAP7_75t_L g855 ( .A1(n_670), .A2(n_856), .A3(n_861), .B1(n_868), .B2(n_871), .B3(n_875), .Y(n_855) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_675), .C(n_679), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g977 ( .A(n_677), .Y(n_977) );
AOI33xp33_ASAP7_75t_L g975 ( .A1(n_679), .A2(n_785), .A3(n_976), .B1(n_978), .B2(n_979), .B3(n_980), .Y(n_975) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_715), .B(n_723), .C(n_728), .D(n_736), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
BUFx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g839 ( .A(n_721), .Y(n_839) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_732), .C(n_735), .Y(n_728) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
BUFx4f_ASAP7_75t_L g740 ( .A(n_733), .Y(n_740) );
INVx1_ASAP7_75t_L g858 ( .A(n_733), .Y(n_858) );
NAND3xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_739), .C(n_743), .Y(n_736) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_801), .B2(n_802), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g800 ( .A(n_748), .Y(n_800) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_784), .Y(n_770) );
AOI33xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .A3(n_776), .B1(n_778), .B2(n_781), .B3(n_783), .Y(n_771) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g912 ( .A(n_783), .B(n_913), .C(n_915), .Y(n_912) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND3xp33_ASAP7_75t_L g815 ( .A(n_816), .B(n_820), .C(n_823), .Y(n_815) );
NAND4xp25_ASAP7_75t_L g825 ( .A(n_826), .B(n_831), .C(n_841), .D(n_846), .Y(n_825) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g991 ( .A(n_849), .Y(n_991) );
XNOR2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_902), .Y(n_849) );
INVx2_ASAP7_75t_SL g850 ( .A(n_851), .Y(n_850) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND3xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_889), .C(n_897), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_876), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .B1(n_859), .B2(n_860), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B1(n_865), .B2(n_866), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_863), .A2(n_866), .B1(n_869), .B2(n_870), .Y(n_868) );
INVx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
OAI22xp33_ASAP7_75t_L g885 ( .A1(n_878), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_885) );
INVx2_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g1256 ( .A(n_887), .Y(n_1256) );
AOI22xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .B1(n_946), .B2(n_990), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
XOR2xp5_ASAP7_75t_L g905 ( .A(n_906), .B(n_945), .Y(n_905) );
NAND3xp33_ASAP7_75t_L g906 ( .A(n_907), .B(n_925), .C(n_935), .Y(n_906) );
AND4x1_ASAP7_75t_L g907 ( .A(n_908), .B(n_912), .C(n_916), .D(n_921), .Y(n_907) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx2_ASAP7_75t_SL g990 ( .A(n_946), .Y(n_990) );
AOI211xp5_ASAP7_75t_SL g947 ( .A1(n_948), .A2(n_961), .B(n_962), .C(n_981), .Y(n_947) );
OAI31xp33_ASAP7_75t_L g1261 ( .A1(n_961), .A2(n_1262), .A3(n_1263), .B(n_1267), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_963), .B(n_975), .Y(n_962) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
OAI21xp33_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_1206), .B(n_1208), .Y(n_992) );
NOR2x1_ASAP7_75t_L g993 ( .A(n_994), .B(n_1172), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_1123), .Y(n_994) );
NOR4xp25_ASAP7_75t_L g995 ( .A(n_996), .B(n_1065), .C(n_1085), .D(n_1101), .Y(n_995) );
AOI21xp33_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_1049), .B(n_1053), .Y(n_996) );
OR2x2_ASAP7_75t_L g997 ( .A(n_998), .B(n_1018), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_998), .B(n_1050), .Y(n_1129) );
INVx1_ASAP7_75t_L g1167 ( .A(n_998), .Y(n_1167) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1127 ( .A(n_999), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_999), .B(n_1131), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_999), .B(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1197 ( .A(n_999), .Y(n_1197) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1000), .B(n_1072), .Y(n_1071) );
INVx2_ASAP7_75t_SL g1084 ( .A(n_1000), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1099 ( .A(n_1000), .B(n_1072), .Y(n_1099) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1001), .Y(n_1063) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1001), .Y(n_1116) );
AND2x4_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1005), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_1002), .B(n_1005), .Y(n_1029) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_1003), .B(n_1005), .Y(n_1007) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_1004), .B(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1006), .Y(n_1014) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1007), .Y(n_1038) );
INVx1_ASAP7_75t_SL g1044 ( .A(n_1007), .Y(n_1044) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1010), .B1(n_1015), .B2(n_1016), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_1010), .A2(n_1016), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
OAI22xp33_ASAP7_75t_L g1056 ( .A1(n_1010), .A2(n_1057), .B1(n_1058), .B2(n_1059), .Y(n_1056) );
BUFx3_ASAP7_75t_L g1120 ( .A(n_1010), .Y(n_1120) );
BUFx6f_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1013), .Y(n_1011) );
OR2x2_ASAP7_75t_L g1016 ( .A(n_1012), .B(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1012), .Y(n_1025) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1013), .Y(n_1024) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1016), .Y(n_1060) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1017), .Y(n_1027) );
A2O1A1Ixp33_ASAP7_75t_L g1065 ( .A1(n_1018), .A2(n_1066), .B(n_1070), .C(n_1075), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1033), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1019), .B(n_1069), .Y(n_1068) );
OAI21xp5_ASAP7_75t_L g1094 ( .A1(n_1019), .A2(n_1095), .B(n_1096), .Y(n_1094) );
NAND3xp33_ASAP7_75t_L g1149 ( .A(n_1019), .B(n_1107), .C(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1156 ( .A(n_1020), .B(n_1034), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1020), .B(n_1040), .Y(n_1177) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1030), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1021), .B(n_1030), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1021), .B(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1021), .Y(n_1089) );
O2A1O1Ixp33_ASAP7_75t_SL g1101 ( .A1(n_1021), .A2(n_1102), .B(n_1105), .C(n_1112), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1021), .B(n_1040), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1028), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .Y(n_1023) );
AND2x4_ASAP7_75t_L g1026 ( .A(n_1025), .B(n_1027), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1281 ( .A(n_1027), .Y(n_1281) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1029), .Y(n_1042) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1030), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1030), .B(n_1039), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1030), .B(n_1089), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1030), .B(n_1033), .Y(n_1128) );
AOI32xp33_ASAP7_75t_L g1159 ( .A1(n_1030), .A2(n_1091), .A3(n_1143), .B1(n_1160), .B2(n_1161), .Y(n_1159) );
A2O1A1Ixp33_ASAP7_75t_L g1163 ( .A1(n_1030), .A2(n_1034), .B(n_1098), .C(n_1133), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1033), .B(n_1052), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1039), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1034), .B(n_1052), .Y(n_1051) );
NOR2xp33_ASAP7_75t_L g1069 ( .A(n_1034), .B(n_1039), .Y(n_1069) );
INVx2_ASAP7_75t_L g1080 ( .A(n_1034), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1034), .B(n_1055), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1034), .B(n_1104), .Y(n_1103) );
INVx4_ASAP7_75t_L g1141 ( .A(n_1034), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1144 ( .A(n_1034), .B(n_1145), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1034), .B(n_1146), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1034), .B(n_1177), .Y(n_1200) );
AND2x6_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
INVx2_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g1114 ( .A1(n_1038), .A2(n_1115), .B1(n_1116), .B2(n_1117), .Y(n_1114) );
NOR2xp33_ASAP7_75t_L g1050 ( .A(n_1039), .B(n_1051), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1039), .B(n_1077), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1135 ( .A(n_1039), .B(n_1078), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1039), .B(n_1111), .Y(n_1169) );
CKINVDCx6p67_ASAP7_75t_R g1039 ( .A(n_1040), .Y(n_1039) );
OR2x2_ASAP7_75t_L g1088 ( .A(n_1040), .B(n_1089), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1040), .B(n_1089), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1040), .B(n_1077), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1040), .B(n_1111), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1040), .B(n_1052), .Y(n_1154) );
OAI211xp5_ASAP7_75t_SL g1158 ( .A1(n_1040), .A2(n_1086), .B(n_1159), .C(n_1163), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1040), .B(n_1166), .Y(n_1165) );
OR2x6_ASAP7_75t_SL g1040 ( .A(n_1041), .B(n_1046), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_1042), .A2(n_1043), .B1(n_1044), .B2(n_1045), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_1044), .A2(n_1062), .B1(n_1063), .B2(n_1064), .Y(n_1061) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1052), .B(n_1141), .Y(n_1166) );
INVx1_ASAP7_75t_SL g1143 ( .A(n_1053), .Y(n_1143) );
INVx3_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1054), .Y(n_1087) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_1054), .B(n_1072), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1054), .B(n_1113), .Y(n_1112) );
OAI211xp5_ASAP7_75t_L g1124 ( .A1(n_1054), .A2(n_1125), .B(n_1129), .C(n_1130), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1054), .B(n_1071), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1054), .B(n_1084), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1054), .B(n_1107), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1054), .B(n_1146), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1054), .B(n_1072), .Y(n_1201) );
INVx3_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1055), .B(n_1072), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1204 ( .A(n_1055), .B(n_1099), .Y(n_1204) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1061), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_1059), .Y(n_1122) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
NOR2xp33_ASAP7_75t_L g1196 ( .A(n_1068), .B(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
AOI221xp5_ASAP7_75t_L g1138 ( .A1(n_1071), .A2(n_1139), .B1(n_1142), .B2(n_1147), .C(n_1148), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1071), .B(n_1140), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_1071), .A2(n_1174), .B1(n_1180), .B2(n_1183), .Y(n_1173) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_1072), .B(n_1084), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1072), .B(n_1084), .Y(n_1104) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1072), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1074), .Y(n_1072) );
OAI21xp5_ASAP7_75t_L g1075 ( .A1(n_1076), .A2(n_1079), .B(n_1082), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_1076), .A2(n_1132), .B1(n_1141), .B2(n_1169), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1076), .B(n_1141), .Y(n_1194) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1077), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1077), .B(n_1140), .Y(n_1139) );
O2A1O1Ixp33_ASAP7_75t_L g1195 ( .A1(n_1079), .A2(n_1126), .B(n_1187), .C(n_1196), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1081), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1080), .B(n_1092), .Y(n_1091) );
NOR2xp33_ASAP7_75t_L g1106 ( .A(n_1080), .B(n_1107), .Y(n_1106) );
INVx2_ASAP7_75t_L g1132 ( .A(n_1080), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1082), .B(n_1087), .Y(n_1086) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx2_ASAP7_75t_SL g1146 ( .A(n_1084), .Y(n_1146) );
OAI221xp5_ASAP7_75t_L g1085 ( .A1(n_1086), .A2(n_1088), .B1(n_1090), .B2(n_1093), .C(n_1094), .Y(n_1085) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1088), .Y(n_1092) );
OAI211xp5_ASAP7_75t_SL g1148 ( .A1(n_1088), .A2(n_1093), .B(n_1149), .C(n_1152), .Y(n_1148) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1100), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1098), .B(n_1141), .Y(n_1183) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_1099), .A2(n_1126), .B1(n_1127), .B2(n_1128), .Y(n_1125) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1104), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1108), .Y(n_1105) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1107), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .Y(n_1108) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
CKINVDCx5p33_ASAP7_75t_R g1152 ( .A(n_1113), .Y(n_1152) );
OR2x6_ASAP7_75t_SL g1113 ( .A(n_1114), .B(n_1118), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_1119), .A2(n_1120), .B1(n_1121), .B2(n_1122), .Y(n_1118) );
BUFx2_ASAP7_75t_SL g1207 ( .A(n_1122), .Y(n_1207) );
OAI32xp33_ASAP7_75t_L g1123 ( .A1(n_1124), .A2(n_1134), .A3(n_1152), .B1(n_1158), .B2(n_1164), .Y(n_1123) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1126), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1133), .Y(n_1131) );
OAI211xp5_ASAP7_75t_SL g1134 ( .A1(n_1135), .A2(n_1136), .B(n_1138), .C(n_1153), .Y(n_1134) );
OAI21xp33_ASAP7_75t_L g1199 ( .A1(n_1135), .A2(n_1141), .B(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1137), .B(n_1154), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1140), .B(n_1147), .Y(n_1203) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
NOR2xp33_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1144), .Y(n_1142) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1144), .Y(n_1188) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
A2O1A1Ixp33_ASAP7_75t_SL g1172 ( .A1(n_1152), .A2(n_1173), .B(n_1184), .C(n_1198), .Y(n_1172) );
OAI21xp5_ASAP7_75t_L g1153 ( .A1(n_1154), .A2(n_1155), .B(n_1157), .Y(n_1153) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
A2O1A1Ixp33_ASAP7_75t_L g1202 ( .A1(n_1156), .A2(n_1203), .B(n_1204), .C(n_1205), .Y(n_1202) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
O2A1O1Ixp33_ASAP7_75t_SL g1164 ( .A1(n_1165), .A2(n_1167), .B(n_1168), .C(n_1170), .Y(n_1164) );
O2A1O1Ixp33_ASAP7_75t_L g1184 ( .A1(n_1169), .A2(n_1185), .B(n_1188), .C(n_1189), .Y(n_1184) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
NOR2xp33_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1178), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
NOR2xp33_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1182), .Y(n_1180) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
A2O1A1Ixp33_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1191), .B(n_1193), .C(n_1195), .Y(n_1189) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
AOI21xp5_ASAP7_75t_L g1198 ( .A1(n_1199), .A2(n_1201), .B(n_1202), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
HB1xp67_ASAP7_75t_L g1275 ( .A(n_1211), .Y(n_1275) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1213), .Y(n_1260) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1220), .Y(n_1253) );
INVxp67_ASAP7_75t_L g1262 ( .A(n_1224), .Y(n_1262) );
INVxp67_ASAP7_75t_L g1267 ( .A(n_1230), .Y(n_1267) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
NAND3xp33_ASAP7_75t_L g1251 ( .A(n_1233), .B(n_1252), .C(n_1261), .Y(n_1251) );
AND4x1_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1237), .C(n_1241), .D(n_1244), .Y(n_1233) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
BUFx2_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
CKINVDCx5p33_ASAP7_75t_R g1277 ( .A(n_1278), .Y(n_1277) );
OAI21xp5_ASAP7_75t_L g1280 ( .A1(n_1279), .A2(n_1281), .B(n_1282), .Y(n_1280) );
endmodule