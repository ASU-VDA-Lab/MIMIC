module fake_aes_8580_n_853 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_853);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_853;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_165;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_522;
wire n_264;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_836;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_44), .Y(n_103) );
BUFx8_ASAP7_75t_SL g104 ( .A(n_76), .Y(n_104) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_33), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_35), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_51), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_89), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_19), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_67), .Y(n_110) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_32), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_101), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_102), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_96), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_97), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_78), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_3), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_48), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_68), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_61), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_4), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_100), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_5), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_27), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_79), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_39), .Y(n_126) );
INVx2_ASAP7_75t_SL g127 ( .A(n_99), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_73), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_13), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_60), .Y(n_130) );
BUFx3_ASAP7_75t_L g131 ( .A(n_70), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_64), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_42), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_58), .Y(n_134) );
INVx2_ASAP7_75t_SL g135 ( .A(n_43), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_2), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_52), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_25), .Y(n_138) );
CKINVDCx16_ASAP7_75t_R g139 ( .A(n_46), .Y(n_139) );
BUFx10_ASAP7_75t_L g140 ( .A(n_26), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_27), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_32), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_57), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_47), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_34), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_36), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_106), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_111), .B(n_0), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_127), .B(n_0), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_104), .Y(n_151) );
INVx2_ASAP7_75t_SL g152 ( .A(n_112), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_106), .Y(n_153) );
BUFx12f_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
INVx5_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_135), .B(n_1), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_117), .B(n_1), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_112), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_111), .Y(n_159) );
INVx2_ASAP7_75t_SL g160 ( .A(n_131), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_117), .B(n_2), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_119), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_135), .B(n_3), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_131), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_131), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_119), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_135), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_104), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_119), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_150), .A2(n_139), .B1(n_123), .B2(n_138), .Y(n_170) );
OAI22xp33_ASAP7_75t_L g171 ( .A1(n_168), .A2(n_123), .B1(n_145), .B2(n_126), .Y(n_171) );
OAI22xp33_ASAP7_75t_L g172 ( .A1(n_168), .A2(n_145), .B1(n_126), .B2(n_129), .Y(n_172) );
OAI22xp5_ASAP7_75t_SL g173 ( .A1(n_151), .A2(n_109), .B1(n_144), .B2(n_124), .Y(n_173) );
INVx8_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_150), .B(n_139), .Y(n_175) );
OR2x6_ASAP7_75t_L g176 ( .A(n_168), .B(n_129), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_159), .B(n_140), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_159), .B(n_149), .Y(n_178) );
OAI22xp33_ASAP7_75t_SL g179 ( .A1(n_157), .A2(n_146), .B1(n_142), .B2(n_141), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_150), .A2(n_121), .B1(n_106), .B2(n_136), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_150), .B(n_136), .Y(n_182) );
BUFx10_ASAP7_75t_L g183 ( .A(n_150), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_149), .B(n_140), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_150), .A2(n_136), .B1(n_140), .B2(n_105), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_150), .A2(n_140), .B1(n_105), .B2(n_137), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_156), .A2(n_105), .B1(n_137), .B2(n_114), .Y(n_187) );
OAI22xp33_ASAP7_75t_R g188 ( .A1(n_163), .A2(n_114), .B1(n_115), .B2(n_122), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_155), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_148), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g191 ( .A1(n_151), .A2(n_115), .B1(n_133), .B2(n_122), .Y(n_191) );
OA22x2_ASAP7_75t_L g192 ( .A1(n_156), .A2(n_128), .B1(n_130), .B2(n_133), .Y(n_192) );
AND2x2_ASAP7_75t_SL g193 ( .A(n_156), .B(n_128), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_157), .A2(n_105), .B1(n_130), .B2(n_132), .Y(n_194) );
OAI22xp33_ASAP7_75t_L g195 ( .A1(n_157), .A2(n_105), .B1(n_134), .B2(n_125), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_148), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_149), .A2(n_156), .B1(n_163), .B2(n_161), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_149), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_156), .B(n_105), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_148), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_156), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
AOI22xp5_ASAP7_75t_SL g203 ( .A1(n_161), .A2(n_143), .B1(n_120), .B2(n_118), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_156), .B(n_105), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_155), .Y(n_207) );
INVx1_ASAP7_75t_SL g208 ( .A(n_161), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_152), .B(n_160), .Y(n_210) );
NAND3xp33_ASAP7_75t_L g211 ( .A(n_148), .B(n_116), .C(n_113), .Y(n_211) );
OAI22xp33_ASAP7_75t_SL g212 ( .A1(n_147), .A2(n_110), .B1(n_108), .B2(n_107), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_154), .B(n_103), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_154), .B(n_155), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_154), .B(n_40), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_208), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_184), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_184), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_177), .B(n_154), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_206), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_206), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_204), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_201), .Y(n_223) );
INVx4_ASAP7_75t_SL g224 ( .A(n_199), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_204), .Y(n_225) );
XOR2xp5_ASAP7_75t_L g226 ( .A(n_173), .B(n_4), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_176), .B(n_152), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_205), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_205), .Y(n_229) );
XOR2xp5_ASAP7_75t_L g230 ( .A(n_198), .B(n_5), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_209), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_174), .B(n_155), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_201), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_174), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_177), .B(n_155), .Y(n_235) );
INVxp33_ASAP7_75t_SL g236 ( .A(n_203), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_178), .B(n_152), .Y(n_237) );
NAND2xp33_ASAP7_75t_SL g238 ( .A(n_198), .B(n_152), .Y(n_238) );
AND2x6_ASAP7_75t_L g239 ( .A(n_201), .B(n_148), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_209), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_170), .B(n_181), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_199), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_199), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_182), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_178), .B(n_155), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_175), .B(n_155), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_175), .B(n_155), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_183), .Y(n_248) );
NOR2xp33_ASAP7_75t_SL g249 ( .A(n_174), .B(n_155), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_197), .B(n_193), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_213), .B(n_155), .Y(n_251) );
XNOR2x2_ASAP7_75t_L g252 ( .A(n_192), .B(n_147), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_176), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_176), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_176), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_210), .A2(n_160), .B(n_167), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_182), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_171), .B(n_147), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_210), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_192), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_192), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_183), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_193), .Y(n_265) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_215), .B(n_167), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_212), .B(n_167), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_185), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_186), .Y(n_270) );
BUFx5_ASAP7_75t_L g271 ( .A(n_174), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_187), .A2(n_160), .B(n_167), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_188), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_188), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_191), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_194), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_179), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_222), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_250), .B(n_172), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_216), .B(n_267), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_225), .Y(n_281) );
AND2x2_ASAP7_75t_SL g282 ( .A(n_227), .B(n_214), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_271), .B(n_160), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_219), .B(n_195), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_228), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_229), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_231), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_240), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_271), .B(n_217), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_253), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_218), .B(n_189), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_265), .B(n_189), .Y(n_292) );
NOR2xp67_ASAP7_75t_R g293 ( .A(n_262), .B(n_167), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_261), .B(n_207), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_241), .B(n_207), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_271), .B(n_167), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_263), .B(n_167), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_223), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_223), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_271), .B(n_167), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_233), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_271), .B(n_167), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_271), .B(n_167), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_271), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_237), .B(n_167), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_239), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_233), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_242), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_239), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_237), .B(n_202), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_245), .B(n_202), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_243), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_227), .B(n_153), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_220), .B(n_202), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_239), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_254), .B(n_162), .Y(n_316) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_227), .B(n_162), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_224), .B(n_221), .Y(n_318) );
OAI21xp5_ASAP7_75t_L g319 ( .A1(n_246), .A2(n_200), .B(n_196), .Y(n_319) );
AND2x2_ASAP7_75t_SL g320 ( .A(n_247), .B(n_169), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_253), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_254), .B(n_169), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_239), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_244), .B(n_169), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_270), .A2(n_200), .B(n_196), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_234), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_248), .B(n_211), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_234), .Y(n_328) );
BUFx4f_ASAP7_75t_L g329 ( .A(n_317), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_278), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
BUFx12f_ASAP7_75t_L g332 ( .A(n_290), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_280), .B(n_273), .Y(n_333) );
NAND2x1_ASAP7_75t_L g334 ( .A(n_278), .B(n_239), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_278), .Y(n_336) );
INVx4_ASAP7_75t_SL g337 ( .A(n_304), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_278), .Y(n_338) );
AND2x6_ASAP7_75t_L g339 ( .A(n_304), .B(n_255), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_317), .B(n_256), .Y(n_340) );
NAND2x1p5_ASAP7_75t_L g341 ( .A(n_304), .B(n_259), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_317), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_280), .B(n_274), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_317), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_313), .B(n_277), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_279), .B(n_256), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_317), .B(n_280), .Y(n_347) );
BUFx6f_ASAP7_75t_SL g348 ( .A(n_317), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_278), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_279), .B(n_260), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_281), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_280), .B(n_248), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_281), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_281), .B(n_258), .Y(n_354) );
OR2x6_ASAP7_75t_L g355 ( .A(n_313), .B(n_257), .Y(n_355) );
OR2x6_ASAP7_75t_L g356 ( .A(n_313), .B(n_232), .Y(n_356) );
INVx5_ASAP7_75t_L g357 ( .A(n_306), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_281), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_281), .Y(n_359) );
AND2x6_ASAP7_75t_L g360 ( .A(n_326), .B(n_269), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_329), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_335), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_330), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_348), .A2(n_282), .B1(n_238), .B2(n_279), .Y(n_364) );
CKINVDCx8_ASAP7_75t_R g365 ( .A(n_342), .Y(n_365) );
BUFx4_ASAP7_75t_SL g366 ( .A(n_330), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_329), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_349), .B(n_285), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_335), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_329), .B(n_288), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_332), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_335), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
CKINVDCx14_ASAP7_75t_R g374 ( .A(n_332), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_349), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_329), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_336), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_336), .Y(n_379) );
BUFx8_ASAP7_75t_L g380 ( .A(n_348), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_332), .Y(n_381) );
BUFx12f_ASAP7_75t_L g382 ( .A(n_342), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_339), .Y(n_383) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_336), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_353), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_339), .Y(n_387) );
BUFx5_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
BUFx4f_ASAP7_75t_SL g389 ( .A(n_339), .Y(n_389) );
AOI22xp33_ASAP7_75t_SL g390 ( .A1(n_389), .A2(n_348), .B1(n_344), .B2(n_347), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_389), .A2(n_348), .B1(n_380), .B2(n_344), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_363), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_388), .B(n_333), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_366), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_363), .Y(n_397) );
CKINVDCx6p67_ASAP7_75t_R g398 ( .A(n_371), .Y(n_398) );
INVx6_ASAP7_75t_L g399 ( .A(n_380), .Y(n_399) );
CKINVDCx11_ASAP7_75t_R g400 ( .A(n_371), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_388), .A2(n_348), .B1(n_342), .B2(n_346), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_388), .A2(n_342), .B1(n_346), .B2(n_345), .Y(n_402) );
INVx6_ASAP7_75t_L g403 ( .A(n_380), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_388), .Y(n_404) );
INVx6_ASAP7_75t_L g405 ( .A(n_380), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_381), .Y(n_406) );
BUFx10_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_364), .A2(n_342), .B1(n_355), .B2(n_346), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_376), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_389), .A2(n_347), .B1(n_342), .B2(n_340), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_388), .A2(n_342), .B1(n_345), .B2(n_347), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_378), .Y(n_412) );
OAI21xp5_ASAP7_75t_SL g413 ( .A1(n_364), .A2(n_226), .B(n_230), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_388), .B(n_353), .Y(n_414) );
BUFx10_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_388), .A2(n_345), .B1(n_333), .B2(n_343), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_388), .A2(n_345), .B1(n_343), .B2(n_236), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_376), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_374), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_381), .Y(n_420) );
AOI22xp33_ASAP7_75t_SL g421 ( .A1(n_380), .A2(n_340), .B1(n_236), .B2(n_290), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_364), .A2(n_355), .B1(n_345), .B2(n_282), .Y(n_422) );
CKINVDCx11_ASAP7_75t_R g423 ( .A(n_374), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_376), .A2(n_355), .B1(n_345), .B2(n_282), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_380), .A2(n_340), .B1(n_360), .B2(n_321), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_388), .A2(n_370), .B1(n_377), .B2(n_380), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_384), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_385), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_388), .B(n_338), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_388), .B(n_350), .Y(n_430) );
CKINVDCx11_ASAP7_75t_R g431 ( .A(n_382), .Y(n_431) );
OAI21xp5_ASAP7_75t_SL g432 ( .A1(n_370), .A2(n_226), .B(n_230), .Y(n_432) );
BUFx12f_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_396), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_422), .A2(n_388), .B1(n_377), .B2(n_373), .Y(n_435) );
BUFx4f_ASAP7_75t_SL g436 ( .A(n_406), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_427), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_429), .B(n_384), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_394), .A2(n_387), .B1(n_386), .B2(n_383), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_424), .A2(n_388), .B1(n_377), .B2(n_373), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_408), .A2(n_388), .B1(n_377), .B2(n_373), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_423), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_400), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_428), .Y(n_444) );
CKINVDCx11_ASAP7_75t_R g445 ( .A(n_406), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_428), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_407), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_425), .A2(n_388), .B1(n_373), .B2(n_367), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_429), .B(n_384), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_427), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_394), .A2(n_387), .B1(n_386), .B2(n_383), .Y(n_451) );
NOR2x1_ASAP7_75t_SL g452 ( .A(n_433), .B(n_383), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_392), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_392), .Y(n_454) );
OR2x2_ASAP7_75t_SL g455 ( .A(n_399), .B(n_385), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_412), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_433), .A2(n_388), .B1(n_367), .B2(n_373), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_398), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_397), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_395), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_395), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_413), .A2(n_383), .B1(n_387), .B2(n_386), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_404), .A2(n_388), .B1(n_361), .B2(n_367), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_409), .Y(n_464) );
OAI211xp5_ASAP7_75t_L g465 ( .A1(n_432), .A2(n_321), .B(n_275), .C(n_260), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_414), .B(n_378), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_404), .A2(n_388), .B1(n_367), .B2(n_361), .Y(n_467) );
OAI21xp5_ASAP7_75t_SL g468 ( .A1(n_421), .A2(n_370), .B(n_321), .Y(n_468) );
OAI21xp33_ASAP7_75t_L g469 ( .A1(n_409), .A2(n_418), .B(n_417), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_412), .B(n_369), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_399), .A2(n_387), .B1(n_386), .B2(n_383), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_414), .B(n_385), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_416), .A2(n_387), .B1(n_386), .B2(n_355), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_419), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_396), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_399), .A2(n_361), .B1(n_367), .B2(n_370), .Y(n_477) );
BUFx3_ASAP7_75t_L g478 ( .A(n_407), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_396), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_396), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_430), .B(n_350), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_396), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_426), .B(n_378), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_399), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g485 ( .A1(n_403), .A2(n_382), .B1(n_361), .B2(n_360), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_403), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_407), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_403), .A2(n_361), .B1(n_355), .B2(n_360), .Y(n_488) );
INVx5_ASAP7_75t_SL g489 ( .A(n_398), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_403), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_405), .A2(n_355), .B1(n_360), .B2(n_356), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_405), .A2(n_360), .B1(n_356), .B2(n_350), .Y(n_492) );
BUFx12f_ASAP7_75t_L g493 ( .A(n_415), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_405), .A2(n_360), .B1(n_356), .B2(n_339), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_401), .A2(n_368), .B1(n_365), .B2(n_356), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_405), .A2(n_360), .B1(n_356), .B2(n_339), .Y(n_496) );
BUFx12f_ASAP7_75t_L g497 ( .A(n_415), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_393), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_402), .A2(n_368), .B1(n_365), .B2(n_356), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_391), .A2(n_368), .B1(n_365), .B2(n_351), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_415), .A2(n_352), .B1(n_360), .B2(n_275), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_431), .A2(n_360), .B1(n_339), .B2(n_382), .Y(n_502) );
NOR2x1_ASAP7_75t_SL g503 ( .A(n_390), .B(n_382), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_411), .A2(n_365), .B1(n_351), .B2(n_358), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_410), .B(n_378), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_420), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_462), .A2(n_360), .B1(n_382), .B2(n_339), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_435), .A2(n_339), .B1(n_238), .B2(n_352), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_468), .A2(n_365), .B1(n_379), .B2(n_378), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_503), .A2(n_419), .B1(n_369), .B2(n_375), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_503), .A2(n_375), .B1(n_372), .B2(n_369), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_474), .A2(n_339), .B1(n_341), .B2(n_331), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_440), .A2(n_341), .B1(n_331), .B2(n_320), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_444), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_499), .A2(n_341), .B1(n_331), .B2(n_320), .Y(n_515) );
AOI21xp33_ASAP7_75t_L g516 ( .A1(n_465), .A2(n_169), .B(n_268), .Y(n_516) );
AOI22xp33_ASAP7_75t_SL g517 ( .A1(n_452), .A2(n_375), .B1(n_372), .B2(n_369), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_495), .A2(n_341), .B1(n_331), .B2(n_320), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_492), .A2(n_331), .B1(n_320), .B2(n_359), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_501), .A2(n_320), .B1(n_338), .B2(n_351), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_468), .A2(n_322), .B1(n_316), .B2(n_358), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_501), .A2(n_320), .B1(n_358), .B2(n_338), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_491), .A2(n_359), .B1(n_322), .B2(n_316), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_469), .A2(n_316), .B1(n_322), .B2(n_359), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_469), .A2(n_316), .B1(n_322), .B2(n_354), .Y(n_525) );
OAI222xp33_ASAP7_75t_L g526 ( .A1(n_485), .A2(n_379), .B1(n_375), .B2(n_372), .C1(n_369), .C2(n_334), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_498), .A2(n_335), .B1(n_375), .B2(n_372), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_455), .A2(n_379), .B1(n_375), .B2(n_372), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_498), .A2(n_335), .B1(n_375), .B2(n_372), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_498), .A2(n_335), .B1(n_372), .B2(n_369), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_506), .A2(n_369), .B1(n_362), .B2(n_252), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_506), .A2(n_362), .B1(n_252), .B2(n_318), .Y(n_532) );
AOI222xp33_ASAP7_75t_L g533 ( .A1(n_436), .A2(n_337), .B1(n_153), .B2(n_379), .C1(n_313), .C2(n_287), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_455), .A2(n_379), .B1(n_282), .B2(n_362), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_466), .B(n_362), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_506), .A2(n_362), .B1(n_318), .B2(n_337), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_452), .A2(n_362), .B1(n_282), .B2(n_313), .Y(n_537) );
NAND3xp33_ASAP7_75t_SL g538 ( .A(n_458), .B(n_153), .C(n_169), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_441), .A2(n_362), .B1(n_318), .B2(n_337), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g540 ( .A1(n_444), .A2(n_295), .B1(n_166), .B2(n_318), .C(n_313), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_483), .A2(n_362), .B1(n_318), .B2(n_337), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_483), .A2(n_362), .B1(n_318), .B2(n_337), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_502), .A2(n_282), .B1(n_362), .B2(n_288), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_500), .A2(n_318), .B1(n_337), .B2(n_313), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_488), .A2(n_318), .B1(n_313), .B2(n_288), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_489), .A2(n_357), .B1(n_354), .B2(n_289), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_484), .A2(n_288), .B1(n_295), .B2(n_285), .Y(n_547) );
AOI221xp5_ASAP7_75t_SL g548 ( .A1(n_446), .A2(n_166), .B1(n_295), .B2(n_148), .C(n_165), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_438), .B(n_148), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_484), .A2(n_288), .B1(n_286), .B2(n_285), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g551 ( .A(n_459), .B(n_166), .C(n_158), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_484), .A2(n_287), .B1(n_286), .B2(n_354), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_481), .A2(n_287), .B1(n_286), .B2(n_289), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_484), .A2(n_284), .B1(n_166), .B2(n_334), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_494), .A2(n_284), .B1(n_166), .B2(n_276), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_466), .B(n_6), .Y(n_556) );
OAI21xp5_ASAP7_75t_SL g557 ( .A1(n_472), .A2(n_326), .B(n_289), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_496), .A2(n_284), .B1(n_166), .B2(n_289), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_438), .B(n_148), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_473), .B(n_6), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_493), .A2(n_166), .B1(n_357), .B2(n_148), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_489), .A2(n_457), .B1(n_448), .B2(n_477), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_446), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_470), .B(n_166), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_489), .A2(n_326), .B1(n_294), .B2(n_298), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_478), .Y(n_566) );
AOI22xp33_ASAP7_75t_SL g567 ( .A1(n_489), .A2(n_357), .B1(n_283), .B2(n_328), .Y(n_567) );
OAI211xp5_ASAP7_75t_L g568 ( .A1(n_445), .A2(n_324), .B(n_166), .C(n_294), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_453), .B(n_7), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_493), .A2(n_166), .B1(n_357), .B2(n_158), .Y(n_570) );
OAI222xp33_ASAP7_75t_L g571 ( .A1(n_447), .A2(n_324), .B1(n_357), .B2(n_283), .C1(n_294), .C2(n_328), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_497), .A2(n_357), .B1(n_158), .B2(n_164), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_497), .A2(n_357), .B1(n_158), .B2(n_164), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_505), .A2(n_357), .B1(n_158), .B2(n_164), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_478), .B(n_158), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_453), .B(n_158), .C(n_165), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_449), .B(n_158), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_505), .A2(n_158), .B1(n_164), .B2(n_165), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_454), .A2(n_158), .B1(n_165), .B2(n_164), .C(n_324), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_449), .B(n_454), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_478), .A2(n_328), .B1(n_291), .B2(n_301), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g582 ( .A1(n_489), .A2(n_283), .B1(n_165), .B2(n_164), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_463), .A2(n_301), .B1(n_299), .B2(n_307), .Y(n_583) );
OAI222xp33_ASAP7_75t_L g584 ( .A1(n_447), .A2(n_7), .B1(n_8), .B2(n_9), .C1(n_10), .C2(n_11), .Y(n_584) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_486), .A2(n_164), .B1(n_165), .B2(n_235), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_467), .A2(n_301), .B1(n_298), .B2(n_299), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_475), .B(n_8), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_487), .A2(n_301), .B1(n_298), .B2(n_299), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_460), .B(n_164), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_490), .A2(n_165), .B1(n_312), .B2(n_299), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_487), .A2(n_165), .B1(n_315), .B2(n_306), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_490), .A2(n_312), .B1(n_298), .B2(n_301), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_439), .A2(n_312), .B1(n_298), .B2(n_307), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_451), .A2(n_306), .B1(n_315), .B2(n_307), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_437), .A2(n_307), .B1(n_291), .B2(n_305), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_461), .A2(n_308), .B1(n_327), .B2(n_319), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_461), .A2(n_308), .B1(n_327), .B2(n_319), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_464), .A2(n_327), .B1(n_319), .B2(n_325), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_471), .A2(n_325), .B1(n_291), .B2(n_266), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_471), .A2(n_325), .B1(n_266), .B2(n_323), .Y(n_600) );
NAND3xp33_ASAP7_75t_L g601 ( .A(n_476), .B(n_180), .C(n_190), .Y(n_601) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_437), .A2(n_305), .B1(n_323), .B2(n_309), .Y(n_602) );
OA21x2_ASAP7_75t_L g603 ( .A1(n_548), .A2(n_476), .B(n_482), .Y(n_603) );
NOR3xp33_ASAP7_75t_L g604 ( .A(n_584), .B(n_442), .C(n_504), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_580), .B(n_450), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_549), .B(n_559), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_557), .A2(n_450), .B1(n_479), .B2(n_482), .C(n_480), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_521), .A2(n_470), .B1(n_443), .B2(n_479), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_514), .B(n_456), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_568), .B(n_480), .C(n_470), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_510), .B(n_456), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_557), .A2(n_470), .B(n_434), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_521), .A2(n_537), .B1(n_587), .B2(n_560), .C(n_511), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_533), .A2(n_434), .B1(n_224), .B2(n_266), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_533), .A2(n_434), .B1(n_224), .B2(n_305), .Y(n_615) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_562), .A2(n_9), .B(n_10), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_563), .B(n_11), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_566), .B(n_306), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_549), .B(n_12), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_538), .B(n_311), .C(n_292), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_559), .B(n_12), .Y(n_621) );
AND2x2_ASAP7_75t_SL g622 ( .A(n_544), .B(n_249), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_577), .B(n_566), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_551), .B(n_180), .C(n_190), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_551), .B(n_323), .C(n_309), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_577), .B(n_13), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_509), .A2(n_310), .B1(n_314), .B2(n_309), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_569), .B(n_323), .C(n_309), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_589), .B(n_14), .Y(n_629) );
NAND3xp33_ASAP7_75t_SL g630 ( .A(n_546), .B(n_14), .C(n_15), .Y(n_630) );
OAI21xp5_ASAP7_75t_SL g631 ( .A1(n_509), .A2(n_296), .B(n_300), .Y(n_631) );
OAI21xp33_ASAP7_75t_SL g632 ( .A1(n_528), .A2(n_296), .B(n_300), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_589), .B(n_15), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_507), .A2(n_310), .B1(n_314), .B2(n_309), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_524), .B(n_16), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_531), .B(n_323), .C(n_272), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_535), .B(n_16), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_564), .B(n_17), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_556), .B(n_18), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_528), .B(n_306), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_564), .B(n_19), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_525), .B(n_20), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_516), .A2(n_20), .B1(n_21), .B2(n_22), .C(n_23), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_564), .B(n_534), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_532), .B(n_21), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_564), .B(n_22), .Y(n_646) );
AOI21xp5_ASAP7_75t_SL g647 ( .A1(n_565), .A2(n_23), .B(n_24), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_541), .B(n_24), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_512), .A2(n_310), .B1(n_314), .B2(n_292), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_515), .B(n_25), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g651 ( .A1(n_565), .A2(n_303), .B(n_302), .Y(n_651) );
OAI21xp5_ASAP7_75t_SL g652 ( .A1(n_517), .A2(n_303), .B(n_302), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_518), .A2(n_520), .B1(n_522), .B2(n_553), .Y(n_653) );
AND2x2_ASAP7_75t_SL g654 ( .A(n_542), .B(n_296), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_553), .A2(n_292), .B1(n_315), .B2(n_306), .Y(n_655) );
OAI21xp5_ASAP7_75t_SL g656 ( .A1(n_567), .A2(n_303), .B(n_302), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_595), .B(n_26), .Y(n_657) );
NOR3xp33_ASAP7_75t_SL g658 ( .A(n_526), .B(n_28), .C(n_29), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_578), .B(n_28), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_548), .B(n_582), .C(n_575), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_598), .B(n_29), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_545), .A2(n_315), .B1(n_306), .B2(n_311), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_576), .B(n_581), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_596), .B(n_30), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_597), .B(n_31), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_574), .B(n_31), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_585), .B(n_251), .C(n_297), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_593), .B(n_33), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_576), .B(n_315), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_527), .B(n_34), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_529), .B(n_35), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_530), .B(n_36), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_552), .B(n_37), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_539), .B(n_37), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_523), .A2(n_224), .B1(n_297), .B2(n_311), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_543), .B(n_38), .Y(n_676) );
NAND3xp33_ASAP7_75t_L g677 ( .A(n_579), .B(n_297), .C(n_303), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_519), .B(n_38), .Y(n_678) );
INVxp67_ASAP7_75t_L g679 ( .A(n_588), .Y(n_679) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_561), .B(n_302), .C(n_300), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_536), .B(n_39), .Y(n_681) );
OAI221xp5_ASAP7_75t_SL g682 ( .A1(n_508), .A2(n_300), .B1(n_296), .B2(n_315), .C(n_293), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_571), .B(n_547), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_550), .A2(n_315), .B1(n_232), .B2(n_293), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_513), .A2(n_293), .B1(n_258), .B2(n_264), .Y(n_685) );
NAND4xp25_ASAP7_75t_L g686 ( .A(n_558), .B(n_41), .C(n_45), .D(n_49), .Y(n_686) );
OAI221xp5_ASAP7_75t_L g687 ( .A1(n_555), .A2(n_50), .B1(n_53), .B2(n_54), .C(n_55), .Y(n_687) );
OAI221xp5_ASAP7_75t_SL g688 ( .A1(n_570), .A2(n_56), .B1(n_59), .B2(n_62), .C(n_63), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_554), .B(n_65), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_572), .B(n_66), .C(n_69), .Y(n_690) );
OAI31xp33_ASAP7_75t_SL g691 ( .A1(n_594), .A2(n_71), .A3(n_72), .B(n_74), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_592), .A2(n_75), .B1(n_77), .B2(n_80), .Y(n_692) );
NOR2xp67_ASAP7_75t_L g693 ( .A(n_601), .B(n_81), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_540), .A2(n_82), .B1(n_83), .B2(n_84), .C(n_85), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_590), .A2(n_239), .B1(n_87), .B2(n_88), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_599), .B(n_86), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_605), .B(n_601), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_623), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_613), .B(n_573), .Y(n_699) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_630), .B(n_586), .C(n_583), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_609), .B(n_600), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_604), .B(n_591), .C(n_602), .Y(n_702) );
OA211x2_ASAP7_75t_L g703 ( .A1(n_612), .A2(n_90), .B(n_91), .C(n_92), .Y(n_703) );
AND2x4_ASAP7_75t_L g704 ( .A(n_644), .B(n_93), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_658), .B(n_94), .C(n_95), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_606), .B(n_98), .Y(n_706) );
BUFx2_ASAP7_75t_L g707 ( .A(n_609), .Y(n_707) );
NOR2xp33_ASAP7_75t_SL g708 ( .A(n_607), .B(n_622), .Y(n_708) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_654), .A2(n_683), .B1(n_644), .B2(n_632), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_608), .A2(n_631), .B1(n_615), .B2(n_683), .Y(n_710) );
AOI211xp5_ASAP7_75t_L g711 ( .A1(n_647), .A2(n_611), .B(n_691), .C(n_653), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_611), .B(n_610), .C(n_660), .Y(n_712) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_654), .A2(n_641), .B1(n_638), .B2(n_651), .Y(n_713) );
AO21x2_ASAP7_75t_L g714 ( .A1(n_617), .A2(n_663), .B(n_693), .Y(n_714) );
OA211x2_ASAP7_75t_L g715 ( .A1(n_663), .A2(n_608), .B(n_640), .C(n_615), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_679), .B(n_637), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_656), .A2(n_652), .B1(n_641), .B2(n_614), .Y(n_717) );
OR2x2_ASAP7_75t_L g718 ( .A(n_619), .B(n_626), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_639), .B(n_621), .Y(n_719) );
OAI211xp5_ASAP7_75t_SL g720 ( .A1(n_614), .A2(n_643), .B(n_650), .C(n_642), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_676), .B(n_640), .Y(n_721) );
OAI211xp5_ASAP7_75t_L g722 ( .A1(n_686), .A2(n_646), .B(n_657), .C(n_675), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_629), .B(n_633), .Y(n_723) );
AND2x4_ASAP7_75t_L g724 ( .A(n_676), .B(n_618), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_603), .B(n_627), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_603), .B(n_670), .Y(n_726) );
OR2x2_ASAP7_75t_L g727 ( .A(n_603), .B(n_635), .Y(n_727) );
INVx4_ASAP7_75t_L g728 ( .A(n_681), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_661), .B(n_664), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_665), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_645), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_674), .A2(n_648), .B1(n_678), .B2(n_673), .Y(n_732) );
OR2x2_ASAP7_75t_L g733 ( .A(n_624), .B(n_669), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_671), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_672), .B(n_659), .Y(n_735) );
AO21x2_ASAP7_75t_L g736 ( .A1(n_696), .A2(n_668), .B(n_666), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_628), .Y(n_737) );
NOR3xp33_ASAP7_75t_SL g738 ( .A(n_682), .B(n_688), .C(n_649), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_625), .B(n_680), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_694), .B(n_687), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_689), .B(n_634), .Y(n_741) );
OR2x2_ASAP7_75t_L g742 ( .A(n_685), .B(n_677), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_675), .A2(n_695), .B1(n_690), .B2(n_684), .Y(n_743) );
AO21x1_ASAP7_75t_SL g744 ( .A1(n_695), .A2(n_692), .B(n_655), .Y(n_744) );
NOR3xp33_ASAP7_75t_L g745 ( .A(n_620), .B(n_667), .C(n_636), .Y(n_745) );
NAND4xp75_ASAP7_75t_L g746 ( .A(n_662), .B(n_622), .C(n_616), .D(n_611), .Y(n_746) );
NAND2x1_ASAP7_75t_L g747 ( .A(n_647), .B(n_528), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_613), .B(n_445), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_604), .A2(n_613), .B1(n_683), .B2(n_653), .Y(n_749) );
NAND4xp75_ASAP7_75t_L g750 ( .A(n_622), .B(n_616), .C(n_611), .D(n_658), .Y(n_750) );
AO21x2_ASAP7_75t_L g751 ( .A1(n_611), .A2(n_617), .B(n_616), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g752 ( .A(n_604), .B(n_658), .C(n_616), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_623), .B(n_644), .Y(n_753) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_604), .B(n_658), .C(n_616), .Y(n_754) );
OAI21xp5_ASAP7_75t_L g755 ( .A1(n_647), .A2(n_663), .B(n_658), .Y(n_755) );
NAND4xp75_ASAP7_75t_L g756 ( .A(n_622), .B(n_616), .C(n_611), .D(n_658), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g757 ( .A(n_611), .B(n_510), .Y(n_757) );
NOR3xp33_ASAP7_75t_L g758 ( .A(n_616), .B(n_630), .C(n_465), .Y(n_758) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_707), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_708), .B(n_712), .Y(n_760) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_749), .B(n_711), .C(n_755), .Y(n_761) );
XNOR2xp5_ASAP7_75t_L g762 ( .A(n_715), .B(n_710), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_709), .A2(n_710), .B1(n_699), .B2(n_745), .Y(n_763) );
NAND4xp25_ASAP7_75t_L g764 ( .A(n_752), .B(n_754), .C(n_755), .D(n_748), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_698), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_727), .Y(n_766) );
XOR2x2_ASAP7_75t_L g767 ( .A(n_750), .B(n_756), .Y(n_767) );
XNOR2x2_ASAP7_75t_L g768 ( .A(n_746), .B(n_757), .Y(n_768) );
XOR2x2_ASAP7_75t_L g769 ( .A(n_717), .B(n_747), .Y(n_769) );
NAND4xp75_ASAP7_75t_SL g770 ( .A(n_740), .B(n_726), .C(n_744), .D(n_741), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_697), .Y(n_771) );
NOR3xp33_ASAP7_75t_L g772 ( .A(n_720), .B(n_745), .C(n_705), .Y(n_772) );
NAND3xp33_ASAP7_75t_L g773 ( .A(n_758), .B(n_709), .C(n_738), .Y(n_773) );
XNOR2xp5_ASAP7_75t_L g774 ( .A(n_713), .B(n_716), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_719), .B(n_728), .Y(n_775) );
XOR2x2_ASAP7_75t_L g776 ( .A(n_702), .B(n_732), .Y(n_776) );
XNOR2xp5_ASAP7_75t_L g777 ( .A(n_718), .B(n_723), .Y(n_777) );
NAND4xp75_ASAP7_75t_L g778 ( .A(n_703), .B(n_730), .C(n_731), .D(n_734), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_701), .B(n_753), .Y(n_779) );
XNOR2x2_ASAP7_75t_L g780 ( .A(n_743), .B(n_742), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_725), .B(n_721), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_725), .B(n_724), .Y(n_782) );
XNOR2xp5_ASAP7_75t_L g783 ( .A(n_735), .B(n_729), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_736), .B(n_751), .Y(n_784) );
XOR2xp5_ASAP7_75t_L g785 ( .A(n_706), .B(n_739), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_720), .B(n_722), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_733), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_737), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_751), .B(n_736), .Y(n_789) );
OR2x2_ASAP7_75t_L g790 ( .A(n_714), .B(n_704), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_759), .Y(n_791) );
INVxp33_ASAP7_75t_L g792 ( .A(n_785), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_782), .B(n_714), .Y(n_793) );
OA22x2_ASAP7_75t_L g794 ( .A1(n_762), .A2(n_704), .B1(n_722), .B2(n_743), .Y(n_794) );
INVx2_ASAP7_75t_SL g795 ( .A(n_765), .Y(n_795) );
XNOR2xp5_ASAP7_75t_L g796 ( .A(n_767), .B(n_700), .Y(n_796) );
INVxp67_ASAP7_75t_L g797 ( .A(n_761), .Y(n_797) );
INVxp67_ASAP7_75t_L g798 ( .A(n_787), .Y(n_798) );
XNOR2x1_ASAP7_75t_L g799 ( .A(n_780), .B(n_767), .Y(n_799) );
XOR2x2_ASAP7_75t_L g800 ( .A(n_773), .B(n_762), .Y(n_800) );
INVxp33_ASAP7_75t_L g801 ( .A(n_785), .Y(n_801) );
BUFx3_ASAP7_75t_L g802 ( .A(n_768), .Y(n_802) );
XNOR2xp5_ASAP7_75t_L g803 ( .A(n_769), .B(n_773), .Y(n_803) );
XOR2x2_ASAP7_75t_L g804 ( .A(n_769), .B(n_780), .Y(n_804) );
INVxp67_ASAP7_75t_L g805 ( .A(n_764), .Y(n_805) );
OR2x2_ASAP7_75t_L g806 ( .A(n_771), .B(n_766), .Y(n_806) );
INVx3_ASAP7_75t_L g807 ( .A(n_790), .Y(n_807) );
OA22x2_ASAP7_75t_L g808 ( .A1(n_803), .A2(n_760), .B1(n_774), .B2(n_783), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_806), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_799), .A2(n_763), .B1(n_786), .B2(n_776), .Y(n_810) );
OA22x2_ASAP7_75t_L g811 ( .A1(n_803), .A2(n_774), .B1(n_783), .B2(n_768), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_806), .Y(n_812) );
XNOR2xp5_ASAP7_75t_L g813 ( .A(n_804), .B(n_770), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_798), .Y(n_814) );
AOI22x1_ASAP7_75t_L g815 ( .A1(n_796), .A2(n_784), .B1(n_790), .B2(n_764), .Y(n_815) );
OAI22x1_ASAP7_75t_L g816 ( .A1(n_796), .A2(n_775), .B1(n_777), .B2(n_784), .Y(n_816) );
AOI22x1_ASAP7_75t_L g817 ( .A1(n_797), .A2(n_766), .B1(n_782), .B2(n_777), .Y(n_817) );
XNOR2x1_ASAP7_75t_L g818 ( .A(n_799), .B(n_776), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_795), .Y(n_819) );
AO22x2_ASAP7_75t_L g820 ( .A1(n_802), .A2(n_789), .B1(n_778), .B2(n_788), .Y(n_820) );
OA22x2_ASAP7_75t_L g821 ( .A1(n_805), .A2(n_766), .B1(n_781), .B2(n_771), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_795), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_814), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_809), .Y(n_824) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_819), .Y(n_825) );
INVxp67_ASAP7_75t_L g826 ( .A(n_822), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_812), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_811), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_811), .Y(n_829) );
BUFx2_ASAP7_75t_L g830 ( .A(n_820), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_828), .A2(n_794), .B1(n_804), .B2(n_808), .Y(n_831) );
NAND4xp25_ASAP7_75t_L g832 ( .A(n_829), .B(n_802), .C(n_810), .D(n_772), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_825), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_830), .A2(n_816), .B1(n_810), .B2(n_813), .C(n_820), .Y(n_834) );
OAI22x1_ASAP7_75t_L g835 ( .A1(n_830), .A2(n_815), .B1(n_817), .B2(n_800), .Y(n_835) );
OAI22x1_ASAP7_75t_L g836 ( .A1(n_831), .A2(n_823), .B1(n_800), .B2(n_818), .Y(n_836) );
A2O1A1Ixp33_ASAP7_75t_SL g837 ( .A1(n_833), .A2(n_823), .B(n_826), .C(n_827), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_832), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_838), .Y(n_839) );
INVxp67_ASAP7_75t_L g840 ( .A(n_836), .Y(n_840) );
INVxp67_ASAP7_75t_L g841 ( .A(n_839), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_840), .Y(n_842) );
AO22x2_ASAP7_75t_L g843 ( .A1(n_842), .A2(n_837), .B1(n_824), .B2(n_827), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_841), .Y(n_844) );
XNOR2xp5_ASAP7_75t_L g845 ( .A(n_843), .B(n_834), .Y(n_845) );
OAI22x1_ASAP7_75t_L g846 ( .A1(n_845), .A2(n_844), .B1(n_835), .B2(n_808), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_846), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_847), .A2(n_801), .B1(n_792), .B2(n_794), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_848), .Y(n_849) );
OAI22xp33_ASAP7_75t_L g850 ( .A1(n_849), .A2(n_794), .B1(n_824), .B2(n_821), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_850), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g852 ( .A1(n_851), .A2(n_820), .B1(n_807), .B2(n_791), .C(n_793), .Y(n_852) );
AOI211xp5_ASAP7_75t_L g853 ( .A1(n_852), .A2(n_791), .B(n_793), .C(n_779), .Y(n_853) );
endmodule