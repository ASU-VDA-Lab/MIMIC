module fake_jpeg_3903_n_109 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

AND2x2_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_24),
.Y(n_35)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_1),
.Y(n_24)
);

HAxp5_ASAP7_75t_SL g25 ( 
.A(n_12),
.B(n_2),
.CON(n_25),
.SN(n_25)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_20),
.B1(n_13),
.B2(n_15),
.Y(n_37)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx5_ASAP7_75t_SL g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2x1_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_20),
.B1(n_12),
.B2(n_14),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_21),
.B1(n_13),
.B2(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_R g39 ( 
.A(n_35),
.B(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_27),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_48),
.B1(n_38),
.B2(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_51),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_56),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_11),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_47),
.B1(n_45),
.B2(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_34),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_23),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_27),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_56),
.B(n_51),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_75),
.B1(n_78),
.B2(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_54),
.B(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_76),
.Y(n_81)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_34),
.A3(n_27),
.B1(n_11),
.B2(n_10),
.C1(n_49),
.C2(n_30),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_63),
.A3(n_62),
.B1(n_69),
.B2(n_66),
.C1(n_61),
.C2(n_22),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_10),
.C(n_15),
.Y(n_82)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_85),
.B1(n_84),
.B2(n_83),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_86),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_28),
.B1(n_17),
.B2(n_33),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_28),
.C(n_33),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_90),
.A2(n_92),
.B1(n_87),
.B2(n_91),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_70),
.B(n_86),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_17),
.B1(n_7),
.B2(n_8),
.Y(n_94)
);

XOR2x2_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_28),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_33),
.C(n_17),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_94),
.C(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_97),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_7),
.B1(n_8),
.B2(n_4),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_96),
.B(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_2),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_95),
.B(n_3),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_2),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_102),
.C(n_106),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_4),
.Y(n_109)
);


endmodule