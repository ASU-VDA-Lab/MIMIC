module fake_jpeg_17826_n_29 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

INVx6_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_12),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.C(n_2),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_21),
.C(n_16),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_11),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_22),
.C(n_16),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_20),
.B2(n_13),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_6),
.C(n_7),
.Y(n_29)
);


endmodule