module fake_ibex_1293_n_2158 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_357, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_366, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_78, n_20, n_69, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_2158);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_357;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_366;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_2158;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_766;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_1930;
wire n_2123;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1954;
wire n_1859;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_1971;
wire n_879;
wire n_1957;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_2112;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_737;
wire n_606;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_395;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_864;
wire n_608;
wire n_412;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_585;
wire n_1982;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_388;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_650;
wire n_409;
wire n_1575;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2095;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_961;
wire n_991;
wire n_634;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_403;
wire n_1353;
wire n_423;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_1830;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_1135;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_934;
wire n_520;
wire n_775;
wire n_950;
wire n_512;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_2078;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_2093;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_753;
wire n_2126;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_383;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_417;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2079;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1385;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2092;
wire n_566;
wire n_581;
wire n_416;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_405;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_414;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_519;
wire n_1843;
wire n_408;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_148),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_131),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_161),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_321),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_121),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_270),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_211),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_367),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_95),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_96),
.Y(n_393)
);

BUFx2_ASAP7_75t_SL g394 ( 
.A(n_223),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_68),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_157),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_11),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_361),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_81),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_196),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_190),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_18),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_86),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_228),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_10),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_L g408 ( 
.A(n_242),
.B(n_296),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_245),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_162),
.B(n_339),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_124),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_212),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_85),
.Y(n_413)
);

BUFx5_ASAP7_75t_L g414 ( 
.A(n_205),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_217),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_87),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_232),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_74),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_264),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_241),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_314),
.Y(n_421)
);

BUFx10_ASAP7_75t_L g422 ( 
.A(n_85),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_61),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_250),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_153),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_309),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_32),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_188),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_257),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_350),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_240),
.B(n_202),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_145),
.Y(n_432)
);

BUFx2_ASAP7_75t_SL g433 ( 
.A(n_362),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_348),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_200),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_283),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_281),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_382),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_80),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_138),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_58),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g442 ( 
.A(n_65),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_187),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_158),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_252),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_44),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_319),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_47),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_124),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_304),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_246),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_139),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_163),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_363),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_59),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_117),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_369),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_364),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_357),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_347),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_322),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_134),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_237),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_103),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_92),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_259),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_130),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_127),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_333),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_25),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_316),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_268),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_197),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_327),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_301),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_274),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_80),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_298),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_276),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_289),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_312),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_288),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_195),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_377),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_79),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_21),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_336),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_230),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_194),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_313),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_265),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_58),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_260),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_30),
.Y(n_495)
);

BUFx8_ASAP7_75t_SL g496 ( 
.A(n_249),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_111),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_98),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_105),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_96),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_147),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_4),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_318),
.Y(n_503)
);

XOR2x2_ASAP7_75t_L g504 ( 
.A(n_109),
.B(n_285),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_208),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_238),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_284),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_253),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_227),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_305),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_179),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_100),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_152),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_66),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_104),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_132),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_14),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_107),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_297),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_287),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_46),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_109),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_375),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_1),
.B(n_278),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_291),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_37),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_75),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_103),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_365),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_300),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_299),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_323),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_20),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_275),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_38),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_277),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_349),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_306),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_6),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_123),
.Y(n_540)
);

CKINVDCx14_ASAP7_75t_R g541 ( 
.A(n_156),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_192),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_43),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_38),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_104),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_273),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_243),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_125),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_102),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_78),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_343),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_52),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_332),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_218),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_112),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_263),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_201),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_235),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_311),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_126),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_79),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_226),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_106),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_140),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_216),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_247),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_99),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_293),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_119),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_52),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_29),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_220),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_368),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_129),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_17),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_91),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_100),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_167),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_63),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_48),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_310),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_222),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_282),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_50),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_114),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_106),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_14),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_213),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_143),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_154),
.Y(n_590)
);

CKINVDCx16_ASAP7_75t_R g591 ( 
.A(n_76),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_126),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_359),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_83),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_272),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_153),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_206),
.Y(n_597)
);

BUFx8_ASAP7_75t_SL g598 ( 
.A(n_302),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_324),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_33),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_162),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_150),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_2),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_340),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_105),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_75),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_320),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_92),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_358),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_23),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g611 ( 
.A(n_308),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_90),
.Y(n_612)
);

BUFx2_ASAP7_75t_SL g613 ( 
.A(n_307),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_219),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_191),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_48),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_239),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_189),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_178),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_225),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_130),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_183),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_145),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_334),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_49),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_244),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_251),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_20),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_381),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_182),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_78),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_355),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_269),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_76),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_41),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_46),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_10),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_255),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_62),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_203),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_271),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_163),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_150),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_7),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_166),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_42),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_121),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_236),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_73),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_116),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_102),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_229),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_84),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_207),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_345),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_28),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_11),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_331),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_87),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_267),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_101),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_15),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_214),
.B(n_317),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_118),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_110),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_142),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_373),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_1),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_8),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_209),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_72),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_49),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_342),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_152),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_290),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_50),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_107),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_147),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_376),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_29),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_338),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_128),
.Y(n_682)
);

BUFx8_ASAP7_75t_SL g683 ( 
.A(n_405),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_525),
.B(n_463),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_403),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_389),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_525),
.B(n_0),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_403),
.Y(n_688)
);

BUFx8_ASAP7_75t_L g689 ( 
.A(n_480),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_402),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_516),
.B(n_0),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_489),
.B(n_2),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_459),
.B(n_3),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_469),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_396),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_396),
.B(n_3),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_442),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_535),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_535),
.Y(n_699)
);

BUFx12f_ASAP7_75t_L g700 ( 
.A(n_422),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_403),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_484),
.Y(n_702)
);

BUFx8_ASAP7_75t_L g703 ( 
.A(n_590),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_389),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_449),
.Y(n_705)
);

BUFx8_ASAP7_75t_SL g706 ( 
.A(n_405),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_403),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_414),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_421),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_496),
.Y(n_710)
);

INVx5_ASAP7_75t_L g711 ( 
.A(n_484),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_421),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_384),
.B(n_5),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_384),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_418),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_449),
.B(n_8),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_499),
.B(n_9),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_430),
.B(n_9),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_419),
.Y(n_719)
);

OA21x2_ASAP7_75t_L g720 ( 
.A1(n_398),
.A2(n_172),
.B(n_171),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_499),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_418),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_491),
.B(n_12),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_417),
.B(n_173),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_421),
.Y(n_725)
);

INVx5_ASAP7_75t_L g726 ( 
.A(n_484),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_486),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_422),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_541),
.Y(n_729)
);

OAI21x1_ASAP7_75t_L g730 ( 
.A1(n_398),
.A2(n_175),
.B(n_174),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_537),
.B(n_12),
.Y(n_731)
);

BUFx8_ASAP7_75t_L g732 ( 
.A(n_612),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_601),
.B(n_13),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_421),
.Y(n_734)
);

OA21x2_ASAP7_75t_L g735 ( 
.A1(n_420),
.A2(n_177),
.B(n_176),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_601),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_541),
.A2(n_16),
.B1(n_13),
.B2(n_15),
.Y(n_737)
);

BUFx8_ASAP7_75t_L g738 ( 
.A(n_616),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_482),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_496),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_385),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_414),
.Y(n_742)
);

CKINVDCx6p67_ASAP7_75t_R g743 ( 
.A(n_568),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_414),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_473),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_393),
.B(n_19),
.Y(n_746)
);

BUFx12f_ASAP7_75t_L g747 ( 
.A(n_637),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_407),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_413),
.B(n_19),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_637),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_414),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_383),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_517),
.B(n_22),
.Y(n_753)
);

INVx5_ASAP7_75t_L g754 ( 
.A(n_568),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_432),
.B(n_22),
.Y(n_755)
);

INVx5_ASAP7_75t_L g756 ( 
.A(n_568),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_549),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_419),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_440),
.Y(n_759)
);

OA21x2_ASAP7_75t_L g760 ( 
.A1(n_420),
.A2(n_181),
.B(n_180),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_441),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_482),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_482),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_637),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_564),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_454),
.Y(n_766)
);

BUFx8_ASAP7_75t_SL g767 ( 
.A(n_471),
.Y(n_767)
);

OA21x2_ASAP7_75t_L g768 ( 
.A1(n_445),
.A2(n_185),
.B(n_184),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_556),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_482),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_388),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_454),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_454),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_558),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_611),
.A2(n_27),
.B1(n_24),
.B2(n_26),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_558),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_468),
.B(n_24),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_478),
.B(n_26),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_666),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_445),
.A2(n_483),
.B(n_455),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_493),
.B(n_27),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_501),
.B(n_28),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_502),
.B(n_513),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_522),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_454),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_558),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_591),
.B(n_30),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_666),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_533),
.B(n_31),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_558),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_495),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_556),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_392),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_540),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_673),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_R g796 ( 
.A(n_710),
.B(n_412),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_695),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_695),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_687),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_683),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_780),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_683),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_706),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_706),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_687),
.Y(n_805)
);

AND3x2_ASAP7_75t_L g806 ( 
.A(n_757),
.B(n_729),
.C(n_705),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_765),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_765),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_700),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_767),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_767),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_740),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_R g813 ( 
.A(n_728),
.B(n_412),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_708),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_713),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_740),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_747),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_743),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_689),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_689),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_703),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_703),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_713),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_684),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_R g825 ( 
.A(n_728),
.B(n_461),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_732),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_732),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_729),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_742),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_738),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_R g831 ( 
.A(n_750),
.B(n_461),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_697),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_721),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_733),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_752),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_752),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_771),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_733),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_684),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_771),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_746),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_793),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_793),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_749),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_795),
.B(n_387),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_744),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_795),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_702),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_L g849 ( 
.A(n_702),
.B(n_406),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_702),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_702),
.Y(n_851)
);

XNOR2xp5_ASAP7_75t_L g852 ( 
.A(n_753),
.B(n_504),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_746),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_711),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_711),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_787),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_696),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_711),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_711),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_726),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_751),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_716),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_726),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_789),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_694),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_698),
.Y(n_866)
);

CKINVDCx6p67_ASAP7_75t_R g867 ( 
.A(n_726),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_685),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_717),
.Y(n_869)
);

CKINVDCx16_ASAP7_75t_R g870 ( 
.A(n_724),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_754),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_754),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_750),
.B(n_666),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_699),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_730),
.A2(n_483),
.B(n_455),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_754),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_756),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_756),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_756),
.B(n_682),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_R g880 ( 
.A(n_764),
.B(n_492),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_779),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_685),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_720),
.A2(n_531),
.B(n_508),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_745),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_690),
.B(n_425),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_775),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_686),
.B(n_395),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_737),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_691),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_788),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_691),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_783),
.Y(n_892)
);

CKINVDCx16_ASAP7_75t_R g893 ( 
.A(n_724),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_783),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_692),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_741),
.B(n_508),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_704),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_718),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_737),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_704),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_718),
.Y(n_901)
);

CKINVDCx16_ASAP7_75t_R g902 ( 
.A(n_692),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_719),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_758),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_758),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_769),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_792),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_792),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_685),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_693),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_693),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_723),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_R g913 ( 
.A(n_748),
.B(n_492),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_759),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_723),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_761),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_784),
.B(n_543),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_714),
.Y(n_918)
);

INVxp33_ASAP7_75t_SL g919 ( 
.A(n_731),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_794),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_755),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_777),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_715),
.B(n_531),
.Y(n_923)
);

BUFx10_ASAP7_75t_L g924 ( 
.A(n_722),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_777),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_727),
.Y(n_926)
);

BUFx10_ASAP7_75t_L g927 ( 
.A(n_736),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_778),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_735),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_778),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_781),
.Y(n_931)
);

BUFx10_ASAP7_75t_L g932 ( 
.A(n_685),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_782),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_782),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_766),
.B(n_415),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_791),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_772),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_773),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_785),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_688),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_688),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_688),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_720),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_720),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_688),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_760),
.Y(n_946)
);

AND2x6_ASAP7_75t_L g947 ( 
.A(n_701),
.B(n_582),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_760),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_760),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_735),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_701),
.Y(n_951)
);

NOR2xp67_ASAP7_75t_L g952 ( 
.A(n_701),
.B(n_426),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_768),
.B(n_673),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_707),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_707),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_709),
.B(n_435),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_709),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_L g958 ( 
.A(n_709),
.B(n_437),
.Y(n_958)
);

AND2x6_ASAP7_75t_L g959 ( 
.A(n_712),
.B(n_582),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_712),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_712),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_712),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_725),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_725),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_725),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_734),
.Y(n_966)
);

BUFx10_ASAP7_75t_L g967 ( 
.A(n_734),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_734),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_734),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_739),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_739),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_739),
.Y(n_972)
);

BUFx10_ASAP7_75t_L g973 ( 
.A(n_739),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_762),
.B(n_763),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_762),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_919),
.B(n_898),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_901),
.B(n_386),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_933),
.Y(n_978)
);

BUFx12f_ASAP7_75t_SL g979 ( 
.A(n_809),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_912),
.B(n_673),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_SL g981 ( 
.A(n_913),
.B(n_509),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_889),
.B(n_446),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_891),
.B(n_519),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_824),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_924),
.Y(n_985)
);

NAND2xp33_ASAP7_75t_L g986 ( 
.A(n_953),
.B(n_390),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_915),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_924),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_925),
.B(n_464),
.Y(n_989)
);

AO221x1_ASAP7_75t_L g990 ( 
.A1(n_913),
.A2(n_825),
.B1(n_880),
.B2(n_831),
.C(n_813),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_SL g991 ( 
.A1(n_805),
.A2(n_552),
.B(n_548),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_817),
.B(n_32),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_918),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_928),
.B(n_474),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_927),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_930),
.B(n_476),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_841),
.A2(n_560),
.B1(n_567),
.B2(n_555),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_914),
.B(n_391),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_931),
.B(n_477),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_920),
.B(n_504),
.Y(n_1000)
);

AO221x1_ASAP7_75t_L g1001 ( 
.A1(n_813),
.A2(n_880),
.B1(n_831),
.B2(n_825),
.C(n_870),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_801),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_916),
.B(n_399),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_927),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_839),
.Y(n_1005)
);

NAND3xp33_ASAP7_75t_L g1006 ( 
.A(n_946),
.B(n_485),
.C(n_479),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_L g1007 ( 
.A(n_943),
.B(n_503),
.C(n_490),
.Y(n_1007)
);

NAND2xp33_ASAP7_75t_L g1008 ( 
.A(n_934),
.B(n_401),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_837),
.B(n_828),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_801),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_929),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_835),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_926),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_917),
.B(n_799),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_865),
.Y(n_1015)
);

OA21x2_ASAP7_75t_L g1016 ( 
.A1(n_883),
.A2(n_875),
.B(n_949),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_897),
.B(n_900),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_903),
.B(n_409),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_904),
.B(n_424),
.Y(n_1019)
);

CKINVDCx11_ASAP7_75t_R g1020 ( 
.A(n_807),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_853),
.B(n_428),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_866),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_905),
.B(n_429),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_906),
.B(n_434),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_874),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_L g1026 ( 
.A(n_902),
.B(n_457),
.C(n_444),
.Y(n_1026)
);

AO221x1_ASAP7_75t_L g1027 ( 
.A1(n_893),
.A2(n_598),
.B1(n_410),
.B2(n_509),
.C(n_530),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_938),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_929),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_853),
.B(n_436),
.Y(n_1030)
);

AND3x1_ASAP7_75t_L g1031 ( 
.A(n_873),
.B(n_570),
.C(n_569),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_836),
.B(n_397),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_847),
.B(n_895),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_845),
.B(n_438),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_815),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_823),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_939),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_887),
.B(n_443),
.Y(n_1038)
);

AND2x4_ASAP7_75t_SL g1039 ( 
.A(n_867),
.B(n_510),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_834),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_907),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_838),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_908),
.B(n_448),
.Y(n_1043)
);

BUFx8_ASAP7_75t_L g1044 ( 
.A(n_885),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_848),
.Y(n_1045)
);

NOR3xp33_ASAP7_75t_L g1046 ( 
.A(n_840),
.B(n_584),
.C(n_578),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_892),
.B(n_451),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_894),
.B(n_452),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_864),
.A2(n_576),
.B1(n_580),
.B2(n_575),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_935),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_947),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_923),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_842),
.B(n_642),
.C(n_587),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_923),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_843),
.B(n_672),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_832),
.B(n_400),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_881),
.B(n_458),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_SL g1058 ( 
.A(n_921),
.B(n_530),
.C(n_510),
.Y(n_1058)
);

INVxp67_ASAP7_75t_SL g1059 ( 
.A(n_961),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_872),
.B(n_532),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_896),
.B(n_538),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_814),
.B(n_542),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_814),
.B(n_546),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_829),
.B(n_581),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_850),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_910),
.B(n_460),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_L g1067 ( 
.A(n_950),
.B(n_588),
.C(n_583),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_849),
.B(n_594),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_911),
.B(n_462),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_833),
.B(n_467),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_796),
.B(n_394),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_879),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_L g1073 ( 
.A(n_812),
.B(n_411),
.C(n_404),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_851),
.B(n_854),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_855),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_922),
.A2(n_599),
.B1(n_640),
.B2(n_532),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_816),
.B(n_416),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_858),
.B(n_470),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_947),
.Y(n_1079)
);

INVxp33_ASAP7_75t_L g1080 ( 
.A(n_852),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_859),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_806),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_860),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_947),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_947),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_890),
.B(n_472),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_863),
.B(n_475),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_821),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_871),
.B(n_481),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_876),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_877),
.B(n_488),
.Y(n_1091)
);

NOR2xp67_ASAP7_75t_L g1092 ( 
.A(n_818),
.B(n_34),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_878),
.B(n_494),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_969),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_846),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_857),
.B(n_862),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_932),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_869),
.B(n_505),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_861),
.B(n_506),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_947),
.Y(n_1100)
);

AND2x6_ASAP7_75t_L g1101 ( 
.A(n_944),
.B(n_652),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_844),
.B(n_507),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_856),
.B(n_423),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_944),
.B(n_511),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_819),
.B(n_820),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_L g1106 ( 
.A(n_822),
.B(n_439),
.C(n_427),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_975),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_SL g1108 ( 
.A(n_948),
.B(n_640),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_952),
.Y(n_1109)
);

INVxp33_ASAP7_75t_L g1110 ( 
.A(n_808),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_936),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_884),
.B(n_520),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_956),
.B(n_523),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_958),
.B(n_529),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_937),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_L g1116 ( 
.A(n_940),
.B(n_604),
.C(n_595),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_886),
.B(n_826),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_827),
.B(n_536),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_932),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_967),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_967),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_959),
.B(n_547),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_959),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_L g1124 ( 
.A(n_830),
.B(n_450),
.C(n_447),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_973),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_797),
.B(n_551),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_888),
.B(n_453),
.Y(n_1127)
);

INVx8_ASAP7_75t_L g1128 ( 
.A(n_959),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_899),
.B(n_456),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_SL g1130 ( 
.A(n_959),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_965),
.A2(n_605),
.B(n_631),
.C(n_600),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_941),
.Y(n_1132)
);

NOR2xp67_ASAP7_75t_L g1133 ( 
.A(n_800),
.B(n_34),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_942),
.B(n_553),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_802),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_945),
.Y(n_1136)
);

INVxp33_ASAP7_75t_SL g1137 ( 
.A(n_803),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_951),
.B(n_554),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_954),
.B(n_557),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_973),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_SL g1141 ( 
.A(n_957),
.B(n_681),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_960),
.B(n_562),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_963),
.B(n_565),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_798),
.B(n_566),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_966),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_968),
.B(n_572),
.Y(n_1146)
);

INVxp33_ASAP7_75t_L g1147 ( 
.A(n_804),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_971),
.B(n_573),
.Y(n_1148)
);

INVxp33_ASAP7_75t_L g1149 ( 
.A(n_810),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_811),
.B(n_465),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_974),
.B(n_597),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_962),
.B(n_607),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_964),
.B(n_609),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_955),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_970),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_972),
.B(n_619),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_955),
.B(n_614),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_955),
.B(n_615),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_955),
.B(n_617),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_868),
.B(n_620),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_882),
.B(n_624),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_909),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_919),
.B(n_626),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_933),
.Y(n_1164)
);

INVx8_ASAP7_75t_L g1165 ( 
.A(n_872),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_898),
.B(n_622),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_915),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_933),
.B(n_466),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_824),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_801),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_933),
.Y(n_1171)
);

NAND2xp33_ASAP7_75t_L g1172 ( 
.A(n_953),
.B(n_632),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_889),
.B(n_681),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_801),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_824),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_898),
.B(n_627),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_889),
.A2(n_643),
.B1(n_644),
.B2(n_635),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_898),
.B(n_629),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_898),
.B(n_633),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_919),
.B(n_638),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_L g1181 ( 
.A(n_817),
.B(n_35),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_L g1182 ( 
.A(n_902),
.B(n_497),
.C(n_487),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_824),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_933),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_801),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_L g1186 ( 
.A(n_953),
.B(n_641),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_898),
.B(n_679),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_919),
.B(n_648),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_824),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_913),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_824),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_824),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_961),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_919),
.B(n_654),
.Y(n_1194)
);

INVxp67_ASAP7_75t_L g1195 ( 
.A(n_915),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_919),
.B(n_658),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1095),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1002),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1002),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1014),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1013),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_976),
.B(n_498),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_985),
.B(n_647),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_988),
.B(n_995),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1012),
.B(n_1076),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1167),
.B(n_471),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1094),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1195),
.B(n_606),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_978),
.A2(n_667),
.B1(n_512),
.B2(n_518),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1002),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1004),
.B(n_670),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1164),
.B(n_514),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1171),
.B(n_606),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1016),
.A2(n_431),
.B(n_408),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1009),
.A2(n_651),
.B1(n_659),
.B2(n_649),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1184),
.B(n_521),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_SL g1217 ( 
.A(n_1190),
.B(n_527),
.C(n_526),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1010),
.B(n_675),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_987),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1033),
.B(n_528),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1015),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1041),
.B(n_668),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_1044),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_983),
.B(n_539),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_991),
.A2(n_674),
.B(n_676),
.C(n_671),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1128),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_SL g1227 ( 
.A(n_1026),
.B(n_545),
.C(n_544),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1193),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_1128),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1022),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1041),
.B(n_677),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1031),
.A2(n_561),
.B1(n_563),
.B2(n_550),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_R g1233 ( 
.A(n_979),
.B(n_571),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_982),
.B(n_574),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_982),
.B(n_577),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1025),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1039),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1166),
.B(n_579),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_1128),
.Y(n_1239)
);

NOR3xp33_ASAP7_75t_L g1240 ( 
.A(n_1058),
.B(n_586),
.C(n_585),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1166),
.B(n_589),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1176),
.B(n_1178),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1031),
.B(n_1075),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1005),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1035),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1176),
.B(n_592),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1081),
.B(n_678),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1178),
.B(n_596),
.Y(n_1248)
);

AND2x4_ASAP7_75t_SL g1249 ( 
.A(n_1071),
.B(n_680),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1044),
.Y(n_1250)
);

NOR3xp33_ASAP7_75t_SL g1251 ( 
.A(n_1117),
.B(n_608),
.C(n_602),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1097),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1100),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1170),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1036),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1168),
.B(n_610),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1170),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1108),
.A2(n_623),
.B1(n_625),
.B2(n_621),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1051),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1108),
.A2(n_634),
.B1(n_636),
.B2(n_628),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1083),
.B(n_663),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_993),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1107),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_SL g1264 ( 
.A(n_1046),
.B(n_645),
.C(n_639),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1174),
.B(n_646),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1174),
.B(n_650),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1173),
.A2(n_656),
.B1(n_657),
.B2(n_653),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1000),
.B(n_661),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1165),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1040),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1042),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_984),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1169),
.Y(n_1273)
);

OR2x6_ASAP7_75t_L g1274 ( 
.A(n_1165),
.B(n_1071),
.Y(n_1274)
);

AO22x1_ASAP7_75t_L g1275 ( 
.A1(n_1060),
.A2(n_598),
.B1(n_664),
.B2(n_662),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1179),
.B(n_665),
.Y(n_1276)
);

INVx5_ASAP7_75t_L g1277 ( 
.A(n_1051),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1127),
.B(n_495),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_R g1279 ( 
.A(n_1020),
.B(n_35),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1180),
.A2(n_524),
.B1(n_613),
.B2(n_433),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1179),
.A2(n_515),
.B1(n_603),
.B2(n_500),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1090),
.B(n_500),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1185),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1045),
.B(n_603),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1165),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1056),
.B(n_1163),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1045),
.B(n_669),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1055),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1131),
.A2(n_559),
.B(n_593),
.C(n_534),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1079),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1175),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1079),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1137),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1188),
.A2(n_618),
.B1(n_630),
.B2(n_593),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1183),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1185),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1187),
.B(n_630),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1079),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1111),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_989),
.B(n_655),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1129),
.B(n_36),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_994),
.B(n_660),
.Y(n_1302)
);

NOR2x2_ASAP7_75t_L g1303 ( 
.A(n_1027),
.B(n_36),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1084),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1032),
.B(n_1077),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1059),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_994),
.B(n_39),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1141),
.Y(n_1308)
);

NAND3xp33_ASAP7_75t_SL g1309 ( 
.A(n_1053),
.B(n_39),
.C(n_40),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_996),
.B(n_40),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_996),
.A2(n_999),
.B1(n_1054),
.B2(n_1052),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1141),
.A2(n_770),
.B1(n_774),
.B2(n_763),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1080),
.A2(n_47),
.B1(n_44),
.B2(n_45),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1068),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1135),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_977),
.B(n_45),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1105),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1068),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1011),
.B(n_770),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1189),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1191),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1192),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1028),
.B(n_51),
.Y(n_1323)
);

BUFx12f_ASAP7_75t_L g1324 ( 
.A(n_1082),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1103),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1115),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1062),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1062),
.Y(n_1328)
);

AND2x6_ASAP7_75t_L g1329 ( 
.A(n_1029),
.B(n_770),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_R g1330 ( 
.A(n_981),
.B(n_51),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1119),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1096),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_980),
.B(n_53),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1088),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1120),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1029),
.B(n_1072),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1084),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1182),
.A2(n_776),
.B1(n_786),
.B2(n_774),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1102),
.Y(n_1339)
);

NOR2x1p5_ASAP7_75t_L g1340 ( 
.A(n_1150),
.B(n_54),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1098),
.Y(n_1341)
);

NAND2x1p5_ASAP7_75t_L g1342 ( 
.A(n_1065),
.B(n_54),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1037),
.B(n_55),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1110),
.A2(n_59),
.B1(n_56),
.B2(n_57),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1085),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1085),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1063),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1063),
.Y(n_1348)
);

AND2x6_ASAP7_75t_L g1349 ( 
.A(n_1085),
.B(n_786),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1064),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1112),
.A2(n_63),
.B1(n_60),
.B2(n_61),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1038),
.B(n_786),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1001),
.A2(n_790),
.B1(n_66),
.B2(n_64),
.Y(n_1353)
);

AND2x6_ASAP7_75t_L g1354 ( 
.A(n_1123),
.B(n_1132),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1064),
.Y(n_1355)
);

AND2x6_ASAP7_75t_L g1356 ( 
.A(n_1136),
.B(n_790),
.Y(n_1356)
);

AND2x4_ASAP7_75t_SL g1357 ( 
.A(n_1073),
.B(n_790),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1126),
.B(n_65),
.Y(n_1358)
);

NAND2x1p5_ASAP7_75t_L g1359 ( 
.A(n_1017),
.B(n_67),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1194),
.B(n_68),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1049),
.B(n_69),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1144),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1152),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1121),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_L g1365 ( 
.A(n_986),
.B(n_70),
.C(n_71),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1118),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1101),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1008),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_998),
.B(n_1003),
.Y(n_1369)
);

AO21x1_ASAP7_75t_L g1370 ( 
.A1(n_1104),
.A2(n_77),
.B(n_82),
.Y(n_1370)
);

INVx5_ASAP7_75t_L g1371 ( 
.A(n_1101),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1156),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1047),
.B(n_83),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1048),
.B(n_84),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1061),
.B(n_86),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1125),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1086),
.B(n_88),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1016),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1140),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1050),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_990),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1021),
.Y(n_1382)
);

AND2x6_ASAP7_75t_SL g1383 ( 
.A(n_1147),
.B(n_89),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1154),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1030),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1109),
.Y(n_1386)
);

AO22x1_ASAP7_75t_L g1387 ( 
.A1(n_1149),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1145),
.Y(n_1388)
);

NOR3xp33_ASAP7_75t_SL g1389 ( 
.A(n_1070),
.B(n_1069),
.C(n_1066),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1074),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1196),
.B(n_94),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1057),
.B(n_97),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1099),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1006),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1172),
.A2(n_110),
.B1(n_101),
.B2(n_108),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1186),
.A2(n_112),
.B1(n_108),
.B2(n_111),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1106),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1034),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1157),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1124),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1089),
.B(n_119),
.Y(n_1401)
);

NOR2xp67_ASAP7_75t_L g1402 ( 
.A(n_1092),
.B(n_120),
.Y(n_1402)
);

CKINVDCx11_ASAP7_75t_R g1403 ( 
.A(n_1133),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_992),
.B(n_120),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1158),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1181),
.B(n_1116),
.Y(n_1406)
);

AOI21xp33_ASAP7_75t_L g1407 ( 
.A1(n_1091),
.A2(n_122),
.B(n_123),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1242),
.A2(n_1007),
.B1(n_1067),
.B2(n_1116),
.Y(n_1408)
);

INVx4_ASAP7_75t_L g1409 ( 
.A(n_1274),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1288),
.B(n_1134),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1378),
.A2(n_1067),
.B(n_1151),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1311),
.B(n_1018),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1268),
.B(n_1093),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1221),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1206),
.B(n_1019),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1233),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1305),
.B(n_1023),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1200),
.B(n_1024),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1327),
.A2(n_1139),
.B1(n_1142),
.B2(n_1138),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1326),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1328),
.B(n_1043),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1347),
.B(n_1101),
.Y(n_1422)
);

NOR2x1_ASAP7_75t_L g1423 ( 
.A(n_1293),
.B(n_1148),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1348),
.A2(n_1146),
.B1(n_1143),
.B2(n_1087),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1350),
.B(n_1355),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1201),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1208),
.B(n_1078),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1207),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1219),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_R g1430 ( 
.A(n_1334),
.B(n_1223),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1390),
.B(n_1113),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1244),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1258),
.B(n_1122),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1279),
.Y(n_1434)
);

OAI21xp33_ASAP7_75t_L g1435 ( 
.A1(n_1300),
.A2(n_1159),
.B(n_1153),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1363),
.A2(n_1114),
.B(n_1161),
.C(n_1160),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1324),
.Y(n_1437)
);

NAND2x1p5_ASAP7_75t_L g1438 ( 
.A(n_1237),
.B(n_1130),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_SL g1439 ( 
.A(n_1330),
.B(n_1162),
.C(n_1155),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1250),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1245),
.B(n_122),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1255),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1270),
.B(n_125),
.Y(n_1443)
);

BUFx12f_ASAP7_75t_L g1444 ( 
.A(n_1274),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1209),
.B(n_127),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1285),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1299),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1275),
.Y(n_1448)
);

BUFx2_ASAP7_75t_SL g1449 ( 
.A(n_1269),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1372),
.A2(n_193),
.B(n_186),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1306),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1271),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1315),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1243),
.B(n_128),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1230),
.Y(n_1455)
);

AOI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1215),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.C(n_133),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1213),
.B(n_133),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1228),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1336),
.A2(n_1385),
.B(n_1382),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1339),
.B(n_134),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1393),
.A2(n_199),
.B(n_198),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1205),
.B(n_135),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1325),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1302),
.A2(n_1352),
.B(n_1297),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_R g1465 ( 
.A(n_1308),
.B(n_136),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1243),
.B(n_137),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1323),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_1467)
);

NOR2xp67_ASAP7_75t_L g1468 ( 
.A(n_1217),
.B(n_141),
.Y(n_1468)
);

AO32x2_ASAP7_75t_L g1469 ( 
.A1(n_1281),
.A2(n_141),
.A3(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1323),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1234),
.B(n_144),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_SL g1472 ( 
.A(n_1226),
.B(n_204),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1235),
.B(n_146),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1260),
.B(n_146),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1370),
.A2(n_148),
.A3(n_149),
.B(n_151),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1238),
.B(n_149),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1241),
.B(n_151),
.Y(n_1477)
);

BUFx12f_ASAP7_75t_L g1478 ( 
.A(n_1383),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1251),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1197),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1332),
.B(n_154),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1249),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1246),
.B(n_155),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1286),
.B(n_155),
.Y(n_1484)
);

CKINVDCx8_ASAP7_75t_R g1485 ( 
.A(n_1373),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1301),
.B(n_156),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1277),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1236),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_SL g1489 ( 
.A1(n_1220),
.A2(n_266),
.B(n_379),
.C(n_378),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1248),
.B(n_157),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1369),
.B(n_158),
.Y(n_1491)
);

NAND2x1p5_ASAP7_75t_L g1492 ( 
.A(n_1226),
.B(n_1229),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_R g1493 ( 
.A(n_1362),
.B(n_159),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1276),
.B(n_159),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1341),
.B(n_160),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1398),
.B(n_160),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1256),
.B(n_161),
.Y(n_1497)
);

BUFx4f_ASAP7_75t_L g1498 ( 
.A(n_1342),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1225),
.B(n_164),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1343),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1317),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1343),
.B(n_165),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1262),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1282),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1313),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_SL g1506 ( 
.A(n_1366),
.B(n_168),
.C(n_169),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1267),
.B(n_170),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1229),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1282),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1277),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1202),
.B(n_170),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1384),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1203),
.B(n_210),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1289),
.A2(n_1307),
.B(n_1310),
.C(n_1375),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1203),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1262),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1369),
.B(n_215),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_SL g1518 ( 
.A(n_1239),
.B(n_1371),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1222),
.B(n_221),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1278),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1222),
.B(n_224),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_SL g1522 ( 
.A(n_1239),
.B(n_231),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1247),
.B(n_233),
.Y(n_1523)
);

OR2x6_ASAP7_75t_SL g1524 ( 
.A(n_1358),
.B(n_234),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1373),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1247),
.B(n_248),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1253),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1263),
.B(n_254),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1272),
.Y(n_1529)
);

BUFx10_ASAP7_75t_L g1530 ( 
.A(n_1374),
.Y(n_1530)
);

OR2x6_ASAP7_75t_L g1531 ( 
.A(n_1314),
.B(n_256),
.Y(n_1531)
);

O2A1O1Ixp33_ASAP7_75t_SL g1532 ( 
.A1(n_1316),
.A2(n_258),
.B(n_261),
.C(n_262),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1273),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1318),
.B(n_380),
.Y(n_1534)
);

INVx4_ASAP7_75t_L g1535 ( 
.A(n_1277),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1291),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1374),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1295),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1198),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1214),
.A2(n_279),
.B(n_280),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1232),
.B(n_286),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1320),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1321),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1231),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1340),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1392),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1389),
.B(n_372),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1322),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1212),
.B(n_1216),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1392),
.B(n_303),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1204),
.B(n_371),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1401),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1377),
.B(n_1401),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1284),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1403),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_R g1556 ( 
.A(n_1381),
.B(n_315),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1331),
.Y(n_1557)
);

A2O1A1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1360),
.A2(n_1391),
.B(n_1406),
.C(n_1365),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1333),
.A2(n_325),
.B(n_326),
.C(n_328),
.Y(n_1559)
);

NOR3xp33_ASAP7_75t_SL g1560 ( 
.A(n_1227),
.B(n_370),
.C(n_329),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1224),
.B(n_1388),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1361),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1284),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1198),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1351),
.A2(n_335),
.B1(n_337),
.B2(n_341),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1287),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1264),
.A2(n_344),
.B1(n_346),
.B2(n_351),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1380),
.B(n_1294),
.Y(n_1568)
);

NAND2x1p5_ASAP7_75t_L g1569 ( 
.A(n_1304),
.B(n_353),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1319),
.A2(n_354),
.B(n_356),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1335),
.B(n_1364),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_L g1572 ( 
.A1(n_1407),
.A2(n_360),
.B(n_1309),
.C(n_1240),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1386),
.Y(n_1573)
);

A2O1A1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1396),
.A2(n_1404),
.B(n_1402),
.C(n_1368),
.Y(n_1574)
);

NOR3xp33_ASAP7_75t_SL g1575 ( 
.A(n_1344),
.B(n_1211),
.C(n_1303),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1359),
.B(n_1387),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1287),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_SL g1578 ( 
.A1(n_1397),
.A2(n_1400),
.B1(n_1353),
.B2(n_1395),
.Y(n_1578)
);

AO21x1_ASAP7_75t_L g1579 ( 
.A1(n_1261),
.A2(n_1312),
.B(n_1280),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1379),
.B(n_1376),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1357),
.Y(n_1581)
);

NOR3xp33_ASAP7_75t_SL g1582 ( 
.A(n_1265),
.B(n_1266),
.C(n_1399),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1376),
.B(n_1261),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1252),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1405),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1354),
.A2(n_1394),
.B1(n_1367),
.B2(n_1218),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1199),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1338),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1199),
.A2(n_1210),
.B(n_1254),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1210),
.B(n_1254),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1259),
.B(n_1298),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_R g1592 ( 
.A(n_1304),
.B(n_1356),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1257),
.A2(n_1296),
.B1(n_1283),
.B2(n_1298),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1259),
.A2(n_1290),
.B1(n_1292),
.B2(n_1337),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1257),
.A2(n_1283),
.B(n_1296),
.Y(n_1595)
);

AOI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1329),
.A2(n_1283),
.B(n_1296),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1337),
.A2(n_1345),
.B(n_1346),
.C(n_1354),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1329),
.A2(n_1242),
.B(n_1010),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1349),
.A2(n_1242),
.B(n_1010),
.Y(n_1599)
);

OA22x2_ASAP7_75t_L g1600 ( 
.A1(n_1349),
.A2(n_1076),
.B1(n_1039),
.B2(n_1027),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1221),
.Y(n_1601)
);

BUFx8_ASAP7_75t_SL g1602 ( 
.A(n_1274),
.Y(n_1602)
);

NOR2xp67_ASAP7_75t_L g1603 ( 
.A(n_1223),
.B(n_1250),
.Y(n_1603)
);

AOI33xp33_ASAP7_75t_L g1604 ( 
.A1(n_1215),
.A2(n_1267),
.A3(n_1177),
.B1(n_997),
.B2(n_1049),
.B3(n_1268),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1242),
.B(n_976),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1242),
.A2(n_1225),
.B(n_1310),
.C(n_1307),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1390),
.B(n_985),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1221),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1207),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1242),
.A2(n_1010),
.B(n_1002),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_SL g1611 ( 
.A(n_1226),
.B(n_1002),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1242),
.B(n_976),
.Y(n_1612)
);

O2A1O1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1242),
.A2(n_1225),
.B(n_1310),
.C(n_1307),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1242),
.A2(n_1006),
.B(n_1007),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1242),
.A2(n_1010),
.B(n_1002),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1242),
.B(n_976),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_R g1617 ( 
.A(n_1334),
.B(n_979),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1242),
.B(n_976),
.Y(n_1618)
);

AND2x6_ASAP7_75t_SL g1619 ( 
.A(n_1274),
.B(n_1000),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1208),
.B(n_1173),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1288),
.B(n_985),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1288),
.B(n_985),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1288),
.B(n_933),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1242),
.A2(n_1311),
.B1(n_1328),
.B2(n_1327),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1221),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1242),
.B(n_976),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1293),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1288),
.B(n_985),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1207),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1242),
.A2(n_1311),
.B1(n_1328),
.B2(n_1327),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1242),
.A2(n_1010),
.B(n_1002),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1242),
.A2(n_1311),
.B1(n_1328),
.B2(n_1327),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1219),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1608),
.Y(n_1634)
);

BUFx2_ASAP7_75t_R g1635 ( 
.A(n_1602),
.Y(n_1635)
);

BUFx2_ASAP7_75t_R g1636 ( 
.A(n_1437),
.Y(n_1636)
);

AO21x2_ASAP7_75t_L g1637 ( 
.A1(n_1514),
.A2(n_1411),
.B(n_1574),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1414),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1595),
.A2(n_1615),
.B(n_1610),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1631),
.A2(n_1598),
.B(n_1599),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1420),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1614),
.A2(n_1613),
.B(n_1606),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1425),
.Y(n_1643)
);

BUFx4f_ASAP7_75t_SL g1644 ( 
.A(n_1444),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1432),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1617),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1623),
.B(n_1451),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1428),
.Y(n_1648)
);

AOI22x1_ASAP7_75t_L g1649 ( 
.A1(n_1461),
.A2(n_1569),
.B1(n_1464),
.B2(n_1450),
.Y(n_1649)
);

BUFx8_ASAP7_75t_L g1650 ( 
.A(n_1478),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1503),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1531),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1624),
.A2(n_1632),
.B(n_1630),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1451),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1605),
.B(n_1612),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1498),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1429),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1442),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1540),
.A2(n_1593),
.B(n_1570),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1501),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1609),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1500),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1452),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1601),
.Y(n_1664)
);

NAND2x1p5_ASAP7_75t_L g1665 ( 
.A(n_1487),
.B(n_1510),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1500),
.Y(n_1666)
);

AO21x2_ASAP7_75t_L g1667 ( 
.A1(n_1489),
.A2(n_1597),
.B(n_1579),
.Y(n_1667)
);

BUFx12f_ASAP7_75t_L g1668 ( 
.A(n_1440),
.Y(n_1668)
);

INVx5_ASAP7_75t_L g1669 ( 
.A(n_1590),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1498),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1620),
.B(n_1616),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1492),
.Y(n_1672)
);

BUFx5_ASAP7_75t_L g1673 ( 
.A(n_1516),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1629),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1625),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1578),
.A2(n_1462),
.B1(n_1600),
.B2(n_1562),
.Y(n_1676)
);

AO21x2_ASAP7_75t_L g1677 ( 
.A1(n_1435),
.A2(n_1558),
.B(n_1532),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1607),
.B(n_1618),
.Y(n_1678)
);

INVx4_ASAP7_75t_L g1679 ( 
.A(n_1531),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1455),
.Y(n_1680)
);

AO21x2_ASAP7_75t_L g1681 ( 
.A1(n_1435),
.A2(n_1422),
.B(n_1408),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1488),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1434),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1492),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1430),
.Y(n_1685)
);

INVx4_ASAP7_75t_L g1686 ( 
.A(n_1535),
.Y(n_1686)
);

AO21x2_ASAP7_75t_L g1687 ( 
.A1(n_1454),
.A2(n_1466),
.B(n_1559),
.Y(n_1687)
);

AO21x2_ASAP7_75t_L g1688 ( 
.A1(n_1459),
.A2(n_1502),
.B(n_1443),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1529),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1533),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1470),
.A2(n_1552),
.B1(n_1525),
.B2(n_1556),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1536),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_SL g1693 ( 
.A1(n_1493),
.A2(n_1491),
.B1(n_1537),
.B2(n_1546),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1607),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1626),
.B(n_1508),
.Y(n_1695)
);

BUFx8_ASAP7_75t_L g1696 ( 
.A(n_1633),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1538),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1508),
.B(n_1534),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1458),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1409),
.Y(n_1700)
);

OAI21x1_ASAP7_75t_SL g1701 ( 
.A1(n_1545),
.A2(n_1467),
.B(n_1565),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1527),
.Y(n_1702)
);

BUFx2_ASAP7_75t_SL g1703 ( 
.A(n_1603),
.Y(n_1703)
);

BUFx8_ASAP7_75t_L g1704 ( 
.A(n_1627),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1446),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1578),
.A2(n_1499),
.B1(n_1457),
.B2(n_1576),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1590),
.Y(n_1707)
);

INVx6_ASAP7_75t_L g1708 ( 
.A(n_1409),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_1416),
.Y(n_1709)
);

AO21x2_ASAP7_75t_L g1710 ( 
.A1(n_1441),
.A2(n_1473),
.B(n_1471),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1572),
.A2(n_1419),
.B(n_1553),
.Y(n_1711)
);

OAI21x1_ASAP7_75t_SL g1712 ( 
.A1(n_1565),
.A2(n_1550),
.B(n_1567),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1549),
.A2(n_1484),
.B1(n_1507),
.B2(n_1497),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1544),
.Y(n_1714)
);

AO21x2_ASAP7_75t_L g1715 ( 
.A1(n_1476),
.A2(n_1483),
.B(n_1477),
.Y(n_1715)
);

AO21x2_ASAP7_75t_L g1716 ( 
.A1(n_1490),
.A2(n_1494),
.B(n_1567),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1542),
.B(n_1543),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1548),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1573),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1517),
.A2(n_1588),
.B(n_1496),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1555),
.Y(n_1721)
);

AOI22x1_ASAP7_75t_L g1722 ( 
.A1(n_1541),
.A2(n_1551),
.B1(n_1547),
.B2(n_1520),
.Y(n_1722)
);

AO21x2_ASAP7_75t_L g1723 ( 
.A1(n_1519),
.A2(n_1521),
.B(n_1474),
.Y(n_1723)
);

INVx8_ASAP7_75t_L g1724 ( 
.A(n_1619),
.Y(n_1724)
);

INVx8_ASAP7_75t_L g1725 ( 
.A(n_1619),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1515),
.B(n_1491),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1539),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1424),
.A2(n_1412),
.B(n_1433),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1453),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1486),
.B(n_1482),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1585),
.Y(n_1731)
);

AO21x2_ASAP7_75t_L g1732 ( 
.A1(n_1523),
.A2(n_1526),
.B(n_1568),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1557),
.B(n_1460),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1426),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1447),
.Y(n_1735)
);

INVx4_ASAP7_75t_L g1736 ( 
.A(n_1581),
.Y(n_1736)
);

AO21x2_ASAP7_75t_L g1737 ( 
.A1(n_1513),
.A2(n_1445),
.B(n_1439),
.Y(n_1737)
);

INVxp67_ASAP7_75t_SL g1738 ( 
.A(n_1512),
.Y(n_1738)
);

BUFx2_ASAP7_75t_SL g1739 ( 
.A(n_1485),
.Y(n_1739)
);

OR2x6_ASAP7_75t_L g1740 ( 
.A(n_1438),
.B(n_1449),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1582),
.B(n_1431),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1530),
.A2(n_1472),
.B1(n_1522),
.B2(n_1576),
.Y(n_1742)
);

INVx8_ASAP7_75t_L g1743 ( 
.A(n_1564),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1554),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1604),
.B(n_1421),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1413),
.B(n_1575),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1431),
.B(n_1417),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1511),
.A2(n_1506),
.B1(n_1456),
.B2(n_1481),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1475),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1423),
.B(n_1418),
.Y(n_1750)
);

OAI21x1_ASAP7_75t_L g1751 ( 
.A1(n_1586),
.A2(n_1591),
.B(n_1580),
.Y(n_1751)
);

INVx6_ASAP7_75t_L g1752 ( 
.A(n_1530),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1583),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1415),
.B(n_1495),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1571),
.B(n_1524),
.Y(n_1755)
);

INVx4_ASAP7_75t_L g1756 ( 
.A(n_1564),
.Y(n_1756)
);

OA21x2_ASAP7_75t_L g1757 ( 
.A1(n_1436),
.A2(n_1560),
.B(n_1551),
.Y(n_1757)
);

AOI22x1_ASAP7_75t_L g1758 ( 
.A1(n_1479),
.A2(n_1509),
.B1(n_1504),
.B2(n_1584),
.Y(n_1758)
);

CKINVDCx11_ASAP7_75t_R g1759 ( 
.A(n_1587),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1561),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1427),
.B(n_1410),
.Y(n_1761)
);

INVx6_ASAP7_75t_SL g1762 ( 
.A(n_1465),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1448),
.Y(n_1763)
);

OAI21x1_ASAP7_75t_L g1764 ( 
.A1(n_1594),
.A2(n_1528),
.B(n_1463),
.Y(n_1764)
);

BUFx12f_ASAP7_75t_L g1765 ( 
.A(n_1563),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1621),
.Y(n_1766)
);

INVx4_ASAP7_75t_L g1767 ( 
.A(n_1566),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1622),
.Y(n_1768)
);

NAND2x1p5_ASAP7_75t_L g1769 ( 
.A(n_1577),
.B(n_1628),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1505),
.B(n_1468),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1592),
.Y(n_1771)
);

OR2x6_ASAP7_75t_L g1772 ( 
.A(n_1518),
.B(n_1611),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1518),
.Y(n_1773)
);

INVx5_ASAP7_75t_L g1774 ( 
.A(n_1469),
.Y(n_1774)
);

OAI21x1_ASAP7_75t_L g1775 ( 
.A1(n_1469),
.A2(n_1596),
.B(n_1589),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1480),
.Y(n_1776)
);

NAND2x1p5_ASAP7_75t_L g1777 ( 
.A(n_1487),
.B(n_1510),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1492),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1428),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1425),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1451),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1623),
.B(n_933),
.Y(n_1782)
);

BUFx2_ASAP7_75t_SL g1783 ( 
.A(n_1501),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1451),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1428),
.Y(n_1785)
);

BUFx4f_ASAP7_75t_L g1786 ( 
.A(n_1444),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1492),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1425),
.Y(n_1788)
);

BUFx3_ASAP7_75t_L g1789 ( 
.A(n_1428),
.Y(n_1789)
);

INVx8_ASAP7_75t_L g1790 ( 
.A(n_1602),
.Y(n_1790)
);

AO21x2_ASAP7_75t_L g1791 ( 
.A1(n_1514),
.A2(n_1214),
.B(n_1411),
.Y(n_1791)
);

INVx2_ASAP7_75t_SL g1792 ( 
.A(n_1498),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1425),
.B(n_1607),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1428),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1655),
.B(n_1782),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1717),
.Y(n_1796)
);

OR2x6_ASAP7_75t_L g1797 ( 
.A(n_1652),
.B(n_1679),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1759),
.Y(n_1798)
);

CKINVDCx6p67_ASAP7_75t_R g1799 ( 
.A(n_1790),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1717),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1706),
.A2(n_1755),
.B1(n_1671),
.B2(n_1676),
.Y(n_1801)
);

CKINVDCx20_ASAP7_75t_R g1802 ( 
.A(n_1650),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1704),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1671),
.B(n_1746),
.Y(n_1804)
);

INVx2_ASAP7_75t_SL g1805 ( 
.A(n_1704),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1706),
.A2(n_1676),
.B1(n_1701),
.B2(n_1724),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1776),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1724),
.A2(n_1725),
.B1(n_1770),
.B2(n_1652),
.Y(n_1808)
);

INVx8_ASAP7_75t_L g1809 ( 
.A(n_1790),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1678),
.B(n_1761),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1638),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1724),
.A2(n_1725),
.B1(n_1679),
.B2(n_1643),
.Y(n_1812)
);

BUFx3_ASAP7_75t_L g1813 ( 
.A(n_1699),
.Y(n_1813)
);

OA21x2_ASAP7_75t_L g1814 ( 
.A1(n_1775),
.A2(n_1653),
.B(n_1642),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1684),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1759),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1790),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1725),
.A2(n_1780),
.B1(n_1788),
.B2(n_1643),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1780),
.A2(n_1788),
.B1(n_1742),
.B2(n_1691),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1641),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1650),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1642),
.B(n_1745),
.Y(n_1822)
);

NAND2x1p5_ASAP7_75t_L g1823 ( 
.A(n_1771),
.B(n_1684),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1647),
.B(n_1678),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1761),
.A2(n_1722),
.B1(n_1713),
.B2(n_1748),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1748),
.A2(n_1713),
.B1(n_1754),
.B2(n_1711),
.Y(n_1826)
);

BUFx12f_ASAP7_75t_L g1827 ( 
.A(n_1646),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1662),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1645),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1762),
.A2(n_1793),
.B1(n_1693),
.B2(n_1695),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1658),
.Y(n_1831)
);

CKINVDCx20_ASAP7_75t_R g1832 ( 
.A(n_1721),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1685),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_SL g1834 ( 
.A1(n_1712),
.A2(n_1774),
.B1(n_1739),
.B2(n_1793),
.Y(n_1834)
);

AO21x2_ASAP7_75t_L g1835 ( 
.A1(n_1791),
.A2(n_1677),
.B(n_1749),
.Y(n_1835)
);

INVx4_ASAP7_75t_L g1836 ( 
.A(n_1644),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1663),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1762),
.A2(n_1693),
.B1(n_1695),
.B2(n_1741),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1664),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1675),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1760),
.B(n_1654),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1711),
.A2(n_1745),
.B1(n_1742),
.B2(n_1728),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1672),
.B(n_1778),
.Y(n_1843)
);

BUFx4_ASAP7_75t_SL g1844 ( 
.A(n_1740),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1786),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1635),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1662),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1691),
.A2(n_1741),
.B1(n_1747),
.B2(n_1774),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1689),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1690),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1654),
.B(n_1781),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1692),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1784),
.Y(n_1853)
);

NAND2x1p5_ASAP7_75t_L g1854 ( 
.A(n_1771),
.B(n_1672),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1786),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1772),
.A2(n_1774),
.B1(n_1651),
.B2(n_1698),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1634),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1743),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1697),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1747),
.A2(n_1710),
.B1(n_1715),
.B2(n_1726),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1710),
.A2(n_1715),
.B1(n_1757),
.B2(n_1753),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1696),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1718),
.B(n_1719),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1680),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1682),
.B(n_1637),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1657),
.Y(n_1866)
);

BUFx4f_ASAP7_75t_SL g1867 ( 
.A(n_1721),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1637),
.B(n_1732),
.Y(n_1868)
);

OAI21x1_ASAP7_75t_L g1869 ( 
.A1(n_1659),
.A2(n_1640),
.B(n_1639),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1772),
.A2(n_1773),
.B1(n_1657),
.B2(n_1744),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1757),
.A2(n_1750),
.B1(n_1714),
.B2(n_1732),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1743),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1772),
.A2(n_1773),
.B1(n_1744),
.B2(n_1666),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1648),
.Y(n_1874)
);

BUFx2_ASAP7_75t_R g1875 ( 
.A(n_1646),
.Y(n_1875)
);

INVx2_ASAP7_75t_SL g1876 ( 
.A(n_1740),
.Y(n_1876)
);

INVx4_ASAP7_75t_L g1877 ( 
.A(n_1644),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1694),
.B(n_1787),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1731),
.B(n_1673),
.Y(n_1879)
);

AOI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1750),
.A2(n_1768),
.B1(n_1766),
.B2(n_1696),
.Y(n_1880)
);

INVx3_ASAP7_75t_L g1881 ( 
.A(n_1686),
.Y(n_1881)
);

NAND2x1p5_ASAP7_75t_L g1882 ( 
.A(n_1669),
.B(n_1686),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1734),
.B(n_1735),
.Y(n_1883)
);

CKINVDCx20_ASAP7_75t_R g1884 ( 
.A(n_1683),
.Y(n_1884)
);

BUFx10_ASAP7_75t_L g1885 ( 
.A(n_1740),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1666),
.Y(n_1886)
);

AO21x2_ASAP7_75t_L g1887 ( 
.A1(n_1791),
.A2(n_1677),
.B(n_1667),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1660),
.B(n_1730),
.Y(n_1888)
);

OAI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1669),
.A2(n_1769),
.B1(n_1767),
.B2(n_1777),
.Y(n_1889)
);

CKINVDCx20_ASAP7_75t_R g1890 ( 
.A(n_1683),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1733),
.B(n_1783),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1795),
.B(n_1648),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1801),
.A2(n_1765),
.B1(n_1737),
.B2(n_1716),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1824),
.B(n_1661),
.Y(n_1894)
);

NOR3xp33_ASAP7_75t_SL g1895 ( 
.A(n_1846),
.B(n_1763),
.C(n_1635),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1866),
.B(n_1767),
.Y(n_1896)
);

CKINVDCx8_ASAP7_75t_R g1897 ( 
.A(n_1809),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1826),
.A2(n_1806),
.B1(n_1825),
.B2(n_1819),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_SL g1899 ( 
.A1(n_1819),
.A2(n_1673),
.B1(n_1752),
.B2(n_1708),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1807),
.Y(n_1900)
);

AO21x2_ASAP7_75t_L g1901 ( 
.A1(n_1869),
.A2(n_1667),
.B(n_1681),
.Y(n_1901)
);

NOR2x1_ASAP7_75t_L g1902 ( 
.A(n_1881),
.B(n_1700),
.Y(n_1902)
);

OR2x6_ASAP7_75t_L g1903 ( 
.A(n_1797),
.B(n_1703),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1863),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1828),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1822),
.B(n_1796),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1828),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1797),
.B(n_1707),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1804),
.B(n_1661),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1841),
.B(n_1674),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1847),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1810),
.B(n_1674),
.Y(n_1912)
);

AO32x2_ASAP7_75t_L g1913 ( 
.A1(n_1873),
.A2(n_1700),
.A3(n_1729),
.B1(n_1756),
.B2(n_1705),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1851),
.B(n_1779),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1883),
.B(n_1779),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_SL g1916 ( 
.A1(n_1867),
.A2(n_1709),
.B1(n_1763),
.B2(n_1668),
.Y(n_1916)
);

NAND2xp33_ASAP7_75t_R g1917 ( 
.A(n_1862),
.B(n_1636),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1822),
.B(n_1720),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1806),
.A2(n_1737),
.B1(n_1687),
.B2(n_1758),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1797),
.B(n_1707),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1800),
.B(n_1673),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1811),
.Y(n_1922)
);

NOR3xp33_ASAP7_75t_SL g1923 ( 
.A(n_1821),
.B(n_1636),
.C(n_1738),
.Y(n_1923)
);

BUFx6f_ASAP7_75t_SL g1924 ( 
.A(n_1803),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1866),
.B(n_1794),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1826),
.B(n_1673),
.Y(n_1926)
);

NAND2xp33_ASAP7_75t_R g1927 ( 
.A(n_1881),
.B(n_1702),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1820),
.Y(n_1928)
);

INVx4_ASAP7_75t_L g1929 ( 
.A(n_1809),
.Y(n_1929)
);

INVx4_ASAP7_75t_L g1930 ( 
.A(n_1809),
.Y(n_1930)
);

NAND2xp33_ASAP7_75t_R g1931 ( 
.A(n_1844),
.B(n_1702),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1847),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1829),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1802),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1799),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1886),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1838),
.A2(n_1687),
.B1(n_1673),
.B2(n_1723),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1813),
.B(n_1794),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1831),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1805),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1842),
.B(n_1688),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1832),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1853),
.B(n_1789),
.Y(n_1943)
);

CKINVDCx20_ASAP7_75t_R g1944 ( 
.A(n_1867),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1874),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1858),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1837),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1839),
.Y(n_1948)
);

INVxp67_ASAP7_75t_L g1949 ( 
.A(n_1886),
.Y(n_1949)
);

OR2x6_ASAP7_75t_L g1950 ( 
.A(n_1882),
.B(n_1665),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1844),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1884),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1840),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1830),
.A2(n_1723),
.B1(n_1688),
.B2(n_1708),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1890),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1842),
.B(n_1751),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1836),
.B(n_1792),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1860),
.B(n_1738),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1817),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1853),
.B(n_1789),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1836),
.B(n_1670),
.Y(n_1961)
);

CKINVDCx20_ASAP7_75t_R g1962 ( 
.A(n_1877),
.Y(n_1962)
);

AOI22xp33_ASAP7_75t_L g1963 ( 
.A1(n_1888),
.A2(n_1708),
.B1(n_1752),
.B2(n_1764),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1885),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1857),
.B(n_1785),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1879),
.B(n_1727),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1860),
.B(n_1861),
.Y(n_1967)
);

AOI22xp33_ASAP7_75t_L g1968 ( 
.A1(n_1818),
.A2(n_1769),
.B1(n_1785),
.B2(n_1649),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1918),
.B(n_1814),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1918),
.B(n_1814),
.Y(n_1970)
);

AND2x4_ASAP7_75t_SL g1971 ( 
.A(n_1903),
.B(n_1885),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1913),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1905),
.B(n_1865),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1907),
.B(n_1868),
.Y(n_1974)
);

OAI31xp33_ASAP7_75t_L g1975 ( 
.A1(n_1898),
.A2(n_1818),
.A3(n_1889),
.B(n_1823),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1913),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1911),
.B(n_1871),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1911),
.Y(n_1978)
);

INVxp67_ASAP7_75t_L g1979 ( 
.A(n_1932),
.Y(n_1979)
);

NAND5xp2_ASAP7_75t_L g1980 ( 
.A(n_1895),
.B(n_1808),
.C(n_1812),
.D(n_1848),
.E(n_1834),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1906),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1932),
.B(n_1887),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1898),
.A2(n_1848),
.B1(n_1834),
.B2(n_1891),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1900),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1922),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1936),
.B(n_1887),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1936),
.B(n_1967),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1928),
.Y(n_1988)
);

NOR2x1_ASAP7_75t_SL g1989 ( 
.A(n_1903),
.B(n_1856),
.Y(n_1989)
);

BUFx2_ASAP7_75t_L g1990 ( 
.A(n_1913),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1967),
.B(n_1835),
.Y(n_1991)
);

BUFx2_ASAP7_75t_L g1992 ( 
.A(n_1966),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1933),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1939),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1947),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1949),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1949),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1926),
.B(n_1870),
.Y(n_1998)
);

AOI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1899),
.A2(n_1808),
.B1(n_1798),
.B2(n_1816),
.Y(n_1999)
);

NOR2x1_ASAP7_75t_L g2000 ( 
.A(n_1903),
.B(n_1873),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1948),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1952),
.B(n_1877),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1896),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1926),
.B(n_1879),
.Y(n_2004)
);

INVx2_ASAP7_75t_SL g2005 ( 
.A(n_1950),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1953),
.B(n_1835),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1904),
.B(n_1849),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_2006),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1984),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_2003),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1981),
.B(n_1925),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1991),
.B(n_1941),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1985),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1989),
.B(n_1958),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2006),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1987),
.B(n_1943),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1991),
.B(n_1987),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1985),
.B(n_1960),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1988),
.B(n_1914),
.Y(n_2019)
);

AND2x4_ASAP7_75t_SL g2020 ( 
.A(n_2005),
.B(n_1929),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1993),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1993),
.B(n_1910),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1974),
.B(n_1956),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1969),
.B(n_1970),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1994),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1974),
.B(n_1956),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1995),
.B(n_1915),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1969),
.B(n_1901),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_2004),
.B(n_1921),
.Y(n_2029)
);

INVxp67_ASAP7_75t_L g2030 ( 
.A(n_1992),
.Y(n_2030)
);

INVx2_ASAP7_75t_SL g2031 ( 
.A(n_2005),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_2024),
.B(n_2017),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2024),
.B(n_1970),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_2017),
.B(n_1982),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2012),
.B(n_1973),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2012),
.B(n_2008),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2028),
.B(n_1982),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2028),
.B(n_2008),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_2020),
.B(n_2000),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2015),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2015),
.B(n_1973),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2016),
.B(n_1986),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_2014),
.A2(n_1980),
.B1(n_1975),
.B2(n_1983),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_2009),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_2023),
.B(n_1986),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2013),
.Y(n_2046)
);

HB1xp67_ASAP7_75t_L g2047 ( 
.A(n_2010),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2023),
.B(n_1977),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_2014),
.A2(n_1980),
.B1(n_1975),
.B2(n_1899),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_2026),
.B(n_1998),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2026),
.B(n_1977),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2014),
.B(n_1998),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_2050),
.B(n_2011),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2046),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_2050),
.B(n_2029),
.Y(n_2055)
);

NOR2xp67_ASAP7_75t_L g2056 ( 
.A(n_2039),
.B(n_1929),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_2052),
.B(n_2000),
.Y(n_2057)
);

OAI31xp33_ASAP7_75t_L g2058 ( 
.A1(n_2043),
.A2(n_2020),
.A3(n_1971),
.B(n_2005),
.Y(n_2058)
);

INVxp67_ASAP7_75t_L g2059 ( 
.A(n_2047),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_2044),
.Y(n_2060)
);

OAI21xp33_ASAP7_75t_SL g2061 ( 
.A1(n_2032),
.A2(n_2031),
.B(n_2030),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2034),
.B(n_2031),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_2035),
.B(n_2029),
.Y(n_2063)
);

INVx2_ASAP7_75t_SL g2064 ( 
.A(n_2032),
.Y(n_2064)
);

OAI221xp5_ASAP7_75t_L g2065 ( 
.A1(n_2049),
.A2(n_1897),
.B1(n_1917),
.B2(n_1895),
.C(n_1999),
.Y(n_2065)
);

INVx1_ASAP7_75t_SL g2066 ( 
.A(n_2033),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_2035),
.B(n_2018),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2040),
.B(n_2021),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_2036),
.B(n_2022),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2040),
.B(n_2025),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2048),
.B(n_2051),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2034),
.B(n_2033),
.Y(n_2072)
);

NAND2x2_ASAP7_75t_L g2073 ( 
.A(n_2036),
.B(n_1940),
.Y(n_2073)
);

OAI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_2073),
.A2(n_1990),
.B1(n_1976),
.B2(n_1972),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2055),
.Y(n_2075)
);

OAI211xp5_ASAP7_75t_SL g2076 ( 
.A1(n_2065),
.A2(n_1923),
.B(n_1812),
.C(n_1963),
.Y(n_2076)
);

O2A1O1Ixp33_ASAP7_75t_L g2077 ( 
.A1(n_2065),
.A2(n_2002),
.B(n_1845),
.C(n_1855),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2059),
.B(n_2048),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2064),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_2073),
.A2(n_1892),
.B1(n_1971),
.B2(n_1909),
.Y(n_2080)
);

AOI21xp5_ASAP7_75t_L g2081 ( 
.A1(n_2061),
.A2(n_1989),
.B(n_1971),
.Y(n_2081)
);

OAI21xp33_ASAP7_75t_L g2082 ( 
.A1(n_2057),
.A2(n_2052),
.B(n_2051),
.Y(n_2082)
);

XNOR2x1_ASAP7_75t_L g2083 ( 
.A(n_2056),
.B(n_1955),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2060),
.Y(n_2084)
);

AOI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_2057),
.A2(n_2045),
.B1(n_2037),
.B2(n_2038),
.Y(n_2085)
);

INVx4_ASAP7_75t_L g2086 ( 
.A(n_2060),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2068),
.Y(n_2087)
);

INVx2_ASAP7_75t_SL g2088 ( 
.A(n_2062),
.Y(n_2088)
);

AOI221xp5_ASAP7_75t_L g2089 ( 
.A1(n_2074),
.A2(n_2059),
.B1(n_2058),
.B2(n_2066),
.C(n_2054),
.Y(n_2089)
);

INVx3_ASAP7_75t_L g2090 ( 
.A(n_2086),
.Y(n_2090)
);

INVx1_ASAP7_75t_SL g2091 ( 
.A(n_2083),
.Y(n_2091)
);

NAND3xp33_ASAP7_75t_L g2092 ( 
.A(n_2077),
.B(n_1923),
.C(n_1893),
.Y(n_2092)
);

INVx2_ASAP7_75t_SL g2093 ( 
.A(n_2079),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_2076),
.A2(n_1972),
.B1(n_1976),
.B2(n_1990),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2085),
.B(n_2072),
.Y(n_2095)
);

OAI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_2081),
.A2(n_1902),
.B(n_2071),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2075),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2088),
.B(n_2071),
.Y(n_2098)
);

OAI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2080),
.A2(n_1962),
.B(n_1919),
.Y(n_2099)
);

OAI211xp5_ASAP7_75t_SL g2100 ( 
.A1(n_2080),
.A2(n_1880),
.B(n_1968),
.C(n_1954),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2087),
.B(n_2078),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_2086),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_2082),
.B(n_1924),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2084),
.B(n_2053),
.Y(n_2104)
);

OAI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_2080),
.A2(n_2063),
.B1(n_2069),
.B2(n_2067),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2097),
.Y(n_2106)
);

OAI322xp33_ASAP7_75t_L g2107 ( 
.A1(n_2091),
.A2(n_2102),
.A3(n_2105),
.B1(n_2103),
.B2(n_2093),
.C1(n_2101),
.C2(n_2090),
.Y(n_2107)
);

AOI221xp5_ASAP7_75t_L g2108 ( 
.A1(n_2089),
.A2(n_1924),
.B1(n_2068),
.B2(n_2070),
.C(n_2045),
.Y(n_2108)
);

NAND3xp33_ASAP7_75t_L g2109 ( 
.A(n_2094),
.B(n_1942),
.C(n_1934),
.Y(n_2109)
);

NOR2x1_ASAP7_75t_L g2110 ( 
.A(n_2090),
.B(n_1930),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2098),
.B(n_2042),
.Y(n_2111)
);

NAND3xp33_ASAP7_75t_L g2112 ( 
.A(n_2099),
.B(n_1816),
.C(n_1798),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2104),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2095),
.B(n_2042),
.Y(n_2114)
);

NOR3x1_ASAP7_75t_L g2115 ( 
.A(n_2096),
.B(n_1876),
.C(n_1656),
.Y(n_2115)
);

NOR3xp33_ASAP7_75t_L g2116 ( 
.A(n_2091),
.B(n_1916),
.C(n_1736),
.Y(n_2116)
);

NAND3xp33_ASAP7_75t_L g2117 ( 
.A(n_2092),
.B(n_1816),
.C(n_1798),
.Y(n_2117)
);

OAI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_2117),
.A2(n_2102),
.B(n_2100),
.Y(n_2118)
);

OAI21xp33_ASAP7_75t_SL g2119 ( 
.A1(n_2108),
.A2(n_1930),
.B(n_1950),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2106),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_2116),
.A2(n_2104),
.B1(n_1944),
.B2(n_1951),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_2110),
.B(n_1935),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2114),
.B(n_2037),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2113),
.Y(n_2124)
);

AOI21xp5_ASAP7_75t_L g2125 ( 
.A1(n_2107),
.A2(n_1959),
.B(n_2070),
.Y(n_2125)
);

NOR3xp33_ASAP7_75t_L g2126 ( 
.A(n_2112),
.B(n_1736),
.C(n_1957),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2111),
.Y(n_2127)
);

OAI21xp33_ASAP7_75t_L g2128 ( 
.A1(n_2109),
.A2(n_1833),
.B(n_1945),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2115),
.B(n_2038),
.Y(n_2129)
);

AOI221xp5_ASAP7_75t_SL g2130 ( 
.A1(n_2125),
.A2(n_1709),
.B1(n_1938),
.B2(n_1961),
.C(n_1912),
.Y(n_2130)
);

AOI321xp33_ASAP7_75t_L g2131 ( 
.A1(n_2124),
.A2(n_1964),
.A3(n_1965),
.B1(n_1894),
.B2(n_1937),
.C(n_1908),
.Y(n_2131)
);

AOI221xp5_ASAP7_75t_L g2132 ( 
.A1(n_2118),
.A2(n_2001),
.B1(n_2007),
.B2(n_1979),
.C(n_1997),
.Y(n_2132)
);

AOI221xp5_ASAP7_75t_L g2133 ( 
.A1(n_2120),
.A2(n_2119),
.B1(n_2127),
.B2(n_2122),
.C(n_2129),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2121),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2126),
.A2(n_1931),
.B1(n_1927),
.B2(n_1964),
.Y(n_2135)
);

OAI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_2123),
.A2(n_2041),
.B1(n_2027),
.B2(n_2019),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2128),
.Y(n_2137)
);

AOI221xp5_ASAP7_75t_L g2138 ( 
.A1(n_2124),
.A2(n_2007),
.B1(n_1979),
.B2(n_1997),
.C(n_1996),
.Y(n_2138)
);

AND2x2_ASAP7_75t_SL g2139 ( 
.A(n_2137),
.B(n_2134),
.Y(n_2139)
);

INVx2_ASAP7_75t_SL g2140 ( 
.A(n_2135),
.Y(n_2140)
);

AOI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_2130),
.A2(n_1827),
.B1(n_1920),
.B2(n_1908),
.Y(n_2141)
);

INVxp67_ASAP7_75t_SL g2142 ( 
.A(n_2133),
.Y(n_2142)
);

OAI22x1_ASAP7_75t_L g2143 ( 
.A1(n_2131),
.A2(n_1823),
.B1(n_1875),
.B2(n_1854),
.Y(n_2143)
);

NOR2x1_ASAP7_75t_L g2144 ( 
.A(n_2136),
.B(n_1875),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2139),
.Y(n_2145)
);

XNOR2x1_ASAP7_75t_L g2146 ( 
.A(n_2144),
.B(n_1854),
.Y(n_2146)
);

NOR3xp33_ASAP7_75t_L g2147 ( 
.A(n_2142),
.B(n_2132),
.C(n_2138),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2140),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_2148),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_2145),
.Y(n_2150)
);

INVx2_ASAP7_75t_SL g2151 ( 
.A(n_2149),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2151),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2152),
.A2(n_2150),
.B1(n_2147),
.B2(n_2146),
.Y(n_2153)
);

OAI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_2153),
.A2(n_2141),
.B1(n_2143),
.B2(n_1950),
.Y(n_2154)
);

AOI21x1_ASAP7_75t_L g2155 ( 
.A1(n_2154),
.A2(n_1815),
.B(n_1878),
.Y(n_2155)
);

AOI222xp33_ASAP7_75t_L g2156 ( 
.A1(n_2155),
.A2(n_1843),
.B1(n_1852),
.B2(n_1859),
.C1(n_1850),
.C2(n_1864),
.Y(n_2156)
);

AOI221xp5_ASAP7_75t_R g2157 ( 
.A1(n_2156),
.A2(n_1996),
.B1(n_1978),
.B2(n_1777),
.C(n_1665),
.Y(n_2157)
);

AOI211xp5_ASAP7_75t_L g2158 ( 
.A1(n_2157),
.A2(n_1872),
.B(n_1858),
.C(n_1946),
.Y(n_2158)
);


endmodule