module fake_jpeg_30989_n_457 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_457);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_457;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_29),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_57),
.Y(n_110)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_53),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_85),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_55),
.Y(n_142)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_29),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_8),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_68),
.B(n_41),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_88),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_30),
.A2(n_37),
.B1(n_44),
.B2(n_32),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_38),
.B1(n_35),
.B2(n_48),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_94),
.Y(n_146)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_92),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_29),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_24),
.B1(n_45),
.B2(n_43),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_18),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_95),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_34),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_24),
.B1(n_41),
.B2(n_48),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_104),
.A2(n_113),
.B1(n_25),
.B2(n_27),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_78),
.A2(n_35),
.B1(n_38),
.B2(n_19),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_106),
.A2(n_137),
.B1(n_110),
.B2(n_146),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_131),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_145),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_46),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_130),
.B(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_28),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_46),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_45),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_135),
.B(n_139),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_84),
.A2(n_19),
.B1(n_26),
.B2(n_33),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_54),
.B(n_43),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_59),
.B(n_40),
.Y(n_143)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_52),
.B(n_40),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_60),
.B(n_33),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_150),
.Y(n_161)
);

AND2x4_ASAP7_75t_L g150 ( 
.A(n_91),
.B(n_26),
.Y(n_150)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_152),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_69),
.B1(n_61),
.B2(n_62),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_153),
.A2(n_192),
.B1(n_80),
.B2(n_101),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx5_ASAP7_75t_SL g212 ( 
.A(n_155),
.Y(n_212)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_27),
.A3(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_182),
.Y(n_209)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_163),
.Y(n_219)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_96),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_168),
.C(n_181),
.Y(n_217)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_135),
.B(n_94),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_169),
.B(n_173),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_170),
.B(n_174),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_92),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_141),
.Y(n_174)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_141),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_179),
.B(n_185),
.Y(n_220)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_55),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_184),
.Y(n_225)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_97),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_186),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_187),
.B(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_58),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_146),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_SL g191 ( 
.A(n_107),
.B(n_82),
.Y(n_191)
);

AOI22x1_ASAP7_75t_SL g232 ( 
.A1(n_191),
.A2(n_190),
.B1(n_173),
.B2(n_181),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_150),
.A2(n_65),
.B1(n_67),
.B2(n_71),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_193),
.B(n_125),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_70),
.B1(n_80),
.B2(n_22),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_146),
.B1(n_129),
.B2(n_105),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_59),
.B1(n_127),
.B2(n_124),
.Y(n_233)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_196),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_197),
.B(n_232),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_206),
.A2(n_138),
.B1(n_184),
.B2(n_177),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_141),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_213),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_158),
.B(n_102),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_215),
.A2(n_226),
.B1(n_229),
.B2(n_196),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_102),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_223),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_161),
.B(n_120),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_161),
.B(n_116),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_168),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_160),
.A2(n_129),
.B1(n_105),
.B2(n_134),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_160),
.A2(n_134),
.B1(n_133),
.B2(n_148),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_233),
.A2(n_172),
.B1(n_187),
.B2(n_191),
.Y(n_239)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_234),
.Y(n_274)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_242),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_239),
.A2(n_245),
.B1(n_247),
.B2(n_253),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_165),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_206),
.Y(n_278)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_248),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_160),
.B1(n_192),
.B2(n_165),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_231),
.A2(n_168),
.B1(n_172),
.B2(n_190),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_230),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_250),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_230),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_223),
.B(n_181),
.CI(n_173),
.CON(n_251),
.SN(n_251)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_251),
.B(n_262),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_224),
.A2(n_169),
.B1(n_183),
.B2(n_133),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_209),
.A2(n_231),
.B(n_232),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_249),
.B(n_246),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_256),
.A2(n_227),
.B1(n_136),
.B2(n_199),
.Y(n_295)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_259),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_208),
.A2(n_156),
.B1(n_151),
.B2(n_114),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_261),
.B1(n_264),
.B2(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_260),
.A2(n_225),
.B1(n_212),
.B2(n_230),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_231),
.A2(n_147),
.B1(n_140),
.B2(n_152),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_171),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_213),
.B(n_186),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_263),
.B(n_202),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_217),
.A2(n_147),
.B1(n_175),
.B2(n_162),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_166),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_204),
.C(n_103),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_197),
.A2(n_178),
.B1(n_154),
.B2(n_182),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_284),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_277),
.B1(n_289),
.B2(n_293),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_256),
.A2(n_215),
.B1(n_226),
.B2(n_229),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_283),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_200),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_288),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_198),
.C(n_202),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_285),
.C(n_251),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_200),
.B(n_205),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_282),
.A2(n_115),
.B(n_26),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_109),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_198),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_286),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_247),
.A2(n_210),
.A3(n_103),
.B1(n_136),
.B2(n_203),
.C1(n_222),
.C2(n_201),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_290),
.Y(n_298)
);

AO21x1_ASAP7_75t_L g288 ( 
.A1(n_246),
.A2(n_252),
.B(n_263),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_245),
.A2(n_204),
.B1(n_203),
.B2(n_201),
.Y(n_289)
);

NAND3xp33_ASAP7_75t_L g290 ( 
.A(n_235),
.B(n_222),
.C(n_1),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_214),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_216),
.Y(n_292)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_260),
.A2(n_227),
.B1(n_115),
.B2(n_216),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_295),
.A2(n_238),
.B1(n_127),
.B2(n_73),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_276),
.A2(n_241),
.B1(n_248),
.B2(n_250),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_299),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_292),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_310),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_267),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_273),
.A2(n_252),
.B(n_234),
.C(n_251),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_303),
.B(n_304),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_258),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_284),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_264),
.C(n_253),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_308),
.B(n_314),
.C(n_317),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_291),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_272),
.A2(n_239),
.B1(n_261),
.B2(n_266),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_312),
.A2(n_296),
.B1(n_274),
.B2(n_272),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_268),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_313),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_236),
.C(n_237),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_289),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_315),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_259),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_199),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_318),
.B(n_19),
.C(n_6),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_288),
.A2(n_257),
.B(n_242),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_319),
.A2(n_324),
.B(n_296),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_271),
.A2(n_155),
.B(n_121),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_320),
.A2(n_270),
.B(n_269),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_275),
.B(n_26),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_321),
.B(n_270),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_268),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_323),
.Y(n_343)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_326),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_315),
.A2(n_277),
.B1(n_293),
.B2(n_275),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_329),
.A2(n_339),
.B1(n_307),
.B2(n_323),
.Y(n_360)
);

OA21x2_ASAP7_75t_L g330 ( 
.A1(n_319),
.A2(n_267),
.B(n_279),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_322),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_331),
.A2(n_342),
.B(n_349),
.Y(n_369)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_347),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_314),
.B(n_274),
.Y(n_336)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_336),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_302),
.Y(n_341)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_341),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_307),
.A2(n_297),
.B1(n_238),
.B2(n_121),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_344),
.A2(n_351),
.B1(n_345),
.B2(n_331),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_297),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_121),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_350),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_11),
.B(n_1),
.Y(n_349)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_121),
.C(n_26),
.Y(n_350)
);

OAI21xp33_ASAP7_75t_SL g351 ( 
.A1(n_322),
.A2(n_11),
.B(n_4),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_311),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_317),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_374),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_360),
.A2(n_312),
.B1(n_330),
.B2(n_327),
.Y(n_393)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_362),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_318),
.C(n_308),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_375),
.C(n_324),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_365),
.A2(n_353),
.B1(n_345),
.B2(n_327),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_340),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_352),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_298),
.B1(n_309),
.B2(n_300),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_368),
.A2(n_371),
.B1(n_354),
.B2(n_357),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_310),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_372),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_339),
.A2(n_313),
.B1(n_301),
.B2(n_305),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_343),
.B(n_320),
.Y(n_373)
);

AOI221xp5_ASAP7_75t_L g384 ( 
.A1(n_373),
.A2(n_349),
.B1(n_335),
.B2(n_321),
.C(n_301),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_347),
.B(n_348),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_334),
.B(n_311),
.C(n_303),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_343),
.B(n_305),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_337),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_350),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_377),
.B(n_382),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_380),
.A2(n_393),
.B1(n_365),
.B2(n_369),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_371),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_342),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g383 ( 
.A(n_375),
.B(n_367),
.CI(n_362),
.CON(n_383),
.SN(n_383)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_383),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_384),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_329),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_388),
.Y(n_399)
);

XNOR2x1_ASAP7_75t_SL g389 ( 
.A(n_361),
.B(n_335),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g397 ( 
.A(n_389),
.B(n_374),
.CI(n_360),
.CON(n_397),
.SN(n_397)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_391),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_341),
.C(n_353),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_355),
.C(n_369),
.Y(n_398)
);

FAx1_ASAP7_75t_SL g394 ( 
.A(n_361),
.B(n_330),
.CI(n_333),
.CON(n_394),
.SN(n_394)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_394),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_393),
.A2(n_370),
.B(n_376),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_398),
.Y(n_417)
);

XOR2x2_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_382),
.Y(n_418)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_402),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_407),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_363),
.Y(n_404)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_385),
.A2(n_372),
.B1(n_386),
.B2(n_359),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_410),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_392),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_404),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_412),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_402),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_391),
.C(n_379),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_419),
.C(n_423),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_400),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_379),
.C(n_387),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g420 ( 
.A(n_395),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_399),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_366),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_421),
.B(n_394),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_383),
.C(n_377),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_416),
.A2(n_396),
.B1(n_405),
.B2(n_403),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_425),
.A2(n_430),
.B1(n_434),
.B2(n_12),
.Y(n_443)
);

AOI21x1_ASAP7_75t_L g442 ( 
.A1(n_426),
.A2(n_12),
.B(n_7),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_419),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_417),
.A2(n_399),
.B(n_397),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_429),
.B(n_433),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_422),
.A2(n_397),
.B1(n_338),
.B2(n_333),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_413),
.B(n_389),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_431),
.A2(n_11),
.B(n_6),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_400),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_326),
.C(n_19),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_435),
.B(n_418),
.C(n_423),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_436),
.B(n_438),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_424),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_439),
.A2(n_440),
.B(n_441),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_431),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_442),
.A2(n_434),
.B(n_7),
.Y(n_447)
);

O2A1O1Ixp33_ASAP7_75t_SL g444 ( 
.A1(n_443),
.A2(n_432),
.B(n_435),
.C(n_8),
.Y(n_444)
);

O2A1O1Ixp33_ASAP7_75t_SL g450 ( 
.A1(n_444),
.A2(n_447),
.B(n_448),
.C(n_12),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_437),
.A2(n_7),
.B(n_10),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_445),
.A2(n_438),
.B(n_440),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_449),
.A2(n_13),
.B(n_14),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_450),
.B(n_451),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_446),
.B(n_12),
.C(n_13),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_452),
.Y(n_454)
);

AOI321xp33_ASAP7_75t_L g455 ( 
.A1(n_454),
.A2(n_0),
.A3(n_15),
.B1(n_453),
.B2(n_437),
.C(n_420),
.Y(n_455)
);

AOI21x1_ASAP7_75t_L g456 ( 
.A1(n_455),
.A2(n_15),
.B(n_0),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_456),
.B(n_0),
.Y(n_457)
);


endmodule