module fake_jpeg_20099_n_185 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_33),
.B(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_30),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_37),
.B1(n_32),
.B2(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_48),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

AOI22x1_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_25),
.B1(n_18),
.B2(n_24),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_29),
.B(n_23),
.C(n_16),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_30),
.B1(n_27),
.B2(n_17),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_39),
.B1(n_2),
.B2(n_3),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_20),
.C(n_16),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_24),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx2_ASAP7_75t_SL g113 ( 
.A(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_79),
.B1(n_80),
.B2(n_52),
.Y(n_94)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_78),
.Y(n_92)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_83),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_26),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_44),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_28),
.B1(n_14),
.B2(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_14),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_10),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_13),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_39),
.C(n_52),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_112),
.C(n_73),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_110),
.B1(n_79),
.B2(n_74),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_54),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_109),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_108),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_71),
.A3(n_80),
.B1(n_76),
.B2(n_67),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_54),
.B1(n_4),
.B2(n_5),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_12),
.C(n_6),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_124),
.Y(n_144)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_122),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_66),
.B(n_83),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_112),
.B(n_97),
.Y(n_135)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_128),
.Y(n_138)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_68),
.B(n_84),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_65),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_70),
.B1(n_77),
.B2(n_12),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_99),
.B1(n_103),
.B2(n_93),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_90),
.B(n_91),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_110),
.B(n_98),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_77),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_1),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_6),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_1),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_140),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_143),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_102),
.C(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_150),
.Y(n_164)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_118),
.B1(n_126),
.B2(n_125),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_118),
.B1(n_125),
.B2(n_131),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_136),
.B(n_121),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_140),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_157),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_135),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_147),
.B(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_160),
.A2(n_151),
.B(n_154),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_143),
.C(n_144),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_132),
.C(n_119),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_155),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_166),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_163),
.B1(n_159),
.B2(n_160),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_148),
.C(n_150),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_170),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_149),
.C(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_164),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_141),
.B(n_8),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_117),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_161),
.A3(n_122),
.B1(n_169),
.B2(n_114),
.C1(n_123),
.C2(n_117),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_176),
.A2(n_175),
.B(n_172),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_177),
.A2(n_178),
.B1(n_116),
.B2(n_129),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_180),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_120),
.B(n_116),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_120),
.B(n_108),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_182),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_102),
.Y(n_185)
);


endmodule