module fake_jpeg_21233_n_141 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_SL g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_1),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_11),
.Y(n_36)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_13),
.B1(n_14),
.B2(n_19),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_13),
.B1(n_19),
.B2(n_16),
.Y(n_49)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_26),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_46),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_28),
.B(n_14),
.C(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_27),
.B1(n_29),
.B2(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_50),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_37),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_22),
.C(n_25),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_31),
.C(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_33),
.B(n_23),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_12),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_12),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_42),
.C(n_2),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_1),
.C(n_2),
.Y(n_97)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_80),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_52),
.Y(n_75)
);

OAI322xp33_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_11),
.A3(n_10),
.B1(n_18),
.B2(n_23),
.C1(n_21),
.C2(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_37),
.B1(n_29),
.B2(n_32),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_82),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_37),
.B1(n_29),
.B2(n_32),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_31),
.C(n_25),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_56),
.Y(n_94)
);

AOI21x1_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_66),
.B(n_57),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_82),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_57),
.B(n_10),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_92),
.B(n_93),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_94),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_65),
.B(n_63),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_18),
.B(n_21),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_72),
.Y(n_107)
);

AOI22x1_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_18),
.B1(n_26),
.B2(n_20),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_107),
.B(n_108),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_106),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_81),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_78),
.C(n_56),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_96),
.B(n_93),
.Y(n_114)
);

OAI21x1_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_116),
.B(n_117),
.Y(n_119)
);

AOI221xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_98),
.B1(n_96),
.B2(n_85),
.C(n_95),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_90),
.B(n_5),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_108),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_35),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_99),
.B1(n_106),
.B2(n_35),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_123),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_122),
.A2(n_116),
.B(n_6),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_35),
.B1(n_5),
.B2(n_6),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_126),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_15),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_128),
.B(n_4),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_4),
.B(n_7),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_7),
.B(n_8),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_133),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_7),
.B(n_8),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_20),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_134),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_130),
.C(n_9),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_138),
.A2(n_139),
.B(n_136),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_9),
.Y(n_141)
);


endmodule