module real_jpeg_11640_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_17;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_1),
.A2(n_19),
.B1(n_30),
.B2(n_31),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_6),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_4),
.B(n_6),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_21),
.C(n_29),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_3),
.B(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_4),
.B(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_22),
.C(n_28),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_18),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_17),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_15),
.B(n_16),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_25),
.B(n_36),
.C(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_34),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_39),
.B(n_40),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B(n_38),
.Y(n_32)
);


endmodule