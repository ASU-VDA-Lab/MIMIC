module fake_netlist_5_863_n_1919 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1919);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1919;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_315;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_119),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_106),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_60),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_162),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_62),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_17),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

BUFx8_ASAP7_75t_SL g196 ( 
.A(n_28),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_177),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_65),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_22),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_42),
.Y(n_202)
);

BUFx8_ASAP7_75t_SL g203 ( 
.A(n_183),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_20),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_187),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_161),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_75),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_37),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_111),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_97),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_38),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_118),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_11),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_18),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_102),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_11),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_40),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_146),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_42),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_73),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_3),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_91),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_145),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_57),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_184),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_110),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_43),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_27),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_46),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_182),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_67),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_133),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_93),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_25),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_41),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_36),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_116),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_59),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_31),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_98),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_5),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_82),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_41),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_96),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_112),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_44),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_109),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_51),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_9),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_44),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_2),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_30),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_103),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_142),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_79),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_174),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_66),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_7),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_159),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_165),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_4),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_81),
.Y(n_267)
);

BUFx2_ASAP7_75t_SL g268 ( 
.A(n_176),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_6),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_14),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_141),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_39),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_72),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_74),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_13),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_51),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_94),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_134),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_12),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_0),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_90),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_151),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_113),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_0),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_185),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_68),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_26),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_52),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_101),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_179),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_23),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_167),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_33),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_137),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_108),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_164),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_114),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_178),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_13),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_125),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_47),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_37),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_69),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_158),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_53),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_117),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_143),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_87),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_4),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_107),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_122),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_36),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_10),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_29),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_131),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_20),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_54),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_121),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_77),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_129),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_28),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_156),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_63),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_15),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_55),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_132),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_140),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_92),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_10),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_21),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_71),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_53),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_6),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_40),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_153),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_54),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_155),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_124),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_173),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_170),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_58),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_45),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_168),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_86),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_21),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_35),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_12),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_52),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_48),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_84),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_105),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_5),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_32),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_78),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_89),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_3),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_19),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_50),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_55),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_99),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_46),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_32),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_22),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_135),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_123),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_126),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_136),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_100),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_24),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_8),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_104),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_17),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_30),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_64),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_130),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_195),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_209),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_209),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_209),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_326),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_337),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_312),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_330),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_347),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_244),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_282),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_209),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_199),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_209),
.Y(n_389)
);

INVxp33_ASAP7_75t_SL g390 ( 
.A(n_194),
.Y(n_390)
);

INVxp33_ASAP7_75t_SL g391 ( 
.A(n_194),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_294),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_209),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_215),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_209),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_196),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_233),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_209),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_251),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_202),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_314),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_295),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_231),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_251),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_251),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_238),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_239),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_251),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_251),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_328),
.Y(n_410)
);

INVxp33_ASAP7_75t_SL g411 ( 
.A(n_215),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_251),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_251),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_251),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_240),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_248),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_243),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_351),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_248),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_203),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_204),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_248),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_358),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_200),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_213),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_375),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_213),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_266),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_224),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_245),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_224),
.Y(n_433)
);

INVxp33_ASAP7_75t_SL g434 ( 
.A(n_216),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_263),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_325),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_269),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_270),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_225),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_325),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_272),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_216),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_199),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_200),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_284),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_352),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_266),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_346),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_352),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_200),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_218),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_287),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g453 ( 
.A(n_346),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_285),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_266),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_266),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_266),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_219),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_219),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_302),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_302),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_288),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_336),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_291),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_336),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_293),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_221),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_254),
.Y(n_468)
);

BUFx8_ASAP7_75t_L g469 ( 
.A(n_388),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_454),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_376),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_397),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_397),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_385),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_455),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_386),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_381),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_447),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_447),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_430),
.Y(n_481)
);

AND2x2_ASAP7_75t_SL g482 ( 
.A(n_428),
.B(n_318),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_377),
.B(n_296),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_430),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_447),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_456),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_457),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_380),
.B(n_229),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_439),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_381),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_419),
.B(n_285),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_416),
.B(n_296),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_388),
.B(n_229),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_427),
.B(n_296),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_429),
.B(n_318),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_377),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_390),
.B(n_212),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_403),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_393),
.A2(n_368),
.B(n_366),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_431),
.B(n_227),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_383),
.A2(n_276),
.B1(n_253),
.B2(n_372),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_387),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_392),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_384),
.A2(n_359),
.B1(n_373),
.B2(n_372),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_387),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_381),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_378),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_389),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_402),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_389),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_406),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_416),
.B(n_366),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_381),
.Y(n_515)
);

BUFx8_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

OR2x6_ASAP7_75t_L g517 ( 
.A(n_396),
.B(n_268),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_422),
.B(n_368),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_395),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_395),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_436),
.B(n_227),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_440),
.B(n_188),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_398),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_442),
.Y(n_524)
);

OA21x2_ASAP7_75t_L g525 ( 
.A1(n_398),
.A2(n_211),
.B(n_201),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_379),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_381),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_399),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_408),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_446),
.B(n_227),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_399),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_404),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_412),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_382),
.A2(n_356),
.B1(n_373),
.B2(n_348),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_413),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_449),
.B(n_222),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_404),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_423),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_414),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_425),
.B(n_223),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_405),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_426),
.B(n_228),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_391),
.B(n_236),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_R g546 ( 
.A(n_407),
.B(n_189),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_405),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_458),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_491),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_482),
.A2(n_444),
.B1(n_450),
.B2(n_421),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_481),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_491),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_SL g553 ( 
.A(n_524),
.B(n_415),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_R g555 ( 
.A(n_472),
.B(n_415),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_497),
.Y(n_556)
);

INVx8_ASAP7_75t_L g557 ( 
.A(n_517),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_497),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_481),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_491),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_488),
.A2(n_411),
.B1(n_434),
.B2(n_394),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_492),
.B(n_458),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_499),
.B(n_401),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_470),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_482),
.B(n_417),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_533),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_498),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_498),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_533),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_544),
.A2(n_453),
.B1(n_256),
.B2(n_257),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_484),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_472),
.Y(n_572)
);

NAND3xp33_ASAP7_75t_SL g573 ( 
.A(n_536),
.B(n_432),
.C(n_417),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_484),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_L g575 ( 
.A1(n_536),
.A2(n_313),
.B1(n_345),
.B2(n_232),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_482),
.B(n_432),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_509),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_524),
.B(n_435),
.Y(n_578)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_477),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_487),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_494),
.B(n_435),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_504),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_504),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_534),
.B(n_437),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_469),
.B(n_437),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_507),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_509),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_469),
.B(n_438),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_502),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_507),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_502),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_510),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_510),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_533),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_491),
.Y(n_595)
);

BUFx8_ASAP7_75t_SL g596 ( 
.A(n_471),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_512),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_526),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_526),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_529),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g601 ( 
.A(n_506),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_529),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_477),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_544),
.B(n_242),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_535),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_L g606 ( 
.A1(n_517),
.A2(n_334),
.B1(n_342),
.B2(n_333),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_473),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_544),
.B(n_459),
.Y(n_608)
);

AO21x2_ASAP7_75t_L g609 ( 
.A1(n_501),
.A2(n_258),
.B(n_247),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_489),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_512),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_533),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_519),
.Y(n_613)
);

INVx8_ASAP7_75t_L g614 ( 
.A(n_517),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_544),
.A2(n_275),
.B1(n_279),
.B2(n_280),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_537),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_519),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_535),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_491),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_534),
.B(n_438),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_520),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_517),
.B(n_265),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_469),
.B(n_441),
.Y(n_623)
);

NOR2x1p5_ASAP7_75t_L g624 ( 
.A(n_540),
.B(n_348),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_508),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_508),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_520),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_475),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_508),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_537),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_521),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_475),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_478),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_478),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_508),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_523),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_523),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g638 ( 
.A(n_546),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_479),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_508),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_534),
.B(n_441),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_534),
.B(n_445),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_537),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_528),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_479),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_480),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_528),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_L g648 ( 
.A(n_500),
.B(n_445),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_532),
.B(n_539),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_521),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_469),
.B(n_452),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_513),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_532),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_539),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_540),
.B(n_459),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_543),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_531),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_543),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_537),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_525),
.A2(n_349),
.B1(n_299),
.B2(n_316),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_547),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_547),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_SL g663 ( 
.A1(n_522),
.A2(n_424),
.B1(n_452),
.B2(n_462),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_501),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_537),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_490),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_486),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_541),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_541),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_480),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_485),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_485),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_486),
.Y(n_673)
);

AO21x2_ASAP7_75t_L g674 ( 
.A1(n_483),
.A2(n_274),
.B(n_271),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_515),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_541),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_531),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_541),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_541),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_530),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_503),
.A2(n_356),
.B1(n_359),
.B2(n_363),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_515),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_514),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_514),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_515),
.Y(n_685)
);

INVx4_ASAP7_75t_SL g686 ( 
.A(n_515),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_490),
.Y(n_687)
);

INVx8_ASAP7_75t_L g688 ( 
.A(n_517),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_493),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_514),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_538),
.B(n_448),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_515),
.Y(n_692)
);

CKINVDCx6p67_ASAP7_75t_R g693 ( 
.A(n_474),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_477),
.B(n_462),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_527),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_527),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_493),
.B(n_464),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_493),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_514),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_564),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_624),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_689),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_689),
.B(n_525),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_698),
.B(n_525),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_638),
.B(n_464),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_589),
.B(n_516),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_698),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_638),
.A2(n_410),
.B1(n_418),
.B2(n_369),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_691),
.B(n_572),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_589),
.B(n_337),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_573),
.B(n_542),
.C(n_451),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_683),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_601),
.B(n_466),
.Y(n_713)
);

NAND2x1p5_ASAP7_75t_L g714 ( 
.A(n_683),
.B(n_684),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_567),
.B(n_568),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_684),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_567),
.B(n_525),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_556),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_584),
.B(n_466),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_568),
.B(n_493),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_655),
.B(n_467),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_582),
.B(n_518),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_591),
.B(n_337),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_596),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_565),
.A2(n_323),
.B1(n_262),
.B2(n_260),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_583),
.B(n_518),
.Y(n_726)
);

O2A1O1Ixp5_ASAP7_75t_L g727 ( 
.A1(n_664),
.A2(n_495),
.B(n_496),
.C(n_518),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_558),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_690),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_690),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_699),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_699),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_583),
.B(n_483),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_681),
.A2(n_400),
.B1(n_329),
.B2(n_353),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_624),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_586),
.B(n_277),
.Y(n_736)
);

AOI221xp5_ASAP7_75t_L g737 ( 
.A1(n_575),
.A2(n_363),
.B1(n_369),
.B2(n_361),
.C(n_357),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_559),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_586),
.B(n_278),
.Y(n_739)
);

O2A1O1Ixp5_ASAP7_75t_L g740 ( 
.A1(n_664),
.A2(n_310),
.B(n_283),
.C(n_354),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_680),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_590),
.B(n_286),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_620),
.B(n_189),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_641),
.B(n_190),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_L g745 ( 
.A(n_642),
.B(n_226),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_590),
.B(n_289),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_576),
.A2(n_255),
.B(n_362),
.C(n_370),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_559),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_592),
.B(n_290),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_571),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_691),
.B(n_190),
.Y(n_751)
);

NOR2x1p5_ASAP7_75t_L g752 ( 
.A(n_693),
.B(n_505),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_667),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_591),
.B(n_191),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_SL g755 ( 
.A(n_666),
.B(n_420),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_631),
.B(n_516),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_697),
.B(n_505),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_667),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_592),
.B(n_297),
.Y(n_759)
);

INVx5_ASAP7_75t_L g760 ( 
.A(n_549),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_631),
.B(n_511),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_608),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_650),
.B(n_516),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_593),
.B(n_298),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_593),
.B(n_304),
.Y(n_765)
);

BUFx8_ASAP7_75t_L g766 ( 
.A(n_650),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_597),
.B(n_306),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_597),
.B(n_611),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_608),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_611),
.Y(n_770)
);

NOR2x1p5_ASAP7_75t_L g771 ( 
.A(n_693),
.B(n_511),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_613),
.B(n_311),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_657),
.B(n_337),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_613),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_617),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_571),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_657),
.B(n_337),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_617),
.B(n_322),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_621),
.B(n_339),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_621),
.B(n_350),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_627),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_571),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_627),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_549),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_636),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_687),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_677),
.B(n_360),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_644),
.B(n_360),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_636),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_581),
.A2(n_267),
.B1(n_230),
.B2(n_234),
.Y(n_790)
);

O2A1O1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_649),
.A2(n_562),
.B(n_647),
.C(n_637),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_562),
.A2(n_468),
.B(n_365),
.C(n_463),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_563),
.B(n_191),
.Y(n_793)
);

OR2x6_ASAP7_75t_L g794 ( 
.A(n_557),
.B(n_468),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_644),
.B(n_360),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_637),
.Y(n_796)
);

AND2x2_ASAP7_75t_SL g797 ( 
.A(n_660),
.B(n_681),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_647),
.B(n_654),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_578),
.B(n_192),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_561),
.B(n_516),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_574),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_654),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_574),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_658),
.B(n_527),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_658),
.B(n_527),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_550),
.B(n_192),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_574),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_694),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_606),
.B(n_193),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_661),
.A2(n_548),
.B(n_341),
.C(n_340),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_607),
.B(n_476),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_661),
.B(n_527),
.Y(n_812)
);

NOR2xp67_ASAP7_75t_L g813 ( 
.A(n_585),
.B(n_548),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_662),
.B(n_235),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_662),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_604),
.B(n_237),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_551),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_673),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_549),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_673),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_663),
.B(n_193),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_SL g822 ( 
.A(n_610),
.B(n_273),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_604),
.B(n_241),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_570),
.B(n_305),
.C(n_301),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_604),
.B(n_246),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_549),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_604),
.B(n_249),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_644),
.B(n_360),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_653),
.B(n_656),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_653),
.Y(n_830)
);

NOR3xp33_ASAP7_75t_L g831 ( 
.A(n_553),
.B(n_648),
.C(n_623),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_653),
.B(n_250),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_656),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_664),
.A2(n_309),
.B1(n_324),
.B2(n_321),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_555),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_622),
.A2(n_197),
.B1(n_198),
.B2(n_205),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_610),
.B(n_197),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_656),
.B(n_252),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_610),
.B(n_652),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_610),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_639),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_645),
.Y(n_842)
);

INVx8_ASAP7_75t_L g843 ( 
.A(n_557),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_549),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_579),
.B(n_259),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_665),
.B(n_668),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_588),
.B(n_261),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_603),
.B(n_264),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_652),
.B(n_465),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_628),
.B(n_292),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_SL g851 ( 
.A(n_651),
.B(n_317),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_632),
.B(n_300),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_645),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_549),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_557),
.B(n_460),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_577),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_652),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_646),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_646),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_712),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_716),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_700),
.B(n_632),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_729),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_709),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_784),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_700),
.B(n_633),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_715),
.B(n_633),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_762),
.B(n_769),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_786),
.Y(n_869)
);

AND2x4_ASAP7_75t_SL g870 ( 
.A(n_811),
.B(n_652),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_741),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_761),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_730),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_797),
.A2(n_614),
.B1(n_557),
.B2(n_688),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_768),
.B(n_634),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_849),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_721),
.Y(n_877)
);

NOR2x1_ASAP7_75t_L g878 ( 
.A(n_757),
.B(n_622),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_731),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_798),
.B(n_770),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_797),
.A2(n_587),
.B1(n_557),
.B2(n_614),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_732),
.Y(n_882)
);

O2A1O1Ixp5_ASAP7_75t_L g883 ( 
.A1(n_740),
.A2(n_727),
.B(n_723),
.C(n_710),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_841),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_721),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_751),
.B(n_622),
.Y(n_886)
);

AND2x6_ASAP7_75t_L g887 ( 
.A(n_717),
.B(n_665),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_701),
.B(n_622),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_774),
.B(n_634),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_842),
.Y(n_890)
);

NOR2x1p5_ASAP7_75t_L g891 ( 
.A(n_724),
.B(n_332),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_775),
.B(n_587),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_781),
.B(n_577),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_714),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_705),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_853),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_830),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_783),
.B(n_577),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_834),
.A2(n_688),
.B1(n_614),
.B2(n_672),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_858),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_766),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_859),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_713),
.A2(n_622),
.B1(n_614),
.B2(n_688),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_835),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_818),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_784),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_833),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_766),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_843),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_714),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_785),
.B(n_598),
.Y(n_911)
);

NOR2x1_ASAP7_75t_R g912 ( 
.A(n_800),
.B(n_198),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_789),
.B(n_598),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_843),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_843),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_820),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_735),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_719),
.B(n_614),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_796),
.B(n_598),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_713),
.A2(n_688),
.B1(n_594),
.B2(n_569),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_817),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_802),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_719),
.A2(n_688),
.B1(n_594),
.B2(n_569),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_815),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_813),
.B(n_670),
.Y(n_925)
);

NAND3xp33_ASAP7_75t_SL g926 ( 
.A(n_831),
.B(n_615),
.C(n_206),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_835),
.Y(n_927)
);

AND2x6_ASAP7_75t_L g928 ( 
.A(n_703),
.B(n_665),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_727),
.A2(n_676),
.B(n_668),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_708),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_834),
.A2(n_711),
.B1(n_758),
.B2(n_753),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_808),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_711),
.A2(n_744),
.B1(n_743),
.B2(n_707),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_702),
.B(n_599),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_743),
.B(n_668),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_718),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_R g937 ( 
.A(n_755),
.B(n_205),
.Y(n_937)
);

AND2x6_ASAP7_75t_SL g938 ( 
.A(n_799),
.B(n_460),
.Y(n_938)
);

INVx5_ASAP7_75t_L g939 ( 
.A(n_784),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_784),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_720),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_728),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_791),
.B(n_599),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_829),
.B(n_599),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_857),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_831),
.A2(n_594),
.B1(n_630),
.B2(n_643),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_819),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_855),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_816),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_722),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_726),
.B(n_600),
.Y(n_951)
);

BUFx10_ASAP7_75t_L g952 ( 
.A(n_793),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_804),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_823),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_704),
.B(n_600),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_738),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_805),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_737),
.A2(n_670),
.B1(n_671),
.B2(n_672),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_793),
.B(n_630),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_708),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_794),
.B(n_671),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_822),
.B(n_676),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_799),
.B(n_678),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_809),
.A2(n_806),
.B1(n_736),
.B2(n_739),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_742),
.B(n_600),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_855),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_746),
.B(n_602),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_832),
.A2(n_745),
.B1(n_827),
.B2(n_825),
.Y(n_968)
);

OR2x2_ASAP7_75t_SL g969 ( 
.A(n_824),
.B(n_461),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_812),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_749),
.B(n_602),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_856),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_840),
.B(n_678),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_759),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_840),
.B(n_678),
.Y(n_975)
);

AND3x1_ASAP7_75t_L g976 ( 
.A(n_754),
.B(n_725),
.C(n_747),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_764),
.B(n_602),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_748),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_754),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_L g980 ( 
.A(n_819),
.B(n_679),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_837),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_819),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_733),
.A2(n_612),
.B(n_554),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_750),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_790),
.B(n_679),
.Y(n_985)
);

NAND2x1p5_ASAP7_75t_L g986 ( 
.A(n_819),
.B(n_630),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_776),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_782),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_801),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_794),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_821),
.B(n_643),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_794),
.A2(n_679),
.B1(n_643),
.B2(n_669),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_765),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_846),
.A2(n_612),
.B(n_554),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_767),
.B(n_605),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_803),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_772),
.B(n_778),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_855),
.B(n_706),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_779),
.B(n_605),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_807),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_847),
.B(n_206),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_756),
.B(n_659),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_839),
.B(n_674),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_780),
.B(n_605),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_SL g1005 ( 
.A1(n_836),
.A2(n_208),
.B1(n_210),
.B2(n_214),
.Y(n_1005)
);

INVx5_ASAP7_75t_L g1006 ( 
.A(n_826),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_710),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_826),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_846),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_723),
.B(n_618),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_851),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_773),
.B(n_618),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_734),
.B(n_763),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_734),
.B(n_659),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_845),
.B(n_669),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_826),
.B(n_554),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_826),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_740),
.A2(n_618),
.B(n_682),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_844),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_850),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_777),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_852),
.B(n_609),
.Y(n_1022)
);

INVxp33_ASAP7_75t_L g1023 ( 
.A(n_752),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_771),
.B(n_609),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_848),
.B(n_207),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_777),
.B(n_609),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_787),
.B(n_580),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_844),
.Y(n_1028)
);

BUFx8_ASAP7_75t_L g1029 ( 
.A(n_844),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_787),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_788),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_788),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_844),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_795),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_854),
.B(n_692),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_838),
.B(n_554),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_795),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_1013),
.A2(n_273),
.B1(n_828),
.B2(n_814),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_860),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_865),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_979),
.B(n_810),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_929),
.A2(n_828),
.B(n_692),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_871),
.Y(n_1043)
);

AOI222xp33_ASAP7_75t_L g1044 ( 
.A1(n_930),
.A2(n_273),
.B1(n_465),
.B2(n_461),
.C1(n_463),
.C2(n_208),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_904),
.B(n_927),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_997),
.A2(n_760),
.B(n_612),
.Y(n_1046)
);

INVx5_ASAP7_75t_L g1047 ( 
.A(n_865),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_879),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_876),
.B(n_854),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_997),
.A2(n_760),
.B(n_612),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_869),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_862),
.B(n_792),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_933),
.A2(n_682),
.B(n_692),
.C(n_696),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_865),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_864),
.Y(n_1055)
);

NOR3xp33_ASAP7_75t_L g1056 ( 
.A(n_886),
.B(n_374),
.C(n_371),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_861),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_994),
.A2(n_695),
.B(n_696),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_952),
.B(n_854),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_863),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_L g1061 ( 
.A(n_894),
.B(n_760),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_895),
.B(n_207),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_932),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_993),
.B(n_210),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_880),
.A2(n_760),
.B(n_616),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_917),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_993),
.B(n_214),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_883),
.A2(n_696),
.B(n_695),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_952),
.B(n_217),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_880),
.A2(n_566),
.B(n_616),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_881),
.A2(n_566),
.B1(n_616),
.B2(n_217),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_926),
.A2(n_367),
.B1(n_281),
.B2(n_343),
.Y(n_1072)
);

CKINVDCx6p67_ASAP7_75t_R g1073 ( 
.A(n_1024),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_862),
.B(n_552),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_873),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_903),
.A2(n_566),
.B1(n_616),
.B2(n_220),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_955),
.A2(n_566),
.B(n_560),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_949),
.A2(n_954),
.B1(n_976),
.B2(n_991),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_882),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_922),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_866),
.B(n_959),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1029),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_866),
.B(n_552),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_872),
.B(n_220),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_867),
.A2(n_675),
.B(n_552),
.C(n_595),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_SL g1086 ( 
.A1(n_1007),
.A2(n_552),
.B(n_675),
.C(n_640),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_924),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1007),
.A2(n_364),
.B1(n_281),
.B2(n_367),
.Y(n_1088)
);

OAI21xp33_ASAP7_75t_L g1089 ( 
.A1(n_931),
.A2(n_344),
.B(n_374),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_974),
.B(n_343),
.Y(n_1090)
);

INVx4_ASAP7_75t_L g1091 ( 
.A(n_909),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_906),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_950),
.B(n_619),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_960),
.B(n_344),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_955),
.A2(n_560),
.B(n_685),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_951),
.A2(n_560),
.B(n_685),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_981),
.B(n_355),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_885),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_877),
.B(n_355),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_941),
.B(n_625),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_951),
.A2(n_560),
.B(n_685),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_892),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1020),
.B(n_364),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_892),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_899),
.A2(n_625),
.B1(n_626),
.B2(n_675),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_867),
.A2(n_560),
.B(n_685),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_1029),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_875),
.A2(n_560),
.B(n_685),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_938),
.B(n_1014),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_1015),
.A2(n_1036),
.B(n_964),
.C(n_968),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_906),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_894),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_889),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_875),
.B(n_625),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_953),
.B(n_626),
.Y(n_1115)
);

BUFx4f_ASAP7_75t_L g1116 ( 
.A(n_998),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_936),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_957),
.B(n_626),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_906),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_874),
.A2(n_626),
.B1(n_629),
.B2(n_640),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_969),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_970),
.B(n_868),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_870),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_965),
.A2(n_685),
.B(n_635),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_SL g1125 ( 
.A(n_937),
.B(n_303),
.C(n_307),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_SL g1126 ( 
.A1(n_1005),
.A2(n_308),
.B1(n_315),
.B2(n_319),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_889),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_R g1128 ( 
.A(n_926),
.B(n_320),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_868),
.B(n_338),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_893),
.Y(n_1130)
);

CKINVDCx8_ASAP7_75t_R g1131 ( 
.A(n_1024),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_901),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_888),
.B(n_629),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_942),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_940),
.Y(n_1135)
);

INVx4_ASAP7_75t_L g1136 ( 
.A(n_914),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_943),
.A2(n_629),
.B(n_2),
.C(n_7),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_L g1138 ( 
.A(n_878),
.B(n_327),
.C(n_331),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_SL g1139 ( 
.A(n_908),
.B(n_335),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_998),
.B(n_635),
.Y(n_1140)
);

NOR2x1_ASAP7_75t_SL g1141 ( 
.A(n_939),
.B(n_635),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_940),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_884),
.B(n_890),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1021),
.A2(n_635),
.B1(n_76),
.B2(n_186),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_990),
.B(n_1),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_965),
.A2(n_971),
.B(n_967),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_943),
.A2(n_1),
.B(n_8),
.C(n_9),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_914),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_896),
.B(n_635),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_940),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_888),
.B(n_14),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_948),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_945),
.B(n_15),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1025),
.B(n_635),
.C(n_18),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1011),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1030),
.A2(n_16),
.B(n_19),
.C(n_23),
.Y(n_1156)
);

AOI222xp33_ASAP7_75t_L g1157 ( 
.A1(n_912),
.A2(n_1001),
.B1(n_1023),
.B2(n_891),
.C1(n_948),
.C2(n_966),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_966),
.B(n_16),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_967),
.A2(n_686),
.B(n_85),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_L g1160 ( 
.A(n_962),
.B(n_24),
.C(n_25),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_900),
.B(n_686),
.Y(n_1161)
);

AOI21x1_ASAP7_75t_L g1162 ( 
.A1(n_935),
.A2(n_686),
.B(n_95),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_902),
.B(n_686),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_910),
.B(n_88),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_905),
.B(n_26),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_916),
.B(n_27),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_958),
.B(n_29),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_982),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_939),
.B(n_120),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_982),
.Y(n_1170)
);

NOR3xp33_ASAP7_75t_SL g1171 ( 
.A(n_973),
.B(n_33),
.C(n_34),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_971),
.A2(n_127),
.B(n_180),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_893),
.B(n_898),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1022),
.A2(n_35),
.B(n_38),
.C(n_39),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_911),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_961),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_956),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_911),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_SL g1179 ( 
.A1(n_1018),
.A2(n_138),
.B(n_172),
.C(n_171),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_987),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1009),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_913),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1003),
.A2(n_139),
.B1(n_169),
.B2(n_61),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_913),
.B(n_49),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_915),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1102),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1120),
.A2(n_992),
.A3(n_983),
.B(n_995),
.Y(n_1187)
);

INVx8_ASAP7_75t_L g1188 ( 
.A(n_1047),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1109),
.A2(n_963),
.B1(n_1002),
.B2(n_918),
.C(n_919),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1081),
.B(n_1002),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1104),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1113),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1078),
.B(n_925),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1146),
.A2(n_1110),
.B(n_1173),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1091),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1095),
.A2(n_1042),
.B(n_1124),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1061),
.A2(n_939),
.B(n_1006),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1127),
.A2(n_920),
.B1(n_923),
.B2(n_946),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1130),
.B(n_999),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1043),
.Y(n_1200)
);

O2A1O1Ixp5_ASAP7_75t_L g1201 ( 
.A1(n_1159),
.A2(n_985),
.B(n_975),
.C(n_1026),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1051),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1055),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1066),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1175),
.B(n_977),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1073),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1045),
.B(n_1006),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1057),
.Y(n_1208)
);

AND2x6_ASAP7_75t_L g1209 ( 
.A(n_1178),
.B(n_1026),
.Y(n_1209)
);

OR2x6_ASAP7_75t_L g1210 ( 
.A(n_1082),
.B(n_1107),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1070),
.A2(n_1004),
.B(n_977),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1053),
.A2(n_983),
.A3(n_995),
.B(n_999),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1055),
.Y(n_1213)
);

AOI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_1044),
.A2(n_1037),
.B(n_1034),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1182),
.B(n_1004),
.Y(n_1215)
);

BUFx10_ASAP7_75t_L g1216 ( 
.A(n_1103),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1060),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1122),
.B(n_944),
.Y(n_1218)
);

NAND3x1_ASAP7_75t_L g1219 ( 
.A(n_1158),
.B(n_947),
.C(n_984),
.Y(n_1219)
);

NAND2xp33_ASAP7_75t_L g1220 ( 
.A(n_1167),
.B(n_1008),
.Y(n_1220)
);

INVxp67_ASAP7_75t_SL g1221 ( 
.A(n_1112),
.Y(n_1221)
);

AOI221x1_ASAP7_75t_L g1222 ( 
.A1(n_1160),
.A2(n_994),
.B1(n_919),
.B2(n_944),
.C(n_934),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1077),
.A2(n_1050),
.B(n_1046),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1041),
.A2(n_1052),
.B(n_1038),
.C(n_1056),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1038),
.A2(n_1032),
.B(n_1031),
.C(n_934),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1077),
.A2(n_1016),
.B(n_980),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1067),
.B(n_921),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1046),
.A2(n_1016),
.B(n_1017),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1075),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1124),
.A2(n_1035),
.B(n_1012),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1056),
.A2(n_972),
.B(n_978),
.C(n_988),
.Y(n_1231)
);

OA22x2_ASAP7_75t_L g1232 ( 
.A1(n_1121),
.A2(n_1033),
.B1(n_1028),
.B2(n_1019),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1154),
.A2(n_989),
.B(n_907),
.C(n_897),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1096),
.A2(n_1035),
.B(n_1010),
.Y(n_1234)
);

AOI21xp33_ASAP7_75t_L g1235 ( 
.A1(n_1062),
.A2(n_1027),
.B(n_1000),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1064),
.B(n_996),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1184),
.A2(n_887),
.B(n_928),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1101),
.A2(n_986),
.B(n_887),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1098),
.B(n_1008),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1080),
.Y(n_1240)
);

AO21x2_ASAP7_75t_L g1241 ( 
.A1(n_1085),
.A2(n_887),
.B(n_928),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1106),
.A2(n_887),
.B(n_928),
.Y(n_1242)
);

OR2x6_ASAP7_75t_L g1243 ( 
.A(n_1155),
.B(n_1008),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1091),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1063),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1064),
.B(n_928),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_SL g1247 ( 
.A1(n_1172),
.A2(n_1017),
.B(n_887),
.Y(n_1247)
);

OAI21xp33_ASAP7_75t_L g1248 ( 
.A1(n_1072),
.A2(n_928),
.B(n_56),
.Y(n_1248)
);

NOR4xp25_ASAP7_75t_L g1249 ( 
.A(n_1147),
.B(n_56),
.C(n_70),
.D(n_80),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1040),
.Y(n_1250)
);

NOR2xp67_ASAP7_75t_SL g1251 ( 
.A(n_1131),
.B(n_83),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1040),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1047),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1097),
.B(n_128),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1087),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1116),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_1256)
);

AND3x4_ASAP7_75t_L g1257 ( 
.A(n_1132),
.B(n_152),
.C(n_154),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1065),
.A2(n_1141),
.B(n_1106),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1143),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1123),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1116),
.A2(n_1049),
.B1(n_1140),
.B2(n_1079),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1039),
.Y(n_1262)
);

AO22x2_ASAP7_75t_L g1263 ( 
.A1(n_1160),
.A2(n_1144),
.B1(n_1165),
.B2(n_1166),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1108),
.A2(n_1114),
.B(n_1085),
.Y(n_1264)
);

AOI21xp33_ASAP7_75t_L g1265 ( 
.A1(n_1089),
.A2(n_1072),
.B(n_1090),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_SL g1266 ( 
.A1(n_1179),
.A2(n_1164),
.B(n_1174),
.C(n_1169),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1112),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1162),
.A2(n_1105),
.B(n_1159),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1074),
.A2(n_1083),
.B(n_1076),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1048),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1115),
.A2(n_1118),
.B(n_1093),
.Y(n_1271)
);

AO31x2_ASAP7_75t_L g1272 ( 
.A1(n_1071),
.A2(n_1172),
.A3(n_1156),
.B(n_1100),
.Y(n_1272)
);

BUFx8_ASAP7_75t_L g1273 ( 
.A(n_1152),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1151),
.B(n_1117),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1069),
.B(n_1084),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1183),
.A2(n_1138),
.B(n_1137),
.C(n_1147),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1157),
.B(n_1128),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1134),
.B(n_1180),
.Y(n_1278)
);

AOI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1088),
.A2(n_1129),
.B(n_1099),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1177),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1133),
.B(n_1185),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1047),
.A2(n_1133),
.B1(n_1181),
.B2(n_1148),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1040),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1142),
.B(n_1153),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1047),
.A2(n_1181),
.B1(n_1148),
.B2(n_1136),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1149),
.A2(n_1163),
.A3(n_1161),
.B(n_1086),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1137),
.A2(n_1171),
.A3(n_1185),
.B(n_1136),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1139),
.B(n_1126),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1054),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1145),
.B(n_1171),
.Y(n_1290)
);

CKINVDCx16_ASAP7_75t_R g1291 ( 
.A(n_1125),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1059),
.B(n_1135),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1054),
.B(n_1092),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1125),
.B(n_1150),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1150),
.A2(n_1054),
.B(n_1092),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_SL g1296 ( 
.A1(n_1092),
.A2(n_1111),
.B(n_1119),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1111),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1111),
.A2(n_1119),
.B(n_1168),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1119),
.A2(n_1168),
.B(n_1170),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1168),
.B(n_1170),
.Y(n_1300)
);

NAND3xp33_ASAP7_75t_SL g1301 ( 
.A(n_1170),
.B(n_490),
.C(n_564),
.Y(n_1301)
);

CKINVDCx16_ASAP7_75t_R g1302 ( 
.A(n_1051),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1146),
.A2(n_1110),
.B(n_1173),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1078),
.B(n_638),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1091),
.B(n_909),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1081),
.B(n_700),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1081),
.B(n_700),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1078),
.B(n_638),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1176),
.B(n_1133),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1043),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1057),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1102),
.Y(n_1312)
);

INVx5_ASAP7_75t_L g1313 ( 
.A(n_1040),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1122),
.B(n_709),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_SL g1315 ( 
.A1(n_1110),
.A2(n_1179),
.B(n_1167),
.C(n_1164),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1058),
.A2(n_1095),
.B(n_1068),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1081),
.B(n_700),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1078),
.B(n_638),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1081),
.A2(n_700),
.B1(n_1078),
.B2(n_979),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1081),
.B(n_700),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1058),
.A2(n_1095),
.B(n_1068),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1094),
.B(n_705),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1040),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1081),
.B(n_700),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1043),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1081),
.B(n_700),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1058),
.A2(n_1095),
.B(n_1068),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1094),
.B(n_705),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1102),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1146),
.A2(n_1110),
.B(n_1173),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_SL g1331 ( 
.A(n_1051),
.B(n_786),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1306),
.A2(n_1320),
.B1(n_1307),
.B2(n_1324),
.Y(n_1332)
);

NOR2x1_ASAP7_75t_SL g1333 ( 
.A(n_1193),
.B(n_1186),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1240),
.Y(n_1334)
);

OR2x6_ASAP7_75t_L g1335 ( 
.A(n_1188),
.B(n_1219),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1267),
.Y(n_1336)
);

NOR2xp67_ASAP7_75t_L g1337 ( 
.A(n_1310),
.B(n_1325),
.Y(n_1337)
);

INVx4_ASAP7_75t_L g1338 ( 
.A(n_1188),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1322),
.B(n_1328),
.Y(n_1339)
);

AOI22x1_ASAP7_75t_SL g1340 ( 
.A1(n_1206),
.A2(n_1202),
.B1(n_1260),
.B2(n_1245),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1303),
.A2(n_1330),
.B(n_1211),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1313),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1319),
.B(n_1189),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1311),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1302),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1226),
.A2(n_1321),
.B(n_1316),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1317),
.A2(n_1326),
.B1(n_1248),
.B2(n_1259),
.Y(n_1347)
);

BUFx2_ASAP7_75t_SL g1348 ( 
.A(n_1200),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1208),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1327),
.A2(n_1230),
.B(n_1234),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1264),
.A2(n_1268),
.B(n_1237),
.Y(n_1351)
);

INVxp67_ASAP7_75t_L g1352 ( 
.A(n_1203),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1273),
.Y(n_1353)
);

CKINVDCx6p67_ASAP7_75t_R g1354 ( 
.A(n_1243),
.Y(n_1354)
);

OR2x6_ASAP7_75t_L g1355 ( 
.A(n_1285),
.B(n_1232),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1288),
.A2(n_1254),
.B1(n_1291),
.B2(n_1290),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1271),
.A2(n_1269),
.B(n_1201),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1213),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1277),
.A2(n_1265),
.B1(n_1263),
.B2(n_1318),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1221),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1262),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1309),
.B(n_1281),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1217),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1190),
.A2(n_1236),
.B1(n_1314),
.B2(n_1218),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1273),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1282),
.B(n_1197),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1309),
.B(n_1281),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1284),
.B(n_1227),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1229),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1274),
.B(n_1304),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1216),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1308),
.A2(n_1205),
.B1(n_1215),
.B2(n_1199),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1261),
.B(n_1294),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1263),
.A2(n_1214),
.B1(n_1279),
.B2(n_1257),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1255),
.Y(n_1375)
);

NAND2x1p5_ASAP7_75t_L g1376 ( 
.A(n_1253),
.B(n_1313),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1198),
.A2(n_1246),
.B(n_1222),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1224),
.B(n_1276),
.C(n_1275),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1270),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1280),
.Y(n_1380)
);

BUFx4f_ASAP7_75t_SL g1381 ( 
.A(n_1250),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1191),
.B(n_1192),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1192),
.Y(n_1383)
);

OAI211xp5_ASAP7_75t_L g1384 ( 
.A1(n_1249),
.A2(n_1301),
.B(n_1266),
.C(n_1315),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1313),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1225),
.A2(n_1231),
.B(n_1220),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1204),
.Y(n_1387)
);

NAND2xp33_ASAP7_75t_L g1388 ( 
.A(n_1209),
.B(n_1305),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1233),
.A2(n_1235),
.B(n_1329),
.Y(n_1389)
);

BUFx4f_ASAP7_75t_L g1390 ( 
.A(n_1210),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1312),
.Y(n_1391)
);

AOI21xp33_ASAP7_75t_L g1392 ( 
.A1(n_1241),
.A2(n_1207),
.B(n_1256),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1243),
.B(n_1239),
.Y(n_1393)
);

BUFx10_ASAP7_75t_L g1394 ( 
.A(n_1210),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1331),
.B(n_1278),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1250),
.Y(n_1396)
);

NAND2x1p5_ASAP7_75t_L g1397 ( 
.A(n_1253),
.B(n_1195),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1300),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1251),
.A2(n_1292),
.B(n_1295),
.C(n_1299),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1298),
.A2(n_1244),
.B(n_1195),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1289),
.Y(n_1401)
);

INVx4_ASAP7_75t_SL g1402 ( 
.A(n_1209),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1244),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1209),
.B(n_1212),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1241),
.A2(n_1296),
.B(n_1293),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1289),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1297),
.A2(n_1272),
.B(n_1323),
.C(n_1250),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1323),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1272),
.A2(n_1187),
.B(n_1286),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1252),
.B(n_1283),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1252),
.A2(n_1283),
.B1(n_1323),
.B2(n_1287),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1287),
.B(n_1187),
.Y(n_1412)
);

INVx3_ASAP7_75t_SL g1413 ( 
.A(n_1252),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1283),
.B(n_1287),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1187),
.A2(n_1242),
.B(n_1238),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1313),
.Y(n_1416)
);

BUFx10_ASAP7_75t_L g1417 ( 
.A(n_1245),
.Y(n_1417)
);

BUFx2_ASAP7_75t_R g1418 ( 
.A(n_1202),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1194),
.A2(n_1110),
.B(n_1303),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1224),
.A2(n_1303),
.B(n_1194),
.Y(n_1420)
);

AO31x2_ASAP7_75t_L g1421 ( 
.A1(n_1258),
.A2(n_1223),
.A3(n_1303),
.B(n_1194),
.Y(n_1421)
);

AO31x2_ASAP7_75t_L g1422 ( 
.A1(n_1223),
.A2(n_1264),
.A3(n_1303),
.B(n_1194),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1200),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1240),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1224),
.A2(n_1303),
.B(n_1194),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1239),
.Y(n_1426)
);

CKINVDCx16_ASAP7_75t_R g1427 ( 
.A(n_1331),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1240),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1200),
.Y(n_1429)
);

BUFx2_ASAP7_75t_R g1430 ( 
.A(n_1202),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1200),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1240),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1306),
.A2(n_700),
.B1(n_1181),
.B2(n_1109),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1277),
.A2(n_700),
.B1(n_960),
.B2(n_930),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1240),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1240),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1200),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1277),
.B(n_700),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1242),
.A2(n_1238),
.B(n_1196),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1224),
.A2(n_1303),
.B(n_1194),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1240),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1319),
.B(n_1078),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1242),
.A2(n_1238),
.B(n_1196),
.Y(n_1443)
);

BUFx2_ASAP7_75t_SL g1444 ( 
.A(n_1260),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1240),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1277),
.A2(n_1013),
.B1(n_1248),
.B2(n_1109),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1194),
.A2(n_1110),
.B(n_1303),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1309),
.B(n_1281),
.Y(n_1448)
);

INVx8_ASAP7_75t_L g1449 ( 
.A(n_1188),
.Y(n_1449)
);

AOI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1226),
.A2(n_918),
.B(n_1228),
.Y(n_1450)
);

BUFx12f_ASAP7_75t_L g1451 ( 
.A(n_1245),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1224),
.A2(n_1303),
.B(n_1194),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1240),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1224),
.A2(n_1303),
.B(n_1194),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_SL g1455 ( 
.A1(n_1247),
.A2(n_1137),
.B(n_1197),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1224),
.A2(n_1303),
.B(n_1194),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1313),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1383),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1347),
.A2(n_1333),
.B(n_1438),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1402),
.B(n_1393),
.Y(n_1460)
);

AOI21x1_ASAP7_75t_SL g1461 ( 
.A1(n_1412),
.A2(n_1414),
.B(n_1404),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1426),
.B(n_1370),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1368),
.B(n_1339),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1342),
.Y(n_1464)
);

NOR2xp67_ASAP7_75t_L g1465 ( 
.A(n_1378),
.B(n_1387),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1420),
.A2(n_1440),
.B(n_1425),
.Y(n_1466)
);

AOI21x1_ASAP7_75t_SL g1467 ( 
.A1(n_1412),
.A2(n_1414),
.B(n_1404),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1426),
.B(n_1336),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1360),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1336),
.B(n_1360),
.Y(n_1470)
);

O2A1O1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1433),
.A2(n_1438),
.B(n_1434),
.C(n_1343),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1446),
.A2(n_1434),
.B1(n_1374),
.B2(n_1359),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1341),
.A2(n_1425),
.B(n_1420),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1341),
.A2(n_1452),
.B(n_1440),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1343),
.A2(n_1442),
.B(n_1433),
.C(n_1372),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1452),
.A2(n_1456),
.B(n_1454),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1347),
.A2(n_1332),
.B(n_1399),
.Y(n_1477)
);

CKINVDCx6p67_ASAP7_75t_R g1478 ( 
.A(n_1345),
.Y(n_1478)
);

CKINVDCx16_ASAP7_75t_R g1479 ( 
.A(n_1427),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1332),
.A2(n_1399),
.B(n_1395),
.Y(n_1480)
);

INVx5_ASAP7_75t_L g1481 ( 
.A(n_1335),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1442),
.A2(n_1372),
.B(n_1446),
.C(n_1384),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1398),
.B(n_1356),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1373),
.B(n_1391),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1352),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1356),
.B(n_1359),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1352),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1364),
.B(n_1382),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1371),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1419),
.A2(n_1447),
.B(n_1409),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1395),
.A2(n_1386),
.B(n_1416),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1406),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1382),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1342),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1451),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1353),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1361),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1409),
.A2(n_1386),
.B(n_1357),
.Y(n_1498)
);

OAI22x1_ASAP7_75t_L g1499 ( 
.A1(n_1349),
.A2(n_1363),
.B1(n_1369),
.B2(n_1375),
.Y(n_1499)
);

O2A1O1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1364),
.A2(n_1374),
.B(n_1392),
.C(n_1455),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1390),
.A2(n_1355),
.B1(n_1334),
.B2(n_1428),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1373),
.B(n_1355),
.Y(n_1502)
);

O2A1O1Ixp5_ASAP7_75t_L g1503 ( 
.A1(n_1392),
.A2(n_1405),
.B(n_1407),
.C(n_1450),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1355),
.B(n_1389),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1362),
.B(n_1367),
.Y(n_1505)
);

CKINVDCx6p67_ASAP7_75t_R g1506 ( 
.A(n_1444),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1415),
.A2(n_1377),
.B(n_1350),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1389),
.B(n_1379),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1344),
.A2(n_1453),
.B1(n_1432),
.B2(n_1435),
.C(n_1445),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1424),
.B(n_1436),
.Y(n_1510)
);

AOI221x1_ASAP7_75t_SL g1511 ( 
.A1(n_1337),
.A2(n_1441),
.B1(n_1401),
.B2(n_1380),
.C(n_1448),
.Y(n_1511)
);

AND2x2_ASAP7_75t_SL g1512 ( 
.A(n_1388),
.B(n_1390),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1423),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1358),
.B(n_1413),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1407),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1413),
.B(n_1410),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1418),
.A2(n_1430),
.B1(n_1354),
.B2(n_1366),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1348),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1411),
.B(n_1405),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1410),
.B(n_1396),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1340),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_R g1522 ( 
.A(n_1381),
.B(n_1449),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1351),
.A2(n_1366),
.B(n_1346),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1385),
.A2(n_1457),
.B(n_1416),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1366),
.B(n_1422),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1411),
.B(n_1422),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1403),
.B(n_1408),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1394),
.B(n_1397),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1394),
.B(n_1397),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1385),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1422),
.B(n_1421),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1418),
.A2(n_1335),
.B1(n_1365),
.B2(n_1381),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1335),
.B(n_1417),
.Y(n_1533)
);

O2A1O1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1437),
.A2(n_1429),
.B(n_1431),
.C(n_1376),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1385),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1439),
.A2(n_1443),
.B(n_1400),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1417),
.B(n_1457),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1402),
.A2(n_1416),
.B(n_1457),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1338),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1338),
.B(n_1449),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1364),
.B(n_1332),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1341),
.A2(n_1110),
.B(n_1420),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1446),
.A2(n_1181),
.B1(n_1438),
.B2(n_700),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1364),
.B(n_1332),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1423),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1420),
.A2(n_1440),
.B(n_1425),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1420),
.A2(n_1440),
.B(n_1425),
.Y(n_1547)
);

O2A1O1Ixp5_ASAP7_75t_L g1548 ( 
.A1(n_1384),
.A2(n_1343),
.B(n_1277),
.C(n_1386),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1368),
.B(n_1339),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1393),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1446),
.A2(n_1181),
.B1(n_1438),
.B2(n_700),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1345),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1360),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1383),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1364),
.B(n_1332),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1420),
.A2(n_1440),
.B(n_1425),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1368),
.B(n_1339),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1446),
.A2(n_1181),
.B1(n_1438),
.B2(n_700),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1368),
.B(n_1339),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1462),
.B(n_1468),
.Y(n_1560)
);

NAND2x1_ASAP7_75t_L g1561 ( 
.A(n_1477),
.B(n_1480),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1496),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1525),
.B(n_1504),
.Y(n_1563)
);

INVxp67_ASAP7_75t_SL g1564 ( 
.A(n_1469),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1508),
.Y(n_1565)
);

AOI21xp33_ASAP7_75t_L g1566 ( 
.A1(n_1475),
.A2(n_1482),
.B(n_1471),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1470),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1508),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1541),
.B(n_1544),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1542),
.A2(n_1503),
.B(n_1474),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1458),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1553),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1548),
.A2(n_1475),
.B(n_1482),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1504),
.B(n_1466),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1526),
.B(n_1531),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1492),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1542),
.A2(n_1473),
.B(n_1523),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1466),
.B(n_1476),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1484),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1493),
.Y(n_1580)
);

NAND2x1p5_ASAP7_75t_L g1581 ( 
.A(n_1481),
.B(n_1546),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1541),
.B(n_1544),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1554),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1499),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1547),
.B(n_1556),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1519),
.A2(n_1526),
.B(n_1515),
.Y(n_1586)
);

OAI31xp33_ASAP7_75t_L g1587 ( 
.A1(n_1472),
.A2(n_1551),
.A3(n_1558),
.B(n_1543),
.Y(n_1587)
);

AOI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1555),
.A2(n_1472),
.B(n_1543),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1533),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1459),
.B(n_1502),
.Y(n_1590)
);

OAI211xp5_ASAP7_75t_L g1591 ( 
.A1(n_1555),
.A2(n_1486),
.B(n_1500),
.C(n_1491),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1551),
.A2(n_1558),
.B(n_1465),
.Y(n_1592)
);

OAI21xp33_ASAP7_75t_SL g1593 ( 
.A1(n_1488),
.A2(n_1512),
.B(n_1509),
.Y(n_1593)
);

INVx5_ASAP7_75t_L g1594 ( 
.A(n_1460),
.Y(n_1594)
);

OR2x6_ASAP7_75t_L g1595 ( 
.A(n_1501),
.B(n_1534),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1536),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1536),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1483),
.B(n_1490),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1485),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1487),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1507),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1511),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1479),
.B(n_1517),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1501),
.B(n_1488),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1498),
.B(n_1559),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1510),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1498),
.B(n_1549),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1550),
.Y(n_1608)
);

NOR2x1_ASAP7_75t_L g1609 ( 
.A(n_1517),
.B(n_1524),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1463),
.B(n_1557),
.Y(n_1610)
);

BUFx12f_ASAP7_75t_L g1611 ( 
.A(n_1562),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1605),
.B(n_1497),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1583),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1601),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1575),
.B(n_1518),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1565),
.B(n_1528),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1583),
.Y(n_1617)
);

INVxp67_ASAP7_75t_SL g1618 ( 
.A(n_1565),
.Y(n_1618)
);

NOR2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1561),
.B(n_1478),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1607),
.B(n_1514),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1568),
.B(n_1529),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1596),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1574),
.B(n_1520),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1574),
.B(n_1537),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1597),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1563),
.B(n_1535),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1598),
.B(n_1461),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1597),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1561),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1598),
.B(n_1467),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1578),
.B(n_1527),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1568),
.B(n_1516),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1606),
.B(n_1539),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1563),
.B(n_1586),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1586),
.B(n_1532),
.Y(n_1635)
);

NOR2x1_ASAP7_75t_L g1636 ( 
.A(n_1595),
.B(n_1532),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1584),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1586),
.B(n_1506),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1578),
.B(n_1460),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1586),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1584),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1571),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1585),
.B(n_1505),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1580),
.B(n_1464),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1636),
.A2(n_1573),
.B1(n_1592),
.B2(n_1591),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1642),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1636),
.A2(n_1573),
.B1(n_1609),
.B2(n_1592),
.Y(n_1647)
);

INVxp67_ASAP7_75t_SL g1648 ( 
.A(n_1618),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1642),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1615),
.B(n_1567),
.Y(n_1650)
);

AOI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1627),
.A2(n_1566),
.B1(n_1593),
.B2(n_1602),
.C(n_1587),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1635),
.B(n_1587),
.C(n_1593),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1632),
.B(n_1599),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1619),
.A2(n_1609),
.B1(n_1595),
.B2(n_1603),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1639),
.B(n_1589),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1611),
.A2(n_1595),
.B1(n_1521),
.B2(n_1552),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1611),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1635),
.A2(n_1588),
.B1(n_1582),
.B2(n_1569),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1615),
.B(n_1567),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1639),
.B(n_1589),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1615),
.B(n_1579),
.Y(n_1661)
);

BUFx3_ASAP7_75t_L g1662 ( 
.A(n_1611),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1642),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1637),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1629),
.A2(n_1590),
.B1(n_1604),
.B2(n_1595),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1613),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1620),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1629),
.A2(n_1595),
.B1(n_1590),
.B2(n_1604),
.C(n_1560),
.Y(n_1668)
);

INVx4_ASAP7_75t_L g1669 ( 
.A(n_1611),
.Y(n_1669)
);

AOI21xp33_ASAP7_75t_L g1670 ( 
.A1(n_1638),
.A2(n_1590),
.B(n_1604),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1614),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1637),
.Y(n_1672)
);

NAND2xp33_ASAP7_75t_R g1673 ( 
.A(n_1638),
.B(n_1522),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1626),
.B(n_1572),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1626),
.B(n_1600),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1626),
.B(n_1564),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1635),
.A2(n_1588),
.B1(n_1604),
.B2(n_1610),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1617),
.Y(n_1678)
);

OAI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1629),
.A2(n_1590),
.B1(n_1604),
.B2(n_1589),
.C(n_1570),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1627),
.A2(n_1581),
.B(n_1538),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1614),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1631),
.B(n_1576),
.Y(n_1682)
);

OAI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1629),
.A2(n_1590),
.B1(n_1638),
.B2(n_1632),
.C(n_1621),
.Y(n_1683)
);

OAI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1616),
.A2(n_1570),
.B1(n_1545),
.B2(n_1513),
.C(n_1581),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1617),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1612),
.Y(n_1686)
);

OAI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1616),
.A2(n_1570),
.B1(n_1581),
.B2(n_1608),
.C(n_1540),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1619),
.A2(n_1594),
.B1(n_1608),
.B2(n_1538),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1617),
.Y(n_1689)
);

OAI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1640),
.A2(n_1570),
.B(n_1577),
.C(n_1585),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1657),
.Y(n_1691)
);

INVx4_ASAP7_75t_SL g1692 ( 
.A(n_1657),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1653),
.B(n_1624),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1671),
.B(n_1641),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1646),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1657),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1649),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1664),
.Y(n_1698)
);

INVx4_ASAP7_75t_L g1699 ( 
.A(n_1669),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1663),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1647),
.B(n_1627),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1672),
.Y(n_1702)
);

OA21x2_ASAP7_75t_L g1703 ( 
.A1(n_1690),
.A2(n_1640),
.B(n_1680),
.Y(n_1703)
);

OA21x2_ASAP7_75t_L g1704 ( 
.A1(n_1680),
.A2(n_1625),
.B(n_1622),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1675),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1671),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1658),
.B(n_1624),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1666),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_1662),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1669),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1648),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1667),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1655),
.B(n_1620),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1658),
.B(n_1634),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1674),
.B(n_1624),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1661),
.B(n_1621),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1678),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1650),
.B(n_1643),
.Y(n_1718)
);

NOR2x1p5_ASAP7_75t_L g1719 ( 
.A(n_1652),
.B(n_1540),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1685),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1656),
.B(n_1489),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1655),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1659),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1689),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1651),
.B(n_1643),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1681),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1681),
.Y(n_1727)
);

INVx4_ASAP7_75t_SL g1728 ( 
.A(n_1656),
.Y(n_1728)
);

OA21x2_ASAP7_75t_L g1729 ( 
.A1(n_1670),
.A2(n_1622),
.B(n_1628),
.Y(n_1729)
);

NOR2xp67_ASAP7_75t_L g1730 ( 
.A(n_1714),
.B(n_1687),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1695),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1704),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1712),
.B(n_1660),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1710),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1712),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1728),
.B(n_1660),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1722),
.B(n_1620),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1695),
.Y(n_1738)
);

INVx3_ASAP7_75t_SL g1739 ( 
.A(n_1692),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1697),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1697),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1722),
.B(n_1623),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1713),
.B(n_1623),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1714),
.B(n_1634),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1713),
.B(n_1710),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1725),
.B(n_1652),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1707),
.B(n_1634),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1728),
.B(n_1630),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1721),
.B(n_1495),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1694),
.B(n_1623),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1700),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1711),
.B(n_1641),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1701),
.B(n_1705),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1694),
.B(n_1631),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1694),
.B(n_1728),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1700),
.B(n_1677),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1702),
.B(n_1682),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1698),
.B(n_1677),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1717),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1704),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1704),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1728),
.B(n_1631),
.Y(n_1762)
);

NOR2x1_ASAP7_75t_L g1763 ( 
.A(n_1699),
.B(n_1619),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1698),
.B(n_1676),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1703),
.B(n_1684),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1704),
.B(n_1630),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1723),
.B(n_1703),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1703),
.B(n_1630),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1719),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1703),
.B(n_1686),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1717),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1708),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1699),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1693),
.B(n_1683),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1727),
.B(n_1643),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1746),
.B(n_1691),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1746),
.B(n_1691),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1734),
.Y(n_1778)
);

NAND4xp25_ASAP7_75t_L g1779 ( 
.A(n_1730),
.B(n_1645),
.C(n_1654),
.D(n_1665),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1734),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1740),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1740),
.Y(n_1782)
);

A2O1A1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1730),
.A2(n_1645),
.B(n_1668),
.C(n_1679),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1735),
.B(n_1715),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1735),
.B(n_1716),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1741),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1741),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1734),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1772),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1731),
.Y(n_1790)
);

CKINVDCx20_ASAP7_75t_R g1791 ( 
.A(n_1749),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1735),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1736),
.B(n_1699),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1734),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1739),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1763),
.B(n_1692),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1731),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1736),
.B(n_1696),
.Y(n_1798)
);

NAND4xp25_ASAP7_75t_L g1799 ( 
.A(n_1769),
.B(n_1765),
.C(n_1753),
.D(n_1763),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1738),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1753),
.B(n_1718),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1736),
.B(n_1696),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1736),
.B(n_1727),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1738),
.Y(n_1804)
);

NAND2x1p5_ASAP7_75t_L g1805 ( 
.A(n_1734),
.B(n_1773),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1734),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1755),
.B(n_1706),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1756),
.B(n_1720),
.Y(n_1808)
);

NAND2x1_ASAP7_75t_L g1809 ( 
.A(n_1748),
.B(n_1706),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1751),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1769),
.B(n_1709),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1751),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1792),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1791),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1801),
.B(n_1784),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1805),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1812),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_L g1818 ( 
.A(n_1799),
.B(n_1765),
.C(n_1773),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1783),
.A2(n_1748),
.B1(n_1774),
.B2(n_1762),
.Y(n_1819)
);

NOR2x1_ASAP7_75t_L g1820 ( 
.A(n_1796),
.B(n_1748),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1779),
.A2(n_1748),
.B1(n_1774),
.B2(n_1745),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1812),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1791),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1798),
.B(n_1739),
.Y(n_1824)
);

CKINVDCx16_ASAP7_75t_R g1825 ( 
.A(n_1811),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1798),
.B(n_1739),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1787),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1787),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1801),
.A2(n_1745),
.B1(n_1768),
.B2(n_1762),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1802),
.B(n_1755),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1805),
.Y(n_1831)
);

OAI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1795),
.A2(n_1756),
.B1(n_1758),
.B2(n_1768),
.C(n_1767),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1776),
.B(n_1777),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1793),
.A2(n_1767),
.B1(n_1758),
.B2(n_1733),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1810),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1789),
.B(n_1743),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1802),
.B(n_1733),
.Y(n_1837)
);

INVxp67_ASAP7_75t_L g1838 ( 
.A(n_1805),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1784),
.B(n_1757),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1813),
.Y(n_1840)
);

OAI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1818),
.A2(n_1819),
.B1(n_1832),
.B2(n_1820),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1814),
.B(n_1778),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1813),
.Y(n_1843)
);

OAI322xp33_ASAP7_75t_L g1844 ( 
.A1(n_1815),
.A2(n_1786),
.A3(n_1782),
.B1(n_1781),
.B2(n_1808),
.C1(n_1785),
.C2(n_1780),
.Y(n_1844)
);

OAI21xp33_ASAP7_75t_L g1845 ( 
.A1(n_1821),
.A2(n_1793),
.B(n_1785),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1827),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1825),
.A2(n_1809),
.B1(n_1673),
.B2(n_1747),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1830),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1823),
.B(n_1807),
.Y(n_1849)
);

NOR3xp33_ASAP7_75t_L g1850 ( 
.A(n_1833),
.B(n_1780),
.C(n_1778),
.Y(n_1850)
);

OAI322xp33_ASAP7_75t_L g1851 ( 
.A1(n_1815),
.A2(n_1839),
.A3(n_1827),
.B1(n_1828),
.B2(n_1838),
.C1(n_1835),
.C2(n_1836),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1837),
.B(n_1788),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1834),
.A2(n_1794),
.B1(n_1788),
.B2(n_1806),
.C(n_1800),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1828),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1817),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1824),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1830),
.B(n_1803),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1822),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1830),
.B(n_1794),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1837),
.A2(n_1807),
.B1(n_1803),
.B2(n_1806),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1842),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1840),
.B(n_1843),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1852),
.B(n_1839),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1856),
.B(n_1824),
.Y(n_1864)
);

XNOR2x1_ASAP7_75t_L g1865 ( 
.A(n_1841),
.B(n_1826),
.Y(n_1865)
);

INVx2_ASAP7_75t_SL g1866 ( 
.A(n_1859),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1848),
.B(n_1829),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1859),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1849),
.B(n_1826),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1845),
.B(n_1831),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1857),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1846),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1854),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1869),
.B(n_1871),
.Y(n_1874)
);

OAI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1865),
.A2(n_1850),
.B(n_1847),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1866),
.B(n_1860),
.Y(n_1876)
);

NOR4xp25_ASAP7_75t_L g1877 ( 
.A(n_1862),
.B(n_1851),
.C(n_1844),
.D(n_1858),
.Y(n_1877)
);

OAI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1870),
.A2(n_1853),
.B(n_1816),
.C(n_1855),
.Y(n_1878)
);

AOI222xp33_ASAP7_75t_L g1879 ( 
.A1(n_1861),
.A2(n_1816),
.B1(n_1766),
.B2(n_1761),
.C1(n_1760),
.C2(n_1732),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1868),
.B(n_1750),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1864),
.A2(n_1809),
.B1(n_1790),
.B2(n_1804),
.Y(n_1881)
);

NAND4xp25_ASAP7_75t_L g1882 ( 
.A(n_1864),
.B(n_1808),
.C(n_1797),
.D(n_1688),
.Y(n_1882)
);

AOI32xp33_ASAP7_75t_L g1883 ( 
.A1(n_1867),
.A2(n_1766),
.A3(n_1732),
.B1(n_1770),
.B2(n_1760),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1863),
.B(n_1873),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1884),
.Y(n_1885)
);

NAND2xp33_ASAP7_75t_R g1886 ( 
.A(n_1874),
.B(n_1862),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1880),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1875),
.A2(n_1872),
.B1(n_1732),
.B2(n_1760),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1876),
.B(n_1750),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1878),
.A2(n_1732),
.B1(n_1761),
.B2(n_1747),
.Y(n_1890)
);

OAI21xp33_ASAP7_75t_L g1891 ( 
.A1(n_1877),
.A2(n_1770),
.B(n_1752),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1889),
.B(n_1881),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1887),
.B(n_1883),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1885),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1891),
.B(n_1882),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1888),
.B(n_1692),
.Y(n_1896)
);

NAND2xp33_ASAP7_75t_L g1897 ( 
.A(n_1890),
.B(n_1752),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1892),
.B(n_1879),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1896),
.B(n_1895),
.Y(n_1899)
);

AOI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1897),
.A2(n_1890),
.B1(n_1886),
.B2(n_1761),
.C(n_1771),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1893),
.A2(n_1771),
.B(n_1759),
.Y(n_1901)
);

NOR2x1_ASAP7_75t_L g1902 ( 
.A(n_1894),
.B(n_1759),
.Y(n_1902)
);

NOR4xp75_ASAP7_75t_SL g1903 ( 
.A(n_1899),
.B(n_1692),
.C(n_1644),
.D(n_1633),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1902),
.Y(n_1904)
);

NAND3xp33_ASAP7_75t_L g1905 ( 
.A(n_1900),
.B(n_1744),
.C(n_1729),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1903),
.B(n_1898),
.Y(n_1906)
);

AOI22x1_ASAP7_75t_L g1907 ( 
.A1(n_1906),
.A2(n_1904),
.B1(n_1901),
.B2(n_1905),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1907),
.Y(n_1908)
);

OA21x2_ASAP7_75t_L g1909 ( 
.A1(n_1907),
.A2(n_1744),
.B(n_1775),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1908),
.A2(n_1764),
.B1(n_1757),
.B2(n_1726),
.Y(n_1910)
);

XNOR2xp5_ASAP7_75t_L g1911 ( 
.A(n_1909),
.B(n_1737),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1911),
.A2(n_1910),
.B1(n_1909),
.B2(n_1764),
.Y(n_1912)
);

AOI22x1_ASAP7_75t_L g1913 ( 
.A1(n_1911),
.A2(n_1909),
.B1(n_1530),
.B2(n_1494),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1913),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1914),
.A2(n_1912),
.B1(n_1530),
.B2(n_1494),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1737),
.B(n_1742),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1775),
.B1(n_1726),
.B2(n_1706),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1917),
.A2(n_1726),
.B1(n_1742),
.B2(n_1754),
.Y(n_1918)
);

OA22x2_ASAP7_75t_L g1919 ( 
.A1(n_1918),
.A2(n_1754),
.B1(n_1720),
.B2(n_1724),
.Y(n_1919)
);


endmodule