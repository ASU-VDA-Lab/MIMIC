module fake_jpeg_22026_n_328 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_37),
.B1(n_26),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_50),
.A2(n_67),
.B1(n_73),
.B2(n_24),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_52),
.B(n_57),
.Y(n_101)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_62),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_21),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_77),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_63),
.Y(n_115)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_34),
.B1(n_35),
.B2(n_17),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_34),
.B1(n_17),
.B2(n_35),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_74),
.B1(n_80),
.B2(n_18),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_79),
.Y(n_86)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_34),
.B1(n_27),
.B2(n_21),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_36),
.B1(n_27),
.B2(n_21),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_27),
.Y(n_76)
);

NOR2x1_ASAP7_75t_R g92 ( 
.A(n_76),
.B(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_33),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_83),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_23),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_95),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_33),
.B1(n_30),
.B2(n_20),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_18),
.B(n_30),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_90),
.A2(n_92),
.B(n_104),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_97),
.B1(n_108),
.B2(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_20),
.B1(n_32),
.B2(n_25),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_98),
.A2(n_105),
.B1(n_64),
.B2(n_72),
.Y(n_136)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_102),
.Y(n_132)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_22),
.B1(n_15),
.B2(n_14),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_0),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_19),
.B(n_24),
.C(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_106),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_24),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_63),
.C(n_57),
.Y(n_124)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_23),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_0),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_8),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_28),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_28),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_28),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_150),
.B1(n_114),
.B2(n_104),
.Y(n_155)
);

BUFx8_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_115),
.C(n_81),
.Y(n_165)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_71),
.B(n_70),
.C(n_52),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_152),
.B(n_83),
.Y(n_169)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_140),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_137),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_138),
.B1(n_139),
.B2(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_58),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_55),
.B1(n_58),
.B2(n_53),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_55),
.B1(n_51),
.B2(n_60),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_145),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_51),
.B1(n_60),
.B2(n_28),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_86),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_94),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_149),
.A2(n_102),
.B1(n_91),
.B2(n_110),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_154),
.A2(n_164),
.B1(n_174),
.B2(n_175),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_173),
.B1(n_184),
.B2(n_142),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_93),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_112),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_171),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_170),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_109),
.B1(n_92),
.B2(n_104),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_152),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_169),
.A2(n_177),
.B(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_88),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_180),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_135),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_124),
.A2(n_82),
.B1(n_117),
.B2(n_118),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_91),
.B1(n_98),
.B2(n_85),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_183),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_139),
.B(n_138),
.C(n_137),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_130),
.A2(n_121),
.B(n_131),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_130),
.A2(n_1),
.B(n_2),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_144),
.B(n_132),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_1),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_3),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_119),
.B1(n_131),
.B2(n_142),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_3),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_134),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_188),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_191),
.B(n_198),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_195),
.B(n_210),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_132),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_214),
.C(n_153),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_141),
.B(n_133),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_161),
.B1(n_174),
.B2(n_164),
.Y(n_218)
);

CKINVDCx10_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_146),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_205),
.B(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_182),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_168),
.B(n_149),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_161),
.A2(n_133),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_177),
.B1(n_155),
.B2(n_171),
.Y(n_225)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_212),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_SL g211 ( 
.A1(n_168),
.A2(n_10),
.A3(n_16),
.B1(n_15),
.B2(n_13),
.C1(n_12),
.C2(n_8),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_123),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_162),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_158),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_221),
.B(n_204),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_224),
.B1(n_209),
.B2(n_200),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_158),
.B(n_169),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_226),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_196),
.A2(n_175),
.B1(n_185),
.B2(n_156),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_231),
.B1(n_191),
.B2(n_198),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_192),
.B(n_195),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_177),
.B1(n_184),
.B2(n_183),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_194),
.C(n_186),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_236),
.Y(n_250)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_157),
.C(n_160),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_215),
.Y(n_247)
);

AOI211xp5_ASAP7_75t_SL g242 ( 
.A1(n_203),
.A2(n_184),
.B(n_176),
.C(n_157),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_242),
.A2(n_206),
.B1(n_212),
.B2(n_207),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

NOR4xp25_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_200),
.C(n_202),
.D(n_213),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_227),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_257),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_259),
.B(n_262),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_189),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_258),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_219),
.B1(n_242),
.B2(n_217),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_217),
.A2(n_227),
.B1(n_231),
.B2(n_225),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_154),
.B1(n_166),
.B2(n_123),
.Y(n_281)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_202),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_221),
.A2(n_187),
.B1(n_184),
.B2(n_204),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_260),
.B(n_261),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_222),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_240),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_226),
.C(n_236),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_270),
.C(n_272),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_268),
.A2(n_253),
.B1(n_245),
.B2(n_11),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_269),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_229),
.C(n_216),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_241),
.C(n_220),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_184),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_277),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_234),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_239),
.C(n_233),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_279),
.C(n_262),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_239),
.C(n_233),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_249),
.B(n_228),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_280),
.B(n_263),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_271),
.B1(n_264),
.B2(n_279),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_292),
.B1(n_270),
.B2(n_272),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_268),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_265),
.B(n_249),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_259),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_294),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_295),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_293),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_253),
.C(n_255),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_252),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_290),
.A2(n_273),
.B(n_276),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_293),
.B(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_303),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_274),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_266),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.C(n_289),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_277),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_291),
.Y(n_306)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_296),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_298),
.B(n_305),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_282),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_123),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_282),
.C(n_123),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_297),
.A2(n_16),
.B1(n_12),
.B2(n_11),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_317),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_311),
.B(n_299),
.Y(n_317)
);

AOI31xp67_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_8),
.A3(n_4),
.B(n_5),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_SL g320 ( 
.A1(n_316),
.A2(n_312),
.B(n_307),
.C(n_16),
.Y(n_320)
);

AOI31xp33_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_321),
.A3(n_3),
.B(n_5),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_318),
.C(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);

OAI221xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_315),
.B1(n_324),
.B2(n_314),
.C(n_7),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_5),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_6),
.B(n_7),
.Y(n_328)
);


endmodule